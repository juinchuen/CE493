VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pid
  CLASS BLOCK ;
  FOREIGN pid ;
  ORIGIN 0.000 0.000 ;
  SIZE 442.700 BY 453.420 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 440.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 440.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 440.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 437.240 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 437.240 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 437.240 337.990 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 440.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 440.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 440.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 437.240 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 437.240 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 437.240 334.690 ;
    END
  END VPWR
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 357.510 449.420 357.790 453.420 ;
    END
  END clock
  PIN iterate_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 360.730 449.420 361.010 453.420 ;
    END
  END iterate_enable
  PIN measurement[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END measurement[0]
  PIN measurement[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END measurement[10]
  PIN measurement[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END measurement[11]
  PIN measurement[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END measurement[12]
  PIN measurement[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END measurement[13]
  PIN measurement[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END measurement[14]
  PIN measurement[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END measurement[15]
  PIN measurement[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END measurement[16]
  PIN measurement[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END measurement[17]
  PIN measurement[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END measurement[18]
  PIN measurement[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END measurement[1]
  PIN measurement[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END measurement[2]
  PIN measurement[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END measurement[3]
  PIN measurement[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END measurement[4]
  PIN measurement[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END measurement[5]
  PIN measurement[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END measurement[6]
  PIN measurement[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END measurement[7]
  PIN measurement[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END measurement[8]
  PIN measurement[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END measurement[9]
  PIN out_clocked[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 438.700 180.240 442.700 180.840 ;
    END
  END out_clocked[0]
  PIN out_clocked[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 438.700 200.640 442.700 201.240 ;
    END
  END out_clocked[10]
  PIN out_clocked[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 438.700 221.040 442.700 221.640 ;
    END
  END out_clocked[11]
  PIN out_clocked[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 438.700 210.840 442.700 211.440 ;
    END
  END out_clocked[12]
  PIN out_clocked[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 438.700 302.640 442.700 303.240 ;
    END
  END out_clocked[13]
  PIN out_clocked[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 438.700 319.640 442.700 320.240 ;
    END
  END out_clocked[14]
  PIN out_clocked[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 438.700 309.440 442.700 310.040 ;
    END
  END out_clocked[15]
  PIN out_clocked[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 438.700 326.440 442.700 327.040 ;
    END
  END out_clocked[16]
  PIN out_clocked[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 438.700 323.040 442.700 323.640 ;
    END
  END out_clocked[17]
  PIN out_clocked[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 438.700 312.840 442.700 313.440 ;
    END
  END out_clocked[18]
  PIN out_clocked[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 438.700 204.040 442.700 204.640 ;
    END
  END out_clocked[1]
  PIN out_clocked[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 438.700 207.440 442.700 208.040 ;
    END
  END out_clocked[2]
  PIN out_clocked[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 438.700 190.440 442.700 191.040 ;
    END
  END out_clocked[3]
  PIN out_clocked[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 438.700 214.240 442.700 214.840 ;
    END
  END out_clocked[4]
  PIN out_clocked[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 438.700 187.040 442.700 187.640 ;
    END
  END out_clocked[5]
  PIN out_clocked[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 438.700 217.640 442.700 218.240 ;
    END
  END out_clocked[6]
  PIN out_clocked[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 438.700 183.640 442.700 184.240 ;
    END
  END out_clocked[7]
  PIN out_clocked[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 438.700 193.840 442.700 194.440 ;
    END
  END out_clocked[8]
  PIN out_clocked[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 438.700 197.240 442.700 197.840 ;
    END
  END out_clocked[9]
  PIN reg_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END reg_addr[0]
  PIN reg_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END reg_addr[10]
  PIN reg_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END reg_addr[11]
  PIN reg_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END reg_addr[12]
  PIN reg_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END reg_addr[13]
  PIN reg_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END reg_addr[14]
  PIN reg_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END reg_addr[15]
  PIN reg_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END reg_addr[16]
  PIN reg_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END reg_addr[17]
  PIN reg_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END reg_addr[18]
  PIN reg_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END reg_addr[2]
  PIN reg_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END reg_addr[3]
  PIN reg_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END reg_addr[4]
  PIN reg_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END reg_addr[5]
  PIN reg_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END reg_addr[6]
  PIN reg_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END reg_addr[7]
  PIN reg_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END reg_addr[8]
  PIN reg_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END reg_addr[9]
  PIN reg_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END reg_data[0]
  PIN reg_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END reg_data[10]
  PIN reg_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END reg_data[11]
  PIN reg_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END reg_data[12]
  PIN reg_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END reg_data[13]
  PIN reg_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END reg_data[14]
  PIN reg_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END reg_data[15]
  PIN reg_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END reg_data[16]
  PIN reg_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END reg_data[17]
  PIN reg_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END reg_data[18]
  PIN reg_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END reg_data[1]
  PIN reg_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END reg_data[2]
  PIN reg_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END reg_data[3]
  PIN reg_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END reg_data[4]
  PIN reg_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END reg_data[5]
  PIN reg_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END reg_data[6]
  PIN reg_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END reg_data[7]
  PIN reg_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END reg_data[8]
  PIN reg_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END reg_data[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 438.700 224.440 442.700 225.040 ;
    END
  END reset
  PIN target[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END target[0]
  PIN target[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END target[10]
  PIN target[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END target[11]
  PIN target[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END target[12]
  PIN target[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END target[13]
  PIN target[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END target[14]
  PIN target[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END target[15]
  PIN target[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END target[16]
  PIN target[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END target[17]
  PIN target[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END target[18]
  PIN target[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END target[1]
  PIN target[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END target[2]
  PIN target[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END target[3]
  PIN target[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END target[4]
  PIN target[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END target[5]
  PIN target[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END target[6]
  PIN target[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END target[7]
  PIN target[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END target[8]
  PIN target[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END target[9]
  PIN write_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END write_enable
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 437.000 440.725 ;
      LAYER met1 ;
        RECT 4.670 9.900 437.390 440.880 ;
      LAYER met2 ;
        RECT 4.690 449.140 357.230 449.420 ;
        RECT 358.070 449.140 360.450 449.420 ;
        RECT 361.290 449.140 437.370 449.420 ;
        RECT 4.690 4.280 437.370 449.140 ;
        RECT 4.690 4.000 167.250 4.280 ;
        RECT 168.090 4.000 170.470 4.280 ;
        RECT 171.310 4.000 173.690 4.280 ;
        RECT 174.530 4.000 176.910 4.280 ;
        RECT 177.750 4.000 180.130 4.280 ;
        RECT 180.970 4.000 183.350 4.280 ;
        RECT 184.190 4.000 186.570 4.280 ;
        RECT 187.410 4.000 189.790 4.280 ;
        RECT 190.630 4.000 193.010 4.280 ;
        RECT 193.850 4.000 196.230 4.280 ;
        RECT 197.070 4.000 199.450 4.280 ;
        RECT 200.290 4.000 202.670 4.280 ;
        RECT 203.510 4.000 205.890 4.280 ;
        RECT 206.730 4.000 209.110 4.280 ;
        RECT 209.950 4.000 212.330 4.280 ;
        RECT 213.170 4.000 215.550 4.280 ;
        RECT 216.390 4.000 218.770 4.280 ;
        RECT 219.610 4.000 221.990 4.280 ;
        RECT 222.830 4.000 225.210 4.280 ;
        RECT 226.050 4.000 228.430 4.280 ;
        RECT 229.270 4.000 231.650 4.280 ;
        RECT 232.490 4.000 234.870 4.280 ;
        RECT 235.710 4.000 238.090 4.280 ;
        RECT 238.930 4.000 241.310 4.280 ;
        RECT 242.150 4.000 244.530 4.280 ;
        RECT 245.370 4.000 247.750 4.280 ;
        RECT 248.590 4.000 250.970 4.280 ;
        RECT 251.810 4.000 254.190 4.280 ;
        RECT 255.030 4.000 257.410 4.280 ;
        RECT 258.250 4.000 260.630 4.280 ;
        RECT 261.470 4.000 263.850 4.280 ;
        RECT 264.690 4.000 267.070 4.280 ;
        RECT 267.910 4.000 270.290 4.280 ;
        RECT 271.130 4.000 273.510 4.280 ;
        RECT 274.350 4.000 276.730 4.280 ;
        RECT 277.570 4.000 279.950 4.280 ;
        RECT 280.790 4.000 283.170 4.280 ;
        RECT 284.010 4.000 286.390 4.280 ;
        RECT 287.230 4.000 289.610 4.280 ;
        RECT 290.450 4.000 437.370 4.280 ;
      LAYER met3 ;
        RECT 3.990 409.040 438.700 440.805 ;
        RECT 4.400 407.640 438.700 409.040 ;
        RECT 3.990 405.640 438.700 407.640 ;
        RECT 4.400 404.240 438.700 405.640 ;
        RECT 3.990 402.240 438.700 404.240 ;
        RECT 4.400 400.840 438.700 402.240 ;
        RECT 3.990 398.840 438.700 400.840 ;
        RECT 4.400 397.440 438.700 398.840 ;
        RECT 3.990 395.440 438.700 397.440 ;
        RECT 4.400 394.040 438.700 395.440 ;
        RECT 3.990 392.040 438.700 394.040 ;
        RECT 4.400 390.640 438.700 392.040 ;
        RECT 3.990 388.640 438.700 390.640 ;
        RECT 4.400 387.240 438.700 388.640 ;
        RECT 3.990 385.240 438.700 387.240 ;
        RECT 4.400 383.840 438.700 385.240 ;
        RECT 3.990 381.840 438.700 383.840 ;
        RECT 4.400 380.440 438.700 381.840 ;
        RECT 3.990 378.440 438.700 380.440 ;
        RECT 4.400 377.040 438.700 378.440 ;
        RECT 3.990 361.440 438.700 377.040 ;
        RECT 4.400 360.040 438.700 361.440 ;
        RECT 3.990 358.040 438.700 360.040 ;
        RECT 4.400 356.640 438.700 358.040 ;
        RECT 3.990 354.640 438.700 356.640 ;
        RECT 4.400 353.240 438.700 354.640 ;
        RECT 3.990 351.240 438.700 353.240 ;
        RECT 4.400 349.840 438.700 351.240 ;
        RECT 3.990 327.440 438.700 349.840 ;
        RECT 3.990 326.040 438.300 327.440 ;
        RECT 3.990 324.040 438.700 326.040 ;
        RECT 3.990 322.640 438.300 324.040 ;
        RECT 3.990 320.640 438.700 322.640 ;
        RECT 4.400 319.240 438.300 320.640 ;
        RECT 3.990 317.240 438.700 319.240 ;
        RECT 4.400 315.840 438.700 317.240 ;
        RECT 3.990 313.840 438.700 315.840 ;
        RECT 4.400 312.440 438.300 313.840 ;
        RECT 3.990 310.440 438.700 312.440 ;
        RECT 4.400 309.040 438.300 310.440 ;
        RECT 3.990 303.640 438.700 309.040 ;
        RECT 3.990 302.240 438.300 303.640 ;
        RECT 3.990 300.240 438.700 302.240 ;
        RECT 4.400 298.840 438.700 300.240 ;
        RECT 3.990 296.840 438.700 298.840 ;
        RECT 4.400 295.440 438.700 296.840 ;
        RECT 3.990 293.440 438.700 295.440 ;
        RECT 4.400 292.040 438.700 293.440 ;
        RECT 3.990 290.040 438.700 292.040 ;
        RECT 4.400 288.640 438.700 290.040 ;
        RECT 3.990 256.040 438.700 288.640 ;
        RECT 4.400 254.640 438.700 256.040 ;
        RECT 3.990 252.640 438.700 254.640 ;
        RECT 4.400 251.240 438.700 252.640 ;
        RECT 3.990 245.840 438.700 251.240 ;
        RECT 4.400 244.440 438.700 245.840 ;
        RECT 3.990 242.440 438.700 244.440 ;
        RECT 4.400 241.040 438.700 242.440 ;
        RECT 3.990 235.640 438.700 241.040 ;
        RECT 4.400 234.240 438.700 235.640 ;
        RECT 3.990 232.240 438.700 234.240 ;
        RECT 4.400 230.840 438.700 232.240 ;
        RECT 3.990 228.840 438.700 230.840 ;
        RECT 4.400 227.440 438.700 228.840 ;
        RECT 3.990 225.440 438.700 227.440 ;
        RECT 4.400 224.040 438.300 225.440 ;
        RECT 3.990 222.040 438.700 224.040 ;
        RECT 4.400 220.640 438.300 222.040 ;
        RECT 3.990 218.640 438.700 220.640 ;
        RECT 4.400 217.240 438.300 218.640 ;
        RECT 3.990 215.240 438.700 217.240 ;
        RECT 4.400 213.840 438.300 215.240 ;
        RECT 3.990 211.840 438.700 213.840 ;
        RECT 4.400 210.440 438.300 211.840 ;
        RECT 3.990 208.440 438.700 210.440 ;
        RECT 3.990 207.040 438.300 208.440 ;
        RECT 3.990 205.040 438.700 207.040 ;
        RECT 3.990 203.640 438.300 205.040 ;
        RECT 3.990 201.640 438.700 203.640 ;
        RECT 3.990 200.240 438.300 201.640 ;
        RECT 3.990 198.240 438.700 200.240 ;
        RECT 3.990 196.840 438.300 198.240 ;
        RECT 3.990 194.840 438.700 196.840 ;
        RECT 3.990 193.440 438.300 194.840 ;
        RECT 3.990 191.440 438.700 193.440 ;
        RECT 3.990 190.040 438.300 191.440 ;
        RECT 3.990 188.040 438.700 190.040 ;
        RECT 3.990 186.640 438.300 188.040 ;
        RECT 3.990 184.640 438.700 186.640 ;
        RECT 3.990 183.240 438.300 184.640 ;
        RECT 3.990 181.240 438.700 183.240 ;
        RECT 4.400 179.840 438.300 181.240 ;
        RECT 3.990 177.840 438.700 179.840 ;
        RECT 4.400 176.440 438.700 177.840 ;
        RECT 3.990 174.440 438.700 176.440 ;
        RECT 4.400 173.040 438.700 174.440 ;
        RECT 3.990 171.040 438.700 173.040 ;
        RECT 4.400 169.640 438.700 171.040 ;
        RECT 3.990 10.715 438.700 169.640 ;
      LAYER met4 ;
        RECT 15.935 11.735 20.640 407.825 ;
        RECT 23.040 11.735 23.940 407.825 ;
        RECT 26.340 11.735 174.240 407.825 ;
        RECT 176.640 11.735 177.540 407.825 ;
        RECT 179.940 11.735 327.840 407.825 ;
        RECT 330.240 11.735 331.140 407.825 ;
        RECT 333.540 11.735 408.185 407.825 ;
  END
END pid
END LIBRARY

