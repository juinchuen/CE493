* NGSPICE file created from fpga_wrapper.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.136 ps=1.1 w=0.65 l=0.15
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258 ps=1.45 w=0.65 l=0.15
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.1 as=0.111 ps=1.37 w=0.42 l=0.15
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.258 pd=1.45 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X2 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.965 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.157 ps=1.32 w=1 l=0.15
X4 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X5 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X9 a_381_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0683 ps=0.86 w=0.65 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.185 ps=1.87 w=0.65 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
X0 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0991 ps=0.955 w=0.65 l=0.15
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X7 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X12 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X17 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.272 ps=2.56 w=1 l=0.15
X15 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X17 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X19 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X24 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.257 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X30 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X35 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X38 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.134 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.118 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.126 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 VPWR a_38_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A1 a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X2 X a_38_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X3 a_141_47# B2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_497_297# A2 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.387 ps=1.77 w=1 l=0.15
X5 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR C1 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.325 ps=2.65 w=1 l=0.15
X7 a_237_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.112 pd=1.23 as=0.165 ps=1.33 w=1 l=0.15
X8 a_38_47# B2 a_237_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.387 pd=1.77 as=0.112 ps=1.23 w=1 l=0.15
X9 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 X a_38_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_141_47# C1 a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.237 ps=2.03 w=0.65 l=0.15
X12 VGND a_38_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_225_47# B1 a_141_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
X0 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X5 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X21 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X35 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X36 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 VPWR A3 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X2 a_352_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.21 ps=1.29 w=0.65 l=0.15
X3 a_549_47# A1 a_21_199# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.08 as=0.107 ps=0.98 w=0.65 l=0.15
X4 X a_21_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_21_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.21 pd=1.29 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.14 ps=1.08 w=0.65 l=0.15
X7 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X8 a_299_297# B1 a_21_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_21_199# B2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND A3 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR a_21_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 X a_21_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_21_199# B1 a_352_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.115 ps=1 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.338 pd=1.67 as=0.135 ps=1.27 w=1 l=0.15
X5 a_1249_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_1249_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.252 pd=1.5 as=0.338 ps=1.67 w=1 l=0.15
X12 a_803_47# A2 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X16 a_803_47# A2 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X20 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X21 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 a_1249_47# A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.133 ps=1.06 w=0.65 l=0.15
X23 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 a_1249_47# A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.252 ps=1.5 w=1 l=0.15
X28 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X30 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X32 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 VGND A3 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X37 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 VGND A3 a_1249_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.106 ps=0.975 w=0.65 l=0.15
X6 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X8 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.275 ps=2.55 w=1 l=0.15
X10 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.162 ps=1.33 w=1 l=0.15
X11 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X18 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 Y A1 a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.119 ps=1.01 w=0.65 l=0.15
X1 a_181_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.0683 ps=0.86 w=0.65 l=0.15
X2 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.106 ps=0.975 w=0.65 l=0.15
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.162 ps=1.33 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.153 ps=1.3 w=1 l=0.15
X6 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_381_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.0683 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
X0 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VGND D_N a_1191_21# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_803_297# a_1191_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_445_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y a_1191_21# a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_803_297# a_1191_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 Y a_1191_21# a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X12 Y a_1191_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR D_N a_1191_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_27_297# B a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 VGND a_1191_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VGND a_1191_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 a_445_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_803_297# C a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 a_27_297# B a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_445_297# C a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_803_297# C a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 Y a_1191_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X32 a_445_297# C a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X33 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.412 pd=1.83 as=0.105 ps=1.21 w=1 l=0.15
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.201 ps=1.92 w=0.65 l=0.15
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0991 ps=0.955 w=0.65 l=0.15
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.412 ps=1.83 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.1 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X16 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X17 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X20 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X21 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X22 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 VGND A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND B2 a_1053_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_804_297# B1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=1.69 as=0.135 ps=1.27 w=1 l=0.15
X3 a_79_21# A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_445_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_804_297# C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_445_297# B1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_1053_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_79_21# C1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X10 a_1053_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_445_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_804_297# B2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X18 a_79_21# B1 a_1053_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_445_297# B2 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.345 ps=1.69 w=1 l=0.15
X21 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 a_445_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 a_445_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VPWR A1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X26 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_56_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR A2 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.101 ps=0.96 w=0.65 l=0.15
X3 a_139_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.266 ps=2.12 w=0.65 l=0.15
X4 a_311_297# B1 a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X5 Y C1 a_311_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X7 Y A1 a_139_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.16 ps=1.32 w=1 l=0.15
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.4 ps=1.8 w=1 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0894 ps=0.925 w=0.65 l=0.15
X3 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_470_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.138 ps=1.27 w=1 l=0.15
X6 a_384_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X7 a_384_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.104 ps=0.97 w=0.65 l=0.15
X8 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_301_47# B2 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND A2 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X2 a_383_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.39 ps=1.78 w=1 l=0.15
X3 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X4 a_301_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X8 VPWR A1 a_579_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X9 a_81_21# B1 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_579_297# A2 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X11 a_81_21# B2 a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.105 ps=1.21 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.127 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=1 w=0.65 l=0.15
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.156 ps=1.36 w=1 l=0.15
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.156 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0852 ps=0.925 w=0.42 l=0.15
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.108 ps=1.36 w=0.42 l=0.15
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.269 pd=2.12 as=0.0921 ps=0.99 w=0.42 l=0.15
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0921 pd=0.99 as=0.109 ps=1.36 w=0.42 l=0.15
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0852 pd=0.925 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0901 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0901 ps=0.995 w=0.42 l=0.15
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.151 ps=1.28 w=0.42 l=0.15
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.151 pd=1.28 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
X0 Y a_251_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y a_251_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X5 VGND a_251_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 VPWR B_N a_251_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X8 VGND B_N a_251_21# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_27_297# a_251_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_286_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2 a_286_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.185 ps=1.87 w=0.65 l=0.15
X3 Y A2 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 VGND A1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X5 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.185 ps=1.87 w=0.65 l=0.15
X6 VGND A2 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 a_487_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_27_47# B1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR A1 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X13 a_487_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X14 a_286_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.151 ps=1.35 w=1 l=0.15
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.151 pd=1.35 as=0.0744 ps=0.815 w=0.42 l=0.15
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.13 ps=1.11 w=0.65 l=0.15
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.11 as=0.0536 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
.ends

.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.127 ps=1.04 w=0.65 l=0.15
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.133 ps=1.06 w=0.65 l=0.15
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.107 ps=0.98 w=0.65 l=0.15
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.213 ps=1.42 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.146 ps=1.34 w=0.42 l=0.15
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0672 ps=0.74 w=0.42 l=0.15
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.209 pd=1.35 as=0.129 ps=1.18 w=0.42 l=0.15
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.209 ps=1.35 w=0.42 l=0.15
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0662 pd=0.735 as=0.0986 ps=0.98 w=0.42 l=0.15
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.0986 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.157 ps=1.17 w=0.42 l=0.15
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
X0 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 a_471_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=2.84 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_27_47# C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X8 a_277_47# B a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.135 ps=1.27 w=1 l=0.15
X10 Y A a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_277_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X13 a_471_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.135 ps=1.07 w=0.65 l=0.15
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.112 ps=0.995 w=0.65 l=0.15
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125 ps=1.03 w=0.65 l=0.15
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.07 as=0.106 ps=0.975 w=0.65 l=0.15
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.207 ps=1.41 w=1 l=0.15
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.207 pd=1.41 as=0.162 ps=1.33 w=1 l=0.15
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.142 ps=1.28 w=1 l=0.15
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.305 ps=1.61 w=1 l=0.15
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.102 ps=0.99 w=0.65 l=0.15
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.111 ps=1.37 w=0.42 l=0.15
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# a_419_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_419_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VGND a_419_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 Y a_419_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 Y a_419_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VGND B_N a_419_21# VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.182 ps=1.86 w=0.65 l=0.15
X13 Y a_419_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VPWR B_N a_419_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.27 ps=2.54 w=1 l=0.15
X15 a_27_297# a_419_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 Y a_419_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.153 ps=1.3 w=1 l=0.15
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.127 ps=1.25 w=1 l=0.15
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.178 ps=1.4 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_806_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.101 ps=0.96 w=0.65 l=0.15
X3 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_47# B1 a_1314_47# VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=2.09 as=0.104 ps=0.97 w=0.65 l=0.15
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X17 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0943 ps=0.94 w=0.65 l=0.15
X19 Y C1 a_978_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 Y C1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X22 a_27_47# B1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 a_806_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.675 pd=3.35 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.091 ps=0.93 w=0.65 l=0.15
X27 a_978_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
X28 a_1314_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X31 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.167 ps=1.39 w=1 l=0.15
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.112 ps=1.04 w=0.65 l=0.15
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.127 ps=1.04 w=0.65 l=0.15
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.184 ps=1.22 w=0.65 l=0.15
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.184 pd=1.22 as=0.161 ps=1.14 w=0.65 l=0.15
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.161 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0452 pd=0.635 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.064 pd=0.725 as=0.0452 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.064 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X1 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.157 ps=1.32 w=1 l=0.15
X3 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.965 w=0.65 l=0.15
X6 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X8 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X9 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X10 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 a_281_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1 a_281_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X9 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.127 ps=1.04 w=0.65 l=0.15
X10 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.198 ps=1.26 w=0.65 l=0.15
X11 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.127 ps=1.04 w=0.65 l=0.15
X12 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 Y A3 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.195 ps=1.39 w=1 l=0.15
X15 a_27_297# A2 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_397_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR B1_N a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X2 Y A2 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VGND A2 a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VGND A1 a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_28_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X6 Y a_28_297# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR a_28_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 a_397_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X9 a_229_47# a_28_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y a_28_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X11 a_229_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_229_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR A1 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X7 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X11 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X12 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X14 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X15 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X16 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X19 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.155 ps=1.31 w=1 l=0.15
X20 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X21 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X22 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X23 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.33 w=1 l=0.15
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 a_316_297# C1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.172 ps=1.35 w=1 l=0.15
X1 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.481 ps=2.78 w=0.65 l=0.15
X2 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.02 as=0.125 ps=1.03 w=0.65 l=0.15
X3 a_420_297# B1 a_316_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=1.58 as=0.185 ps=1.37 w=1 l=0.15
X4 VPWR A1 a_420_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.29 ps=1.58 w=1 l=0.15
X5 VGND A2 a_568_47# VNB sky130_fd_pr__nfet_01v8 ad=0.192 pd=1.89 as=0.0845 ps=0.91 w=0.65 l=0.15
X6 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.192 pd=1.24 as=0.12 ps=1.02 w=0.65 l=0.15
X7 a_420_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.138 ps=1.27 w=1 l=0.15
X8 a_217_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.755 ps=3.51 w=1 l=0.15
X9 a_568_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0845 pd=0.91 as=0.192 ps=1.24 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
X0 Y a_74_47# a_265_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B_N a_74_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.39 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_265_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.157 ps=1.39 w=1 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X4 VGND B_N a_74_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VGND a_74_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND A1 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_926_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A3 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X4 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A2 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_926_297# A2 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_102_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X8 a_496_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0975 ps=0.95 w=0.65 l=0.15
X10 a_102_21# B1 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X11 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.15 ps=1.3 w=1 l=0.15
X14 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X15 a_672_297# A3 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_496_47# B1 a_102_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_102_21# A3 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X18 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X20 a_496_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VPWR B1 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.145 ps=1.29 w=1 l=0.15
X22 a_496_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 a_672_297# A2 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 a_600_345# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1 a_788_316# S1 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VPWR A3 a_372_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.164 ps=1.33 w=0.64 l=0.15
X3 a_872_316# a_600_345# a_788_316# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X4 VPWR S0 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 a_1279_413# S0 a_872_316# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND a_788_316# X VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_1060_369# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.16 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_872_316# a_27_47# a_1060_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.138 ps=1.16 w=0.42 l=0.15
X9 a_1281_47# a_27_47# a_872_316# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.072 ps=0.76 w=0.36 l=0.15
X10 a_193_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1064_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0786 pd=0.805 as=0.109 ps=1.36 w=0.42 l=0.15
X12 a_872_316# S1 a_788_316# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.6 as=0.0729 ps=0.81 w=0.54 l=0.15
X13 a_872_316# S0 a_1064_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0786 ps=0.805 w=0.36 l=0.15
X14 X a_788_316# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=1 w=0.65 l=0.15
X15 a_788_316# a_600_345# a_288_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.14 ps=1.6 w=0.54 l=0.15
X16 a_372_413# a_27_47# a_288_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.164 pd=1.33 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VGND A3 a_397_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.0671 ps=0.75 w=0.42 l=0.15
X18 a_600_345# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0819 ps=0.81 w=0.42 l=0.15
X19 a_193_369# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0957 pd=0.965 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 VPWR a_788_316# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.135 ps=1.27 w=1 l=0.15
X21 a_288_47# S0 a_193_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0957 ps=0.965 w=0.42 l=0.15
X22 a_397_47# S0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X23 VGND A0 a_1281_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.066 ps=0.745 w=0.42 l=0.15
X24 a_288_47# a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X25 X a_788_316# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.154 ps=1.34 w=1 l=0.15
X26 VGND S0 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X27 VPWR A0 a_1279_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.105 ps=0.995 w=0.64 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
X0 a_121_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.115 ps=1 w=0.65 l=0.15
X4 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.177 ps=1.36 w=1 l=0.15
X7 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.36 as=0.105 ps=1.21 w=1 l=0.15
X9 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=0.99 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.162 pd=1.15 as=0.111 ps=0.99 w=0.65 l=0.15
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.162 ps=1.15 w=0.65 l=0.15
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.14 ps=1.28 w=1 l=0.15
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.123 ps=1.03 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.119 ps=1.01 w=0.65 l=0.15
X1 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.62 as=0.26 ps=2.52 w=1 l=0.15
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.203 pd=1.27 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.312 ps=1.62 w=1 l=0.15
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X7 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.137 ps=1.07 w=0.65 l=0.15
X8 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.203 ps=1.27 w=0.65 l=0.15
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.21 ps=1.42 w=1 l=0.15
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.138 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_79_21# C1 a_635_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.21 ps=1.42 w=1 l=0.15
X1 VPWR A2 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.17 ps=1.34 w=1 l=0.15
X2 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.08 as=0.133 ps=1.06 w=0.65 l=0.15
X3 a_417_47# A2 a_319_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.02 as=0.111 ps=0.99 w=0.65 l=0.15
X4 a_79_21# A1 a_417_47# VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.12 ps=1.02 w=0.65 l=0.15
X5 a_319_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=0.99 as=0.156 ps=1.13 w=0.65 l=0.15
X6 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.24 pd=1.48 as=0.135 ps=1.27 w=1 l=0.15
X7 a_319_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.185 ps=1.37 w=1 l=0.15
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.156 pd=1.13 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_319_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.34 as=0.24 ps=1.48 w=1 l=0.15
X10 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.14 ps=1.08 w=0.65 l=0.15
X11 a_635_297# B1 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.21 ps=1.42 w=1 l=0.15
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=1.77 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X9 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.385 ps=1.77 w=1 l=0.15
X14 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X21 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X31 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.28 ps=1.62 w=1 l=0.15
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0619 ps=0.715 w=0.42 l=0.15
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0746 pd=0.775 as=0.109 ps=1.36 w=0.42 l=0.15
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.62 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.175 ps=1.26 w=0.65 l=0.15
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0746 ps=0.775 w=0.42 l=0.15
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.172 ps=1.83 w=0.65 l=0.15
X2 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X5 a_326_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.127 ps=1.04 w=0.65 l=0.15
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.635 pd=3.27 as=0.195 ps=1.39 w=1 l=0.15
X7 Y C1 a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=0.393 pd=2.51 as=0.0683 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_223_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 Y A1 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X3 a_223_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X4 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 VGND A2 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_223_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X7 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.123 ps=1.03 w=0.65 l=0.15
X8 VPWR A2 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 a_658_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.201 ps=1.27 w=0.65 l=0.15
X10 VPWR A1 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_223_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_658_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X13 Y a_27_47# a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14 a_223_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15 VPWR A2 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.155 ps=1.31 w=1 l=0.15
X16 VPWR A1 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 a_658_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 VGND B1_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.27 ps=2.13 w=0.65 l=0.15
X19 a_223_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X20 a_658_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X21 VGND A2 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X22 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.27 as=0.091 ps=0.93 w=0.65 l=0.15
X23 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X24 Y A1 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X25 Y a_27_47# a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 Y B1 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_301_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_301_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND B2 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A1 a_735_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_27_297# B2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR A1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_735_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_301_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.176 ps=1.84 w=0.65 l=0.15
X12 VPWR A2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X13 a_383_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X14 a_383_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_735_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X16 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X17 a_301_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X18 a_735_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_109_47# B1 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.165 ps=1.82 w=0.65 l=0.15
X1 Y B2 a_295_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.12 ps=1.24 w=1 l=0.15
X2 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3 a_213_123# B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_295_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12 pd=1.24 as=0.38 ps=1.76 w=1 l=0.15
X5 a_493_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.225 ps=1.45 w=1 l=0.15
X6 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=1.76 as=0.28 ps=2.56 w=1 l=0.15
X7 VGND A2 a_213_123# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X8 a_213_123# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_109_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 Y A1 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_453_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y B1 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.25 ps=1.42 w=0.65 l=0.15
X3 Y A1 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_471_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X6 Y B1 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND A2 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X11 a_453_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_471_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND B2 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_1241_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_27_297# B2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 a_453_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_1241_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_1241_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X21 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VPWR A2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 a_471_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X24 a_471_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_471_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR A1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X28 a_27_297# B1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND A2 a_1241_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 a_471_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_27_297# B1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_1241_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X33 a_471_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 VPWR A1 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X35 a_27_297# B2 a_471_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 a_471_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X38 a_453_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X39 VGND B2 a_453_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 Y A2 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_300_47# B2 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 a_300_47# B1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_300_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_734_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X7 a_28_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y C1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR B1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X11 a_382_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_28_47# B1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_28_47# B2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VGND A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X15 Y B2 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VPWR A1 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND A2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_382_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X19 a_734_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X3 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X5 a_1228_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X6 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X7 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X8 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X10 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X11 VPWR a_1602_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1028_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VGND a_1602_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1028_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X20 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X21 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0441 ps=0.63 w=0.42 l=0.15
X23 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X24 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.223 pd=2.21 as=0.121 ps=1.16 w=0.84 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_1300_47# a_1178_261# a_1228_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X29 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X30 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X31 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.121 pd=1.16 as=0.109 ps=1.36 w=0.42 l=0.15
X32 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X33 VGND SET_B a_1300_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0441 ps=0.63 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.107 ps=0.98 w=0.65 l=0.15
X5 a_277_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
X0 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_475_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_762_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.31 ps=1.62 w=1 l=0.15
X5 a_475_47# B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X6 VGND A2 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X10 a_80_21# A2 a_762_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_80_21# B1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X12 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15 ps=1.3 w=1 l=0.15
X13 a_475_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.117 ps=1.01 w=0.65 l=0.15
X14 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 VPWR A1 a_934_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X16 a_934_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 VPWR B1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=1.62 as=0.14 ps=1.28 w=1 l=0.15
X18 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND A1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.117 ps=1.01 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_467_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_109_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VPWR A a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_555_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_197_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_197_297# B a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 Y a_27_47# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y a_27_47# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X16 a_555_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_555_297# B a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_197_297# B a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 a_555_297# B a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A a_197_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X23 a_197_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X25 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 a_676_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.213 ps=1.42 w=1 l=0.15
X1 a_512_47# B1 a_409_47# VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.119 ps=1.01 w=0.65 l=0.15
X2 a_306_47# D1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.198 ps=1.91 w=0.65 l=0.15
X3 VGND A2 a_512_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.198 ps=1.26 w=0.65 l=0.15
X4 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.218 ps=1.43 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.305 ps=1.61 w=1 l=0.15
X6 VPWR A1 a_676_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X7 a_512_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_409_47# C1 a_306_47# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.119 ps=1.01 w=0.65 l=0.15
X9 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.382 pd=1.76 as=0.26 ps=2.52 w=1 l=0.15
X10 a_79_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=1.43 as=0.382 ps=1.76 w=1 l=0.15
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.148 ps=1.34 w=0.42 l=0.15
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.102 ps=0.99 w=0.42 l=0.15
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 Y a_61_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.183 ps=1.24 w=0.65 l=0.15
X1 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_217_297# a_61_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_479_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X4 a_217_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5 Y a_61_47# a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VPWR A1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 a_61_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X8 VGND A2 a_637_47# VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND a_61_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y A1 a_479_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0683 ps=0.86 w=0.65 l=0.15
X11 VGND B1_N a_61_47# VNB sky130_fd_pr__nfet_01v8 ad=0.183 pd=1.24 as=0.126 ps=1.44 w=0.42 l=0.15
X12 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X13 a_637_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_484_297# B2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND B2 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_96_21# B1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X8 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_484_297# B1 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_484_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A2 a_918_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_96_21# B2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 a_96_21# B1 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_484_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR A1 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_96_21# A1 a_918_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VPWR A2 a_484_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X18 a_566_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X19 a_918_47# A1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_566_47# B1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 a_918_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X22 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.0829 ps=0.905 w=0.65 l=0.15
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.101 ps=0.96 w=0.65 l=0.15
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.125 ps=1.25 w=1 l=0.15
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.214 ps=1.96 w=0.65 l=0.15
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.25 as=0.385 ps=2.77 w=1 l=0.15
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.56 as=0.18 ps=1.36 w=1 l=0.15
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.135 ps=1.27 w=1 l=0.15
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0.0829 pd=0.905 as=0.185 ps=1.22 w=0.65 l=0.15
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.275 ps=1.5 w=0.65 l=0.15
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=1.56 w=1 l=0.15
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.22 as=0.117 ps=1.01 w=0.65 l=0.15
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
X0 a_398_413# a_206_93# a_316_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR a_316_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_316_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X3 X a_316_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X4 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.32 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND a_27_410# a_316_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X7 VGND A a_316_413# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND a_316_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_566_297# B a_494_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0598 pd=0.705 as=0.0441 ps=0.63 w=0.42 l=0.15
X10 a_206_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0619 ps=0.715 w=0.42 l=0.15
X11 a_316_413# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_206_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.123 ps=1.32 w=0.42 l=0.15
X13 a_494_297# a_27_410# a_398_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.122 ps=1.33 w=0.42 l=0.15
X14 a_316_413# a_206_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X15 VPWR A a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0598 ps=0.705 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.0683 ps=0.745 w=0.42 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.09 as=0.0696 ps=0.765 w=0.42 l=0.15
X8 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X10 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0683 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X11 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0767 ps=0.785 w=0.42 l=0.15
X12 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.09 w=0.64 l=0.15
X13 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.08 as=0.179 ps=1.26 w=0.75 l=0.15
X14 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.08 w=0.42 l=0.15
X18 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X19 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X20 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X21 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X22 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X23 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X25 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X6 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.123 ps=1.17 w=0.84 l=0.15
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 a_39_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR A1 a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X4 a_125_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X5 a_125_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_125_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_1163_47# B1 a_125_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_39_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_1163_47# B1 a_125_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VGND A3 a_125_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND A1 a_125_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND A3 a_125_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_39_297# A2 a_461_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A1 a_125_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_125_47# B1 a_1163_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X17 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 a_125_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X19 VGND A2 a_125_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_125_47# B1 a_1163_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VGND A2 a_125_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y C1 a_1163_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 Y C1 a_1163_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 a_461_297# A2 a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y A3 a_461_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y A3 a_461_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_125_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 VPWR A1 a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X31 a_461_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_461_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X33 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 a_125_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 a_1163_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 a_1163_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X37 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 a_39_297# A2 a_461_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 a_461_297# A2 a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.91 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.192 ps=1.38 w=1 l=0.15
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.192 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125 ps=1.03 w=0.65 l=0.15
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_108_21# B1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 a_346_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X2 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.263 ps=2.11 w=0.65 l=0.15
X3 a_108_21# A3 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4 a_430_297# A2 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.175 ps=1.35 w=1 l=0.15
X6 a_346_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.405 ps=2.81 w=1 l=0.15
X9 VPWR B1 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.213 ps=1.42 w=1 l=0.15
X10 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.114 ps=1 w=0.65 l=0.15
X11 a_346_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 Y A1 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.377 ps=1.75 w=1 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.305 ps=1.61 w=1 l=0.15
X3 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.335 ps=1.67 w=1 l=0.15
X4 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.138 ps=1.27 w=1 l=0.15
X5 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.377 pd=1.75 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_478_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_478_47# A2 a_730_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VGND A3 a_730_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12 ps=1.02 w=0.65 l=0.15
X10 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_730_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.02 as=0.205 ps=1.93 w=0.65 l=0.15
X16 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.15 ps=1.3 w=1 l=0.15
X18 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X19 a_730_47# A2 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_82_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 a_646_47# B2 a_82_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_574_369# a_313_47# a_82_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0976 pd=0.945 as=0.166 ps=1.8 w=0.64 l=0.15
X3 a_574_369# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4 VGND a_82_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR B2 a_574_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0976 ps=0.945 w=0.64 l=0.15
X6 X a_82_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X7 X a_82_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X8 a_313_47# A2_N a_313_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17 pd=1.81 as=0.0672 ps=0.85 w=0.64 l=0.15
X9 a_313_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X10 a_313_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.186 ps=1.43 w=0.64 l=0.15
X11 VGND A2_N a_313_47# VNB sky130_fd_pr__nfet_01v8 ad=0.142 pd=1.1 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_82_21# a_313_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.142 ps=1.1 w=0.42 l=0.15
X13 VGND B1 a_646_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.159 ps=1.14 w=0.65 l=0.15
X3 a_1139_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.245 pd=1.49 as=0.135 ps=1.27 w=1 l=0.15
X4 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_109_297# B1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_1139_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_109_297# B1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_1139_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 Y C1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_1139_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.159 pd=1.14 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X32 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y C1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.245 ps=1.49 w=1 l=0.15
X35 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X38 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X39 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.131 ps=1.05 w=0.64 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.41 as=0.135 ps=1.27 w=1 l=0.15
X3 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.05 as=0.229 ps=1.36 w=0.64 l=0.15
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0578 ps=0.695 w=0.42 l=0.15
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.36 as=0.178 ps=1.41 w=0.64 l=0.15
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.173 pd=1.25 as=0.0683 ps=0.745 w=0.42 l=0.15
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.173 ps=1.25 w=0.42 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
X0 VPWR A a_304_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X1 a_304_297# B a_220_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND C a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X3 a_220_297# C a_114_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X4 a_32_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_32_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X11 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X13 a_114_297# D a_32_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X14 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
X0 VGND B1 a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_741_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.101 ps=0.96 w=0.65 l=0.15
X2 a_84_21# A1 a_741_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0747 ps=0.88 w=0.65 l=0.15
X3 VGND A2 a_901_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR A2 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_483_297# B1 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.185 ps=1.87 w=0.65 l=0.15
X8 a_84_21# B1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.265 pd=1.47 as=0.091 ps=0.93 w=0.65 l=0.15
X10 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_483_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=2.79 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR A1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X14 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.285 ps=2.57 w=1 l=0.15
X15 a_84_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.265 ps=1.47 w=0.65 l=0.15
X16 a_483_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X18 a_901_47# A1 a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
X0 VPWR A a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_218_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.156 ps=1.16 w=0.42 l=0.15
X2 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.156 pd=1.16 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_300_297# a_27_53# a_218_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X4 X a_218_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X5 VPWR a_218_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_218_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND a_218_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_218_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X1 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.194 pd=1.95 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VGND B a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y a_27_93# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_229_47# a_27_93# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.147 ps=1.34 w=1 l=0.15
X6 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.165 ps=1.33 w=1 l=0.15
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X8 a_229_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0943 pd=0.94 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0943 ps=0.94 w=0.65 l=0.15
X4 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0959 ps=0.945 w=0.65 l=0.15
X7 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.147 ps=1.29 w=1 l=0.15
X10 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0959 ps=0.945 w=0.65 l=0.15
X18 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X20 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.237 pd=1.48 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.237 ps=1.48 w=1 l=0.15
X28 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X32 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X33 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X34 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.0878 ps=0.92 w=0.65 l=0.15
X37 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X39 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.63 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.14 ps=1.28 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.305 ps=2.61 w=1 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.139 ps=1.5 w=0.42 l=0.15
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
X0 Y a_27_47# a_432_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y a_27_47# a_432_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_850_47# a_193_47# a_432_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND D a_1266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.555 ps=2.11 w=1 l=0.15
X8 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X10 a_432_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_432_47# a_193_47# a_850_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_432_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_432_47# a_193_47# a_850_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR a_193_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.555 pd=2.11 as=0.135 ps=1.27 w=1 l=0.15
X16 a_193_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.495 pd=2.99 as=0.135 ps=1.27 w=1 l=0.15
X17 Y a_193_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_193_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.322 pd=2.29 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_850_47# C a_1266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.189 ps=1.88 w=0.65 l=0.15
X22 a_850_47# a_193_47# a_432_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 a_850_47# C a_1266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VGND D a_1266_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 VPWR a_193_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_1266_47# C a_850_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 Y a_193_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_1266_47# C a_850_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 a_1266_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X32 a_1266_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X34 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X35 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_294_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0662 pd=0.735 as=0.0986 ps=0.98 w=0.42 l=0.15
X1 VPWR A2_N a_295_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.227 pd=1.35 as=0.173 ps=1.4 w=0.64 l=0.15
X2 VPWR B1 a_665_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0986 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.185 ps=1.87 w=0.65 l=0.15
X5 a_581_47# a_295_369# a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X7 a_665_369# B2 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0928 ps=0.93 w=0.64 l=0.15
X8 VGND B2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_295_369# A2_N a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0662 ps=0.735 w=0.42 l=0.15
X10 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.285 ps=2.57 w=1 l=0.15
X11 a_84_21# a_295_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0928 pd=0.93 as=0.227 ps=1.35 w=0.64 l=0.15
X12 a_295_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.4 as=0.154 ps=1.34 w=0.64 l=0.15
X13 a_581_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
X0 VGND A a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VPWR A a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0598 ps=0.705 w=0.42 l=0.15
X2 a_393_413# a_205_93# a_311_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.122 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.32 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_311_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.148 ps=1.34 w=1 l=0.15
X6 VGND a_27_410# a_311_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0598 ps=0.705 w=0.42 l=0.15
X7 a_561_297# B a_489_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0598 pd=0.705 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 a_205_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0619 ps=0.715 w=0.42 l=0.15
X9 a_205_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.123 ps=1.32 w=0.42 l=0.15
X10 a_489_297# a_27_410# a_393_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.122 ps=1.33 w=0.42 l=0.15
X11 a_311_413# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_311_413# a_205_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0598 pd=0.705 as=0.109 ps=1.36 w=0.42 l=0.15
X13 X a_311_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.102 ps=0.99 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 a_27_47# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.368 pd=1.74 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.231 pd=2.01 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3 VPWR A1 a_373_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X4 a_182_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.165 ps=1.82 w=0.65 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.195 ps=1.39 w=1 l=0.15
X6 a_182_47# B1 a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X8 a_373_297# A2 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.368 ps=1.74 w=1 l=0.15
X9 a_110_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X10 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11 VGND A1 a_182_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
X0 a_429_297# A2 a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND A2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.08 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_345_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.14 ps=1.08 w=0.65 l=0.15
X5 a_345_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=1.61 w=1 l=0.15
X6 a_629_297# B2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR B1 a_629_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.19 ps=1.38 w=1 l=0.15
X8 a_79_21# B2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_345_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.123 ps=1.03 w=0.65 l=0.15
X10 a_79_21# A3 a_429_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X12 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_345_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.198 ps=1.26 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 Y A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.109 ps=0.985 w=0.65 l=0.15
X4 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_949_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y C1 a_949_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.15 ps=1.3 w=1 l=0.15
X10 a_781_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_27_297# B1 a_781_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 Y A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_781_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_1301_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.15 ps=1.3 w=1 l=0.15
X16 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 Y C1 a_781_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.14 ps=1.28 w=1 l=0.15
X18 a_109_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_109_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 a_109_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X27 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X28 a_27_297# B1 a_1301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X29 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0894 ps=0.925 w=0.65 l=0.15
X30 a_109_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_465_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_204_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0699 pd=0.865 as=0.106 ps=0.975 w=0.65 l=0.15
X4 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.91 as=0.0991 ps=0.955 w=0.65 l=0.15
X5 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X6 Y B1 a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0699 ps=0.865 w=0.65 l=0.15
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.153 ps=1.3 w=1 l=0.15
X8 a_109_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1 a_277_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2 a_79_21# B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3 a_277_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_361_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_277_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.127 ps=1.04 w=0.65 l=0.15
X9 a_79_21# A1 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.107 ps=0.98 w=0.65 l=0.15
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.115 ps=1 w=0.65 l=0.15
X1 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.0926 ps=0.935 w=0.65 l=0.15
X2 VPWR A1 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.105 ps=1.21 w=1 l=0.15
X3 a_307_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.233 ps=1.47 w=1 l=0.15
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.233 pd=1.47 as=0.112 ps=1.23 w=1 l=0.15
X6 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.112 pd=1.23 as=0.26 ps=2.52 w=1 l=0.15
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 Y A3 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_449_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 Y A3 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y B1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_449_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.263 ps=2.57 w=1 l=0.15
X8 Y B1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_31_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_27_297# A2 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.261 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND A1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_31_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 a_31_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_31_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_449_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X20 VGND A2 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VGND A2 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 VGND A3 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.223 pd=1.34 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 a_31_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.223 ps=1.34 w=0.65 l=0.15
X25 a_27_297# A2 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND A3 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 a_31_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
X28 a_449_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_31_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_31_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
X0 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X17 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X23 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X5 a_277_47# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_193_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_361_47# A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VGND A3 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X15 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X16 a_277_47# A1 a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_445_47# A2 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.5 pd=3 as=0.135 ps=1.27 w=1 l=0.15
X22 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X23 a_277_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
X0 VPWR a_193_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND D a_781_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y a_193_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X6 a_591_47# C a_781_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 a_781_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_781_47# C a_591_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR B_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X10 a_193_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.197 pd=1.78 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 Y a_193_47# a_341_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_591_47# a_27_47# a_341_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X14 a_341_47# a_193_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_341_47# a_27_47# a_591_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X17 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 a_193_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.197 pd=1.78 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VGND B_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 a_79_21# A1 a_348_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.133 ps=1.06 w=0.65 l=0.15
X1 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.26 as=0.091 ps=0.93 w=0.65 l=0.15
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_79_21# C1 a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X5 VPWR A2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X6 a_299_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.195 ps=1.39 w=1 l=0.15
X7 a_585_297# B1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_348_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.2 ps=1.26 w=0.65 l=0.15
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.115 ps=1 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X4 a_215_297# a_109_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.165 ps=1.82 w=0.65 l=0.15
X5 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X6 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X8 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_109_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X10 VPWR A a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X11 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_487_297# B a_403_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_403_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X14 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X16 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_297_297# a_109_93# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.198 ps=1.26 w=0.65 l=0.15
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.393 pd=1.78 as=0.135 ps=1.27 w=1 l=0.15
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.393 ps=1.78 w=1 l=0.15
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 VPWR B1 a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X1 a_484_47# B1 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_566_297# B2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X8 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_96_21# B2 a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A1 a_918_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X11 a_484_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_566_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X13 a_484_47# B2 a_96_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_96_21# A2 a_918_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_918_297# A2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 a_484_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_918_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X18 a_96_21# B1 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X19 VGND A2 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_96_21# B2 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VGND A1 a_484_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X22 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X23 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
X0 VGND A2 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 VPWR A1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 a_37_297# B1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4 a_485_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_292_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X7 VPWR A2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_485_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X11 a_37_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 Y A1 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X13 Y C1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X14 a_292_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X15 a_292_297# B1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
X0 VGND B1_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VGND A2 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.106 ps=0.975 w=0.65 l=0.15
X2 a_478_47# a_27_93# a_174_21# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_478_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X5 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X6 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X7 VPWR A1 a_574_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X8 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR B1_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X10 a_574_297# A2 a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X11 a_174_21# a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.395 ps=1.79 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14 ps=1.28 w=1 l=0.15
X1 VGND A3 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X2 a_309_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0715 pd=0.87 as=0.153 ps=1.12 w=0.65 l=0.15
X3 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.153 pd=1.12 as=0.0747 ps=0.88 w=0.65 l=0.15
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X5 a_383_47# A2 a_309_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0715 ps=0.87 w=0.65 l=0.15
X6 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X7 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 VGND A4 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_321_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.123 ps=1.03 w=0.65 l=0.15
X2 a_103_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_103_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.425 ps=2.85 w=1 l=0.15
X4 VGND a_103_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.247 ps=2.06 w=0.65 l=0.15
X5 VGND A2 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X6 a_321_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.127 ps=1.04 w=0.65 l=0.15
X7 a_511_297# A3 a_393_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.22 ps=1.44 w=1 l=0.15
X8 a_619_297# A2 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 a_321_47# B1 a_103_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_393_297# A4 a_103_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.26 ps=1.52 w=1 l=0.15
X11 VPWR A1 a_619_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
X0 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.117 ps=1.01 w=0.65 l=0.15
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=1.82 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.175 ps=1.35 w=1 l=0.15
X4 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.41 ps=1.82 w=1 l=0.15
X10 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.18 ps=1.36 w=1 l=0.15
X11 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X13 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0975 ps=0.95 w=0.65 l=0.15
X14 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
X0 VGND B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X2 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VGND B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_215_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.254 pd=2.08 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_215_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X17 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
X0 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X3 a_91_199# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_245_297# B a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_91_199# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.146 ps=1.34 w=0.42 l=0.15
X7 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
X0 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.36 as=0.14 ps=1.28 w=1 l=0.15
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138 ps=1.08 w=0.65 l=0.15
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND B a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.08 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X8 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.177 ps=1.36 w=1 l=0.15
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
X0 a_176_21# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 VGND D_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.5 as=0.135 ps=1.27 w=1 l=0.15
X5 a_555_297# C a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_176_21# a_27_53# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.169 ps=1.5 w=1 l=0.15
X8 a_387_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.168 ps=1.5 w=0.42 l=0.15
X9 a_483_297# B a_387_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X11 VGND a_27_53# a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 VPWR D_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.169 pd=1.5 as=0.109 ps=1.36 w=0.42 l=0.15
X13 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1 ps=0.985 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.14 ps=1.28 w=1 l=0.15
X1 a_235_47# C1 a_163_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.0683 ps=0.86 w=0.65 l=0.15
X2 a_343_47# B1 a_235_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.05 as=0.127 ps=1.04 w=0.65 l=0.15
X3 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.203 pd=1.4 as=0.195 ps=1.39 w=1 l=0.15
X4 a_454_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.203 ps=1.4 w=1 l=0.15
X5 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6 VPWR A1 a_454_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.195 ps=1.39 w=1 l=0.15
X7 a_163_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X8 VGND A2 a_343_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.132 ps=1.05 w=0.65 l=0.15
X9 a_343_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.127 ps=1.04 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
X0 VPWR A1 a_485_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_485_297# a_297_93# a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 a_297_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.108 ps=1.01 w=0.42 l=0.15
X3 a_581_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.01 as=0.091 ps=0.93 w=0.65 l=0.15
X5 a_79_21# a_297_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VGND A2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.51 as=0.14 ps=1.28 w=1 l=0.15
X8 a_297_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.182 ps=1.51 w=0.42 l=0.15
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X10 a_485_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_33_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.182 ps=1.86 w=0.65 l=0.15
X4 Y a_33_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7 Y a_33_297# a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VGND A2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X11 a_225_47# a_33_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_225_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VPWR A1 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 a_561_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR B1_N a_33_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X20 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y A2 a_561_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X24 a_561_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 VPWR a_33_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 a_33_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND A1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VGND A2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_33_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_797_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_797_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y B2 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR B1 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_33_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VGND A1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_33_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_33_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_33_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_797_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.16 ps=1.32 w=1 l=0.15
X17 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR B1 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 a_33_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 a_797_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.135 ps=1.27 w=1 l=0.15
X24 Y B2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 Y B2 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 Y B1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.104 ps=0.97 w=0.65 l=0.15
X27 Y B2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 Y B1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 a_33_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.229 ps=1.75 w=1 l=0.15
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0767 ps=0.785 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.75 as=0.0609 ps=0.71 w=0.42 l=0.15
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0894 ps=0.925 w=0.65 l=0.15
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.119 ps=1.01 w=0.65 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 Y A1 a_194_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_194_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X2 Y C1 a_376_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.35 w=1 l=0.15
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.112 ps=0.995 w=0.65 l=0.15
X5 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.115 ps=1 w=0.65 l=0.15
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X7 a_376_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.165 ps=1.33 w=1 l=0.15
X8 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
X0 Y C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X6 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X10 a_281_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X3 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 Y A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X17 a_803_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X30 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X31 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
X0 Y A a_150_67# VNB sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.67 as=0.066 ps=0.79 w=0.55 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0.14 ps=1.28 w=1 l=0.25
X2 a_150_67# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.79 as=0.157 ps=1.67 w=0.55 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
.ends

.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 X a_91_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X1 a_91_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X2 a_360_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.137 ps=1.07 w=0.65 l=0.15
X3 VPWR B1 a_91_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.138 ps=1.27 w=1 l=0.15
X4 a_360_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.312 ps=1.62 w=1 l=0.15
X5 VGND A2 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0.137 pd=1.07 as=0.114 ps=1 w=0.65 l=0.15
X6 a_360_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.203 ps=1.27 w=0.65 l=0.15
X7 VPWR a_91_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.62 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND a_91_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.203 pd=1.27 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 X a_91_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.208 ps=1.94 w=0.65 l=0.15
X10 a_677_47# B1 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.119 ps=1.01 w=0.65 l=0.15
X11 a_460_297# A2 a_360_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.175 ps=1.35 w=1 l=0.15
X12 a_91_21# C1 a_677_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X13 a_91_21# A3 a_460_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.21 ps=1.42 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_471_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_471_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_471_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X5 a_471_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_471_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_1241_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X10 a_27_47# B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR B1 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND A2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_553_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X14 a_27_47# B2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VGND A2 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VGND A1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X19 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_1241_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR B1 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A1 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 Y B2 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_1241_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X26 a_553_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_471_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 Y A2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_553_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_27_47# B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 VGND A1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X32 Y B2 a_553_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_1241_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 a_27_47# B1 a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 a_553_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X36 Y A2 a_1241_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X38 a_471_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 a_471_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 a_298_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VGND A1 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3 a_664_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.14 ps=1.28 w=1 l=0.15
X4 VGND A2 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 a_298_47# B1 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.176 ps=1.84 w=0.65 l=0.15
X7 a_497_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X8 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.224 ps=1.99 w=0.65 l=0.15
X9 a_497_47# B1 a_298_47# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 Y A2 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.295 ps=2.59 w=1 l=0.15
X12 a_27_47# C1 a_298_47# VNB sky130_fd_pr__nfet_01v8 ad=0.192 pd=1.89 as=0.091 ps=0.93 w=0.65 l=0.15
X13 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X14 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X16 a_497_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.091 ps=0.93 w=0.65 l=0.15
X17 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X18 VPWR A1 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 a_664_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_27_47# a_415_21# a_193_297# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VPWR A2_N a_415_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_415_21# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X3 a_415_21# A2_N a_717_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_193_297# a_415_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR a_193_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_193_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_109_297# B2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_193_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_717_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_717_47# A2_N a_415_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_193_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_27_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_27_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VGND a_193_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VGND A1_N a_717_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND a_193_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 VGND B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_193_297# a_415_21# a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VPWR a_193_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR a_415_21# a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X23 X a_193_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A1_N a_415_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 a_415_21# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 VGND B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_475_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR A1 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X9 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.27 pd=1.48 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X12 a_475_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 Y A2 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X14 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.27 ps=1.48 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 a_236_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.163 ps=1.17 w=0.65 l=0.15
X1 a_428_47# A2 a_336_47# VNB sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.08 as=0.101 ps=0.96 w=0.65 l=0.15
X2 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.37 pd=2.74 as=0.213 ps=1.42 w=1 l=0.15
X3 Y A1 a_428_47# VNB sky130_fd_pr__nfet_01v8 ad=0.241 pd=2.04 as=0.138 ps=1.08 w=0.65 l=0.15
X4 a_336_47# A3 a_236_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X5 VPWR A4 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.213 ps=1.42 w=1 l=0.15
X6 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.26 ps=2.52 w=1 l=0.15
X7 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.205 ps=1.41 w=1 l=0.15
X8 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.155 ps=1.31 w=1 l=0.15
X9 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.163 pd=1.17 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_27_47# B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_109_47# A2 a_717_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_717_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X3 VGND A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_277_297# B2 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_47# B2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_277_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 a_277_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_277_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR C1 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 a_27_47# C1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_27_47# B2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VGND A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_277_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_277_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X23 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A1 a_717_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_109_47# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 a_717_297# A2 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_109_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X15 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
X0 a_27_47# C a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_47# C a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_445_47# B a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_445_47# B a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 Y A a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X14 Y A a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_803_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X17 a_803_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_445_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_803_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X24 a_445_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 a_803_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X30 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X31 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.247 ps=2.06 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.43 ps=2.86 w=1 l=0.15
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_109_47# A2_N a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 a_397_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B2 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A2_N a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.283 pd=1.52 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_397_297# a_109_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.34 ps=2.68 w=1 l=0.15
X5 a_481_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.283 ps=1.52 w=0.65 l=0.15
X7 VGND B1 a_481_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_109_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
X0 VPWR a_193_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1 a_297_47# a_27_413# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.104 ps=1 w=0.65 l=0.15
X4 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.143 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=1 as=0.0619 ps=0.715 w=0.42 l=0.15
X7 VGND a_193_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0991 ps=0.955 w=0.65 l=0.15
X8 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X9 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X10 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.143 ps=1.33 w=1 l=0.15
X11 a_193_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.715 as=0.0735 ps=0.77 w=0.42 l=0.15
X13 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
X0 a_408_47# B a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_408_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y a_27_47# a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176 pd=1.39 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND C a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_218_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.12 ps=1.04 w=0.65 l=0.15
X7 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_218_47# B a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.176 ps=1.39 w=1 l=0.15
X12 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.04 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 VGND A2 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.114 ps=1 w=0.65 l=0.15
X1 a_496_297# A4 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.36 as=0.303 ps=1.61 w=1 l=0.15
X2 a_393_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.115 ps=1 w=0.65 l=0.15
X3 VPWR A1 a_697_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=2.82 as=0.175 ps=1.35 w=1 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.303 pd=1.61 as=0.305 ps=1.61 w=1 l=0.15
X7 VGND A4 a_393_47# VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.119 ps=1.01 w=0.65 l=0.15
X8 a_697_297# A2 a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.175 ps=1.35 w=1 l=0.15
X9 a_393_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.266 pd=2.12 as=0.114 ps=1 w=0.65 l=0.15
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_393_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.208 ps=1.94 w=0.65 l=0.15
X12 a_597_297# A3 a_496_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.177 ps=1.36 w=1 l=0.15
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_1224_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VPWR A1 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.183 ps=1.37 w=1 l=0.15
X2 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_806_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.205 ps=1.28 w=0.65 l=0.15
X8 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.205 pd=1.28 as=0.14 ps=1.08 w=0.65 l=0.15
X10 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_806_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A3 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 Y A3 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X19 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.119 ps=1.01 w=0.65 l=0.15
X22 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0926 ps=0.935 w=0.65 l=0.15
X24 a_806_297# A2 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X25 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.142 ps=1.28 w=1 l=0.15
X28 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.08 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 a_1224_297# A2 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_1224_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.183 pd=1.37 as=0.135 ps=1.27 w=1 l=0.15
X32 a_806_297# A2 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 VPWR A1 a_1224_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X37 a_1224_297# A2 a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X39 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2 a_80_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.365 ps=1.73 w=1 l=0.15
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4 VPWR C1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.14 ps=1.28 w=1 l=0.15
X5 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X6 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X7 a_674_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X8 a_386_47# D1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X9 VPWR A1 a_674_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.195 ps=1.39 w=1 l=0.15
X10 a_566_47# B1 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X11 VGND A2 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X12 a_566_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.127 ps=1.04 w=0.65 l=0.15
X13 a_458_47# C1 a_386_47# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.0683 ps=0.86 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_641_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_109_297# B1 a_641_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X5 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.17 w=0.65 l=0.15
X11 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X12 a_641_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0975 ps=0.95 w=0.65 l=0.15
X15 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 Y C1 a_641_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=1.52 w=1 l=0.15
X18 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X19 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 Y B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VGND a_751_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_751_21# A2_N a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_1139_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VPWR B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND A2_N a_751_21# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_27_297# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A1_N a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y a_751_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_1139_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 a_27_297# a_751_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X13 Y a_751_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR A1_N a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 a_751_21# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X16 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_27_297# a_751_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VGND B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 Y B2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X20 Y a_751_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_1139_297# A2_N a_751_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X22 a_751_21# A2_N a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VGND A1_N a_751_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 VGND A1_N a_751_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 a_109_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VGND A2_N a_751_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 a_109_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 VPWR B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_109_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 Y a_751_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X32 a_27_297# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 a_751_21# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X34 a_751_21# A2_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X36 a_1139_297# A2_N a_751_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 a_109_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X38 VGND a_751_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 a_751_21# A2_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt fpga_wrapper VGND VPWR clk_mosi clk_sys cs pwmA pwmB pwmC ready rstb spi_mosi
XFILLER_0_20_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18869_ _10718_ _10716_ VGND VGND VPWR VPWR _10844_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20900_ _12681_ _11788_ _12683_ VGND VGND VPWR VPWR _12748_ sky130_fd_sc_hd__mux2_1
X_21880_ _01441_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__inv_2
X_20831_ _12198_ _12200_ _12203_ VGND VGND VPWR VPWR _12680_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23550_ _02941_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__clkbuf_1
X_20762_ net300 net292 VGND VGND VPWR VPWR _12611_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22501_ net111 _02020_ _02018_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__o21a_1
X_23481_ _02905_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20693_ _12539_ _12541_ _12535_ VGND VGND VPWR VPWR _12542_ sky130_fd_sc_hd__a21o_1
X_25220_ _04565_ _04566_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__and2b_1
XFILLER_0_175_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22432_ _01885_ _01941_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25151_ _04437_ _04439_ _04371_ _03687_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__o211a_1
XFILLER_0_162_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22363_ net125 net120 _01778_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24102_ _03458_ _03459_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__xnor2_1
X_21314_ _13138_ _13136_ _13139_ VGND VGND VPWR VPWR _13156_ sky130_fd_sc_hd__a21bo_1
X_25082_ _04429_ _04430_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22294_ net91 _01848_ _01851_ net95 _01853_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24033_ _03388_ _03389_ _03390_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21245_ _12606_ _12578_ _13086_ VGND VGND VPWR VPWR _13089_ sky130_fd_sc_hd__or3_1
XFILLER_0_103_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21176_ net252 _12982_ VGND VGND VPWR VPWR _13020_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20127_ top0.cordic0.slte0.opA\[16\] VGND VGND VPWR VPWR _11983_ sky130_fd_sc_hd__inv_2
X_25984_ top0.pid_q.out\[6\] _12032_ _05014_ spi0.data_packed\[54\] VGND VGND VPWR
+ VPWR _05188_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_0_clk_sys clknet_3_2__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_0_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_24935_ _04187_ _04193_ _04185_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__a21bo_1
X_20058_ _11918_ _11920_ VGND VGND VPWR VPWR _11921_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24866_ _03765_ _03908_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26605_ clknet_leaf_67_clk_sys _00228_ net660 VGND VGND VPWR VPWR top0.pid_q.curr_int\[15\]
+ sky130_fd_sc_hd__dfrtp_2
X_23817_ _03170_ _03171_ _03174_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__a21o_1
XFILLER_0_169_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24797_ _04149_ _04147_ _04032_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14550_ net44 _06268_ VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__and2_1
XFILLER_0_184_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26536_ clknet_leaf_60_clk_sys _00159_ net652 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_23748_ _03066_ _03067_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__nor2_4
XFILLER_0_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13501_ _05676_ _05713_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14481_ _06687_ _06674_ _06672_ VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__mux2_1
X_26467_ clknet_leaf_18_clk_sys net575 net612 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23679_ net572 top0.matmul0.matmul_stage_inst.d\[4\] top0.matmul0.matmul_stage_inst.c\[4\]
+ net556 VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__a22o_2
XFILLER_0_165_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16220_ _08220_ VGND VGND VPWR VPWR _08312_ sky130_fd_sc_hd__clkbuf_4
X_25418_ _04663_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__inv_2
X_13432_ _05582_ _05592_ _05644_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__o21a_1
XFILLER_0_153_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26398_ clknet_leaf_79_clk_sys _00039_ net588 VGND VGND VPWR VPWR top0.kpd\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16151_ top0.pid_q.curr_int\[6\] VGND VGND VPWR VPWR _08243_ sky130_fd_sc_hd__inv_2
X_25349_ _04692_ _04693_ _04518_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__a21oi_2
X_13363_ _05571_ _05572_ _05575_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15102_ _07197_ _07200_ VGND VGND VPWR VPWR _07201_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_107_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16082_ _08115_ _08117_ _08113_ VGND VGND VPWR VPWR _08175_ sky130_fd_sc_hd__a21bo_1
X_13294_ _05502_ _05506_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27019_ clknet_leaf_17_clk_sys _00636_ net611 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_15033_ top0.pid_d.prev_int\[3\] _07140_ _07144_ top0.pid_d.curr_int\[3\] VGND VGND
+ VPWR VPWR _00120_ sky130_fd_sc_hd__a22o_1
X_19910_ _11783_ VGND VGND VPWR VPWR _11784_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19841_ _11702_ _11700_ VGND VGND VPWR VPWR _11719_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16984_ top0.currT_r\[11\] _09033_ VGND VGND VPWR VPWR _09039_ sky130_fd_sc_hd__or2_1
X_19772_ _11573_ VGND VGND VPWR VPWR _11654_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15935_ _08028_ _08029_ VGND VGND VPWR VPWR _08030_ sky130_fd_sc_hd__xnor2_1
X_18723_ _10694_ _10699_ VGND VGND VPWR VPWR _10700_ sky130_fd_sc_hd__xor2_1
X_18654_ net331 _10545_ VGND VGND VPWR VPWR _10632_ sky130_fd_sc_hd__xor2_4
XFILLER_0_188_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15866_ _07944_ _07961_ VGND VGND VPWR VPWR _07962_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_188_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14817_ _05666_ _07016_ _06867_ net26 VGND VGND VPWR VPWR _07017_ sky130_fd_sc_hd__o211a_1
X_17605_ _09574_ _09579_ _09591_ VGND VGND VPWR VPWR _09592_ sky130_fd_sc_hd__a21oi_1
X_18585_ _10103_ _10563_ VGND VGND VPWR VPWR _10564_ sky130_fd_sc_hd__xnor2_1
X_15797_ _07892_ _07893_ VGND VGND VPWR VPWR _07894_ sky130_fd_sc_hd__and2b_1
XFILLER_0_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17536_ net340 net425 VGND VGND VPWR VPWR _09523_ sky130_fd_sc_hd__nand2_1
X_14748_ _06896_ _06916_ _06917_ VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_86_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17467_ _09376_ _09379_ VGND VGND VPWR VPWR _09454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14679_ _06217_ _05626_ _06882_ _06106_ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__o22a_1
XFILLER_0_157_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16418_ _08495_ _08506_ VGND VGND VPWR VPWR _08507_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19206_ _11154_ _11145_ _11155_ VGND VGND VPWR VPWR _11156_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17398_ _09379_ _09384_ VGND VGND VPWR VPWR _09385_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19137_ top0.kid\[3\] _11098_ _11100_ top0.kpd\[3\] VGND VGND VPWR VPWR _11104_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16349_ _08436_ _08438_ VGND VGND VPWR VPWR _08439_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19068_ _11017_ _11021_ VGND VGND VPWR VPWR _11040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18019_ _09941_ _09946_ _09939_ VGND VGND VPWR VPWR _10004_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21030_ _12749_ _12746_ _12876_ VGND VGND VPWR VPWR _12877_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_11_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout105 net106 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_8
Xfanout116 net1031 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_4
Xfanout127 net128 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout138 net140 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_2
XFILLER_0_201_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout149 top0.cordic0.vec\[1\]\[3\] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_4
X_22981_ top0.svm0.counter\[8\] _02483_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__nor2_1
X_24720_ _02994_ _02996_ _03150_ _03151_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__o22a_1
X_21932_ net151 net137 VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24651_ _04001_ _04002_ _04003_ _04004_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__a211o_1
XFILLER_0_96_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21863_ _01379_ _01423_ _01424_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_171_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23602_ net1024 _09296_ net559 VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20814_ _12579_ _12662_ _12546_ VGND VGND VPWR VPWR _12663_ sky130_fd_sc_hd__a21o_1
X_24582_ _03824_ _03935_ _03936_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__o21ai_1
X_21794_ net166 net161 VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26321_ _05392_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23533_ _02932_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20745_ _11407_ _12491_ _12590_ _12591_ VGND VGND VPWR VPWR _12594_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_148_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26252_ spi0.data_packed\[24\] spi0.data_packed\[25\] net698 VGND VGND VPWR VPWR
+ _05358_ sky130_fd_sc_hd__mux2_1
X_23464_ _02896_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__clkbuf_1
X_20676_ net249 _12499_ VGND VGND VPWR VPWR _12525_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25203_ _04548_ _04549_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22415_ _01972_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__inv_2
X_26183_ spi0.data_packed\[10\] _05318_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__xor2_1
X_23395_ net215 _11560_ _02833_ _11654_ _02834_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__o221a_2
XFILLER_0_6_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25134_ _03474_ _03936_ _04421_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__and3_1
XFILLER_0_162_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22346_ _01845_ _01904_ _01230_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25065_ _04412_ _04413_ _04258_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__mux2_1
X_22277_ _01113_ _01412_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__nor2_1
X_24016_ _03320_ _03373_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__xnor2_4
X_21228_ _13070_ _13071_ _13067_ VGND VGND VPWR VPWR _13072_ sky130_fd_sc_hd__mux2_1
Xhold170 top0.matmul0.matmul_stage_inst.c\[1\] VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _00317_ VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 top0.pid_d.prev_error\[2\] VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__dlygate4sd3_1
X_21159_ _13000_ _13003_ VGND VGND VPWR VPWR _13004_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout650 net653 VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__clkbuf_4
Xfanout661 net663 VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__clkbuf_2
Xfanout672 net673 VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__buf_2
Xfanout683 net685 VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__buf_2
X_13981_ _05657_ _05718_ _05720_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__or3_1
X_25967_ _05175_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__clkbuf_1
Xfanout694 net695 VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15720_ _07813_ _07816_ VGND VGND VPWR VPWR _07817_ sky130_fd_sc_hd__xnor2_2
X_24918_ _04198_ _04210_ _04195_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__o21ba_1
X_25898_ net429 _05113_ _05114_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15651_ _07743_ _07748_ VGND VGND VPWR VPWR _07749_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_186_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24849_ net1017 _03112_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14602_ _06689_ _06806_ VGND VGND VPWR VPWR _06807_ sky130_fd_sc_hd__nor2_1
XFILLER_0_185_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18370_ net391 net317 VGND VGND VPWR VPWR _10351_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_1_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15582_ _07680_ _07588_ _07293_ VGND VGND VPWR VPWR _07681_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_200_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17321_ top0.matmul0.matmul_stage_inst.mult1\[11\] top0.matmul0.matmul_stage_inst.mult2\[11\]
+ VGND VGND VPWR VPWR _09313_ sky130_fd_sc_hd__xor2_1
X_14533_ _06699_ _06739_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_185_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26519_ clknet_leaf_66_clk_sys _00142_ net659 VGND VGND VPWR VPWR top0.pid_q.out\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17252_ top0.matmul0.matmul_stage_inst.mult1\[1\] top0.matmul0.matmul_stage_inst.mult2\[1\]
+ VGND VGND VPWR VPWR _09254_ sky130_fd_sc_hd__xor2_1
X_14464_ _06661_ _06671_ VGND VGND VPWR VPWR _06672_ sky130_fd_sc_hd__xor2_4
XFILLER_0_153_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16203_ net468 net501 _08289_ _08294_ net497 VGND VGND VPWR VPWR _08295_ sky130_fd_sc_hd__a32o_2
X_13415_ _05623_ _05627_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17183_ _09193_ _09187_ _08324_ VGND VGND VPWR VPWR _09194_ sky130_fd_sc_hd__o21a_1
XFILLER_0_183_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14395_ _06481_ _06487_ VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__xnor2_1
X_16134_ _08140_ _08147_ _08226_ VGND VGND VPWR VPWR _08227_ sky130_fd_sc_hd__o21a_1
X_13346_ _05509_ _05558_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_144_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16065_ top0.pid_q.out\[5\] _08158_ _07700_ VGND VGND VPWR VPWR _08159_ sky130_fd_sc_hd__mux2_1
X_13277_ top0.matmul0.beta_pass\[1\] _05466_ _05470_ _05464_ top0.c_out_calc\[1\]
+ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__a32oi_4
X_15016_ _07133_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19824_ _11514_ _11700_ _11702_ VGND VGND VPWR VPWR _11703_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_166_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19755_ _11612_ _11637_ VGND VGND VPWR VPWR _11638_ sky130_fd_sc_hd__nand2_1
X_16967_ net455 _08861_ VGND VGND VPWR VPWR _09024_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18706_ _10676_ VGND VGND VPWR VPWR _10683_ sky130_fd_sc_hd__inv_2
X_15918_ net455 net521 VGND VGND VPWR VPWR _08013_ sky130_fd_sc_hd__nand2_1
X_16898_ _08957_ _08958_ _05601_ VGND VGND VPWR VPWR _08959_ sky130_fd_sc_hd__a21o_1
X_19686_ _11419_ VGND VGND VPWR VPWR _11572_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18637_ net316 _10613_ _10614_ _10208_ VGND VGND VPWR VPWR _10615_ sky130_fd_sc_hd__a22o_1
X_15849_ _07839_ _07838_ VGND VGND VPWR VPWR _07945_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_56_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18568_ _10544_ _10546_ VGND VGND VPWR VPWR _10547_ sky130_fd_sc_hd__xor2_2
XFILLER_0_75_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17519_ _09424_ VGND VGND VPWR VPWR _09506_ sky130_fd_sc_hd__inv_2
XFILLER_0_185_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18499_ _10477_ _10478_ VGND VGND VPWR VPWR _10479_ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20530_ _12283_ _12314_ VGND VGND VPWR VPWR _12379_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20461_ net288 _12308_ _12309_ net303 VGND VGND VPWR VPWR _12310_ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22200_ net104 net100 net95 VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__and3b_1
X_23180_ _02647_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__buf_6
XFILLER_0_171_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20392_ _12233_ _12240_ VGND VGND VPWR VPWR _12241_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_65_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22131_ _01692_ _01691_ _01221_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22062_ _01557_ _01621_ _01622_ _01623_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_101_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21013_ _12858_ _12859_ VGND VGND VPWR VPWR _12860_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26870_ clknet_leaf_36_clk_sys _00487_ net678 VGND VGND VPWR VPWR top0.svm0.tA\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25821_ top0.matmul0.alpha_pass\[2\] top0.matmul0.beta_pass\[2\] VGND VGND VPWR VPWR
+ _05046_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25752_ net69 top0.matmul0.cos\[4\] _05458_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22964_ top0.svm0.delta\[6\] _02474_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_74_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24703_ _04053_ _04056_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__xor2_1
X_21915_ _01472_ _01475_ _01471_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__a21bo_1
X_25683_ _04884_ _04951_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__and2_1
X_22895_ top0.svm0.tC\[3\] _02412_ _02339_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__a21o_1
X_24634_ _03984_ _03987_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_139_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21846_ _01122_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24565_ _03916_ _03917_ _03918_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__and3_1
X_21777_ net135 _01338_ _01330_ _01327_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__a211o_1
X_26304_ spi0.data_packed\[50\] spi0.data_packed\[51\] net697 VGND VGND VPWR VPWR
+ _05384_ sky130_fd_sc_hd__mux2_1
X_23516_ _02923_ VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__clkbuf_1
X_20728_ _12501_ _12576_ VGND VGND VPWR VPWR _12577_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27284_ clknet_3_2__leaf_clk_mosi _00898_ VGND VGND VPWR VPWR spi0.data_packed\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24496_ _03663_ _03849_ _03850_ _03676_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_65_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26235_ _05349_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23447_ _11650_ _02882_ _11954_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__a21o_1
XFILLER_0_191_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20659_ _12156_ _12506_ net294 VGND VGND VPWR VPWR _12508_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_83_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13200_ spi0.cs_sync\[2\] _05428_ _05429_ spi0.cs_sync\[1\] VGND VGND VPWR VPWR _05430_
+ sky130_fd_sc_hd__nor4b_4
XFILLER_0_162_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14180_ _06356_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__inv_2
X_26166_ _05305_ top0.cordic0.slte0.opB\[8\] _12006_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23378_ net1014 _02819_ net178 VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25117_ _04405_ _04408_ _04465_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22329_ _01745_ _01867_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26097_ _05274_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__dlymetal6s2s_1
X_25048_ _04306_ _04392_ _04394_ _04397_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__a31o_1
X_17870_ _09843_ _09856_ VGND VGND VPWR VPWR _09857_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16821_ net496 _08861_ VGND VGND VPWR VPWR _08888_ sky130_fd_sc_hd__or2_1
X_26999_ clknet_leaf_24_clk_sys _00616_ net626 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout480 net481 VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_92_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout491 net492 VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__clkbuf_4
X_16752_ _08453_ _08835_ VGND VGND VPWR VPWR _08836_ sky130_fd_sc_hd__nor2_1
X_19540_ _11429_ VGND VGND VPWR VPWR _11430_ sky130_fd_sc_hd__clkbuf_4
X_13964_ _05799_ _06083_ _05857_ _06176_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__a211o_1
X_15703_ _05443_ VGND VGND VPWR VPWR _07800_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16683_ _08764_ _08767_ VGND VGND VPWR VPWR _08768_ sky130_fd_sc_hd__xnor2_1
X_19471_ top0.pid_d.prev_int\[10\] VGND VGND VPWR VPWR _11366_ sky130_fd_sc_hd__inv_2
X_13895_ _06105_ _06107_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__xor2_2
XFILLER_0_201_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18422_ net406 net402 _09967_ VGND VGND VPWR VPWR _10403_ sky130_fd_sc_hd__and3_1
X_15634_ _07723_ _07731_ VGND VGND VPWR VPWR _07732_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_150_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18353_ top0.pid_d.out\[5\] _10334_ net14 VGND VGND VPWR VPWR _10335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15565_ _07557_ _07558_ _07559_ VGND VGND VPWR VPWR _07664_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17304_ top0.matmul0.matmul_stage_inst.mult2\[8\] VGND VGND VPWR VPWR _09298_ sky130_fd_sc_hd__inv_2
X_14516_ net30 _06717_ _06719_ _05822_ _06722_ VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__o221a_1
X_18284_ _10260_ _10265_ VGND VGND VPWR VPWR _10266_ sky130_fd_sc_hd__xor2_2
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15496_ _07586_ _07587_ _07593_ VGND VGND VPWR VPWR _07595_ sky130_fd_sc_hd__or3b_1
X_17235_ top0.pid_q.prev_int\[14\] _09239_ VGND VGND VPWR VPWR _09240_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14447_ net49 _06131_ _06562_ _06563_ VGND VGND VPWR VPWR _06655_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17166_ top0.pid_q.curr_int\[6\] top0.pid_q.prev_int\[6\] VGND VGND VPWR VPWR _09179_
+ sky130_fd_sc_hd__xnor2_1
X_14378_ _06583_ _06586_ VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_49_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16117_ _08207_ _08209_ VGND VGND VPWR VPWR _08210_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13329_ top0.matmul0.alpha_pass\[7\] _05434_ _05467_ VGND VGND VPWR VPWR _05542_
+ sky130_fd_sc_hd__and3_1
X_17097_ top0.pid_q.curr_error\[7\] _08860_ _09117_ VGND VGND VPWR VPWR _09125_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16048_ net483 _08003_ net499 VGND VGND VPWR VPWR _08142_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_161_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19807_ net1013 _11686_ _11673_ VGND VGND VPWR VPWR _11688_ sky130_fd_sc_hd__a21oi_1
X_17999_ top0.pid_d.out\[2\] top0.pid_d.curr_int\[2\] VGND VGND VPWR VPWR _09984_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_193_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19738_ _11584_ _11619_ VGND VGND VPWR VPWR _11622_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_55_clk_sys clknet_3_4__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_55_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_196_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19669_ net103 net98 net200 VGND VGND VPWR VPWR _11556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21700_ net131 _01259_ _01261_ _01080_ _01079_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__a221o_4
XFILLER_0_56_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22680_ _02228_ _02208_ _02231_ net210 VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_59_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21631_ _01085_ _01192_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_176_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24350_ _03703_ _03704_ _03705_ _03706_ VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_173_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21562_ net132 _01122_ _01123_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23301_ _11650_ _02747_ net1020 VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20513_ _12280_ _12360_ _12361_ VGND VGND VPWR VPWR _12362_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24281_ _03450_ _03618_ _03638_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__or3_1
X_21493_ _01044_ _01053_ _01056_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26020_ top0.pid_q.out\[14\] _05198_ _05199_ spi0.data_packed\[62\] VGND VGND VPWR
+ VPWR _05216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20444_ net271 net265 VGND VGND VPWR VPWR _12293_ sky130_fd_sc_hd__nand2_1
X_23232_ _02680_ _02681_ _11511_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23163_ _02641_ _06380_ _02645_ net795 VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20375_ net283 _12127_ VGND VGND VPWR VPWR _12224_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22114_ _01637_ _01675_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__nor2_1
X_23094_ net171 _07114_ _02594_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__o21a_2
XFILLER_0_100_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22045_ _01334_ _01347_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__nor2_1
X_26922_ clknet_leaf_3_clk_sys _00539_ net581 VGND VGND VPWR VPWR top0.matmul0.cos\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_26853_ clknet_leaf_47_clk_sys _00470_ net676 VGND VGND VPWR VPWR top0.svm0.delta\[13\]
+ sky130_fd_sc_hd__dfrtp_2
X_25804_ top0.matmul0.alpha_pass\[0\] top0.matmul0.beta_pass\[0\] VGND VGND VPWR VPWR
+ _05032_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26784_ clknet_leaf_109_clk_sys _00401_ net578 VGND VGND VPWR VPWR top0.cordic0.sin\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_23996_ _02993_ _02995_ _03063_ _03064_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__o22a_2
XFILLER_0_97_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25735_ top0.matmul0.sin\[12\] _04987_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__xnor2_1
X_22947_ _02459_ _02447_ _02452_ _02339_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13680_ _05488_ _05490_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25666_ top0.matmul0.sin\[7\] _04931_ _04884_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__o21a_1
X_22878_ net169 _02381_ _02396_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24617_ _03968_ _03969_ _03967_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__a21o_1
X_21829_ _01385_ _01387_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_78_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25597_ net71 top0.matmul0.cos\[2\] VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15350_ net482 _07443_ _07446_ _07448_ VGND VGND VPWR VPWR _07449_ sky130_fd_sc_hd__a2bb2o_1
X_24548_ _02994_ _02996_ _03018_ _03019_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14301_ _06442_ _06443_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15281_ _07333_ _07378_ _07379_ VGND VGND VPWR VPWR _07380_ sky130_fd_sc_hd__nand3_1
X_27267_ clknet_3_6__leaf_clk_mosi _00881_ VGND VGND VPWR VPWR spi0.data_packed\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24479_ _03833_ _03834_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17020_ _09053_ _09071_ _09072_ VGND VGND VPWR VPWR _09073_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14232_ net28 _06331_ _06332_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_124_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26218_ spi0.data_packed\[7\] spi0.data_packed\[8\] net694 VGND VGND VPWR VPWR _05341_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27198_ clknet_leaf_32_clk_sys _00812_ net664 VGND VGND VPWR VPWR top0.currT_r\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14163_ _06256_ _06266_ _06374_ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__a21oi_1
X_26149_ spi0.data_packed\[0\] spi0.data_packed\[15\] spi0.data_packed\[1\] spi0.data_packed\[2\]
+ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__and4_1
XFILLER_0_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14094_ _05688_ _05531_ _05532_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__nor3_1
X_18971_ _09395_ net368 _09356_ VGND VGND VPWR VPWR _10945_ sky130_fd_sc_hd__a21oi_1
X_17922_ _09827_ _09828_ _09829_ VGND VGND VPWR VPWR _09908_ sky130_fd_sc_hd__o21ai_1
X_17853_ _09831_ _09839_ VGND VGND VPWR VPWR _09840_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16804_ net509 _08855_ _08858_ net713 _08875_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14996_ spi0.data_packed\[4\] top0.periodTop\[4\] _07108_ VGND VGND VPWR VPWR _07123_
+ sky130_fd_sc_hd__mux2_1
X_17784_ _09688_ _09706_ VGND VGND VPWR VPWR _09771_ sky130_fd_sc_hd__nor2_2
XFILLER_0_191_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19523_ _11412_ VGND VGND VPWR VPWR _11413_ sky130_fd_sc_hd__buf_2
X_13947_ _06157_ _06159_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_163_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16735_ _08764_ _08762_ _08818_ VGND VGND VPWR VPWR _08819_ sky130_fd_sc_hd__o21a_1
XFILLER_0_199_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16666_ _07213_ _08711_ net459 VGND VGND VPWR VPWR _08751_ sky130_fd_sc_hd__o21a_1
X_19454_ top0.pid_d.prev_int\[8\] VGND VGND VPWR VPWR _11351_ sky130_fd_sc_hd__inv_2
X_13878_ _05565_ _05534_ _05775_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_147_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18405_ net348 _10384_ _10385_ VGND VGND VPWR VPWR _10386_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15617_ _07714_ _07686_ _07677_ VGND VGND VPWR VPWR _07715_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_69_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16597_ _08542_ _08607_ _08605_ VGND VGND VPWR VPWR _08684_ sky130_fd_sc_hd__a21o_1
X_19385_ net437 _07136_ _05441_ VGND VGND VPWR VPWR _11291_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18336_ _10304_ _10317_ VGND VGND VPWR VPWR _10318_ sky130_fd_sc_hd__xnor2_1
X_15548_ _07644_ _07646_ VGND VGND VPWR VPWR _07647_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18267_ _10246_ _10247_ VGND VGND VPWR VPWR _10249_ sky130_fd_sc_hd__or2_1
XFILLER_0_170_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15479_ net540 net451 VGND VGND VPWR VPWR _07578_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17218_ _09217_ _09223_ _09224_ VGND VGND VPWR VPWR _09225_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18198_ _10174_ _10179_ VGND VGND VPWR VPWR _10181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17149_ _09163_ _09154_ _09156_ _08076_ VGND VGND VPWR VPWR _09164_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout7 _08403_ VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__buf_2
X_20160_ net209 net206 VGND VGND VPWR VPWR _12012_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_139_Left_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20091_ _11942_ _11950_ VGND VGND VPWR VPWR _11951_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23850_ _03037_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22801_ _02311_ _02312_ _02320_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23781_ _03035_ _03138_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__or2_1
XFILLER_0_196_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20993_ net267 _12836_ _12838_ _12778_ _12839_ VGND VGND VPWR VPWR _12840_ sky130_fd_sc_hd__a221o_1
X_25520_ _05456_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__buf_4
X_22732_ _01877_ _02278_ _02277_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_148_Left_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25451_ _04791_ _04793_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22663_ _02153_ _02213_ _02214_ _02154_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24402_ _03029_ _03030_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__or2_2
XFILLER_0_133_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21614_ net158 _01175_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__xnor2_1
X_25382_ _04722_ _04725_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_168_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22594_ _01798_ _02147_ _01074_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_30_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27121_ clknet_3_6__leaf_clk_sys _00735_ net665 VGND VGND VPWR VPWR top0.c_out_calc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_24333_ _03045_ _03046_ _03029_ _03030_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__o22a_1
X_21545_ net155 _01105_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27052_ clknet_leaf_20_clk_sys _00669_ net611 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.d\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24264_ _03442_ _03436_ _03621_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__a21o_1
X_21476_ _01014_ _00994_ net1021 VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_161_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26003_ _05168_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__buf_2
X_23215_ net301 net297 net292 net286 net198 net191 VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__mux4_1
X_20427_ _12271_ _12275_ VGND VGND VPWR VPWR _12276_ sky130_fd_sc_hd__xnor2_2
X_24195_ _03010_ _03549_ _03552_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_157_Left_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23146_ _02440_ _02632_ _02596_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__o21ai_1
X_20358_ net246 net239 VGND VGND VPWR VPWR _12207_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_30_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23077_ net64 _02352_ _02574_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__or3b_1
X_20289_ net250 net244 VGND VGND VPWR VPWR _12138_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22028_ _01560_ _01589_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__xnor2_2
X_26905_ clknet_leaf_4_clk_sys _00522_ net580 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold30 top0.matmul0.matmul_stage_inst.a\[13\] VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold41 top0.periodTop\[4\] VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 top0.matmul0.matmul_stage_inst.d\[11\] VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ _07044_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__clkbuf_1
X_26836_ clknet_leaf_36_clk_sys _00453_ net678 VGND VGND VPWR VPWR top0.svm0.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold63 top0.cordic0.cos\[7\] VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 top0.svm0.tB\[10\] VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 top0.cordic0.cos\[9\] VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ net68 _06010_ _06012_ _06013_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__o211ai_2
Xhold96 top0.kpq\[10\] VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ _06981_ VGND VGND VPWR VPWR _06982_ sky130_fd_sc_hd__inv_2
X_26767_ clknet_leaf_4_clk_sys _00384_ net580 VGND VGND VPWR VPWR top0.cordic0.cos\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23979_ _03027_ _03028_ VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__or2_2
XFILLER_0_202_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16520_ _08542_ _08605_ _08607_ VGND VGND VPWR VPWR _08608_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_168_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13732_ _05889_ _05944_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__xnor2_1
X_25718_ net764 _04964_ _04936_ _04976_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26698_ clknet_leaf_64_clk_sys _00315_ net648 VGND VGND VPWR VPWR top0.pid_d.prev_error\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16451_ _08532_ _08539_ VGND VGND VPWR VPWR _08540_ sky130_fd_sc_hd__xnor2_2
X_13663_ _05828_ _05809_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__xor2_1
X_25649_ _04890_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15402_ _07414_ _07500_ VGND VGND VPWR VPWR _07501_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19170_ net440 _11118_ _11121_ top0.matmul0.alpha_pass\[0\] _11123_ VGND VGND VPWR
+ VPWR _11124_ sky130_fd_sc_hd__a221o_1
X_16382_ _08142_ _08383_ _08381_ _08386_ VGND VGND VPWR VPWR _08472_ sky130_fd_sc_hd__or4_1
X_13594_ net66 _05641_ _05806_ _05731_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18121_ _10103_ _10010_ _10104_ VGND VGND VPWR VPWR _10105_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_54_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15333_ _07425_ _07431_ VGND VGND VPWR VPWR _07432_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18052_ _10022_ _10036_ VGND VGND VPWR VPWR _10037_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15264_ _07355_ _07360_ _07362_ VGND VGND VPWR VPWR _07363_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17003_ top0.matmul0.beta_pass\[12\] _09042_ _05436_ top0.matmul0.beta_pass\[11\]
+ VGND VGND VPWR VPWR _09057_ sky130_fd_sc_hd__o211a_1
X_14215_ net27 _05523_ _05524_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__and3_2
XFILLER_0_22_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_5 _03020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15195_ _07193_ _07191_ VGND VGND VPWR VPWR _07294_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14146_ _06344_ _06357_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_46_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14077_ net45 _05602_ _05603_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__and3_1
X_18954_ _10857_ _10890_ VGND VGND VPWR VPWR _10928_ sky130_fd_sc_hd__and2b_1
X_17905_ _09823_ _09891_ VGND VGND VPWR VPWR _09892_ sky130_fd_sc_hd__nand2_1
X_18885_ _09356_ net360 _10781_ _10859_ VGND VGND VPWR VPWR _10860_ sky130_fd_sc_hd__a31o_1
XFILLER_0_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17836_ _09746_ _09821_ _09822_ VGND VGND VPWR VPWR _09823_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17767_ _09662_ _09682_ VGND VGND VPWR VPWR _09754_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14979_ spi0.data_packed\[31\] top0.kiq\[15\] _07108_ VGND VGND VPWR VPWR _07112_
+ sky130_fd_sc_hd__mux2_1
X_19506_ _10993_ _11027_ _11077_ VGND VGND VPWR VPWR _11397_ sky130_fd_sc_hd__o21a_1
X_16718_ _08754_ _08777_ _08778_ VGND VGND VPWR VPWR _08802_ sky130_fd_sc_hd__a21o_1
X_17698_ _09647_ _09684_ VGND VGND VPWR VPWR _09685_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19437_ _11334_ _11330_ _11335_ VGND VGND VPWR VPWR _11336_ sky130_fd_sc_hd__a21o_1
X_16649_ _08732_ _08734_ VGND VGND VPWR VPWR _08735_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19368_ net961 _11285_ _11288_ top0.pid_d.curr_error\[1\] VGND VGND VPWR VPWR _00311_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18319_ _10299_ _10300_ VGND VGND VPWR VPWR _10301_ sky130_fd_sc_hd__nor2_1
X_19299_ top0.matmul0.alpha_pass\[11\] top0.matmul0.alpha_pass\[12\] _11221_ VGND
+ VGND VPWR VPWR _11241_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21330_ _13001_ _13170_ VGND VGND VPWR VPWR _13172_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21261_ _13103_ _13104_ VGND VGND VPWR VPWR _13105_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23000_ _06277_ _02505_ net171 VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20212_ net304 net281 VGND VGND VPWR VPWR _12061_ sky130_fd_sc_hd__xnor2_1
X_21192_ net213 _13035_ VGND VGND VPWR VPWR _13036_ sky130_fd_sc_hd__nand2_2
XFILLER_0_60_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20143_ net1020 _11983_ _11991_ _11992_ _11998_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__o32a_1
XFILLER_0_25_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24951_ _04270_ _04301_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__xor2_2
X_20074_ net913 _11934_ _11935_ _11933_ VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23902_ _03237_ _03242_ _03256_ _03259_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__a2bb2o_1
X_24882_ _04214_ _04233_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__xnor2_1
X_26621_ clknet_leaf_25_clk_sys _00238_ net627 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_23833_ _03184_ _03190_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_174_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26552_ clknet_leaf_51_clk_sys _00175_ net671 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23764_ _03090_ _03091_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20976_ _12072_ _12820_ VGND VGND VPWR VPWR _12823_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25503_ _04837_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22715_ _02207_ _02224_ _02264_ _02265_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__o31a_1
XFILLER_0_165_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26483_ clknet_leaf_11_clk_sys _00114_ net604 VGND VGND VPWR VPWR top0.periodTop\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_23695_ _03042_ _03044_ _03052_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__o21a_1
XFILLER_0_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25434_ _04726_ _04730_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22646_ _02192_ _02198_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_192_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25365_ _04661_ _04709_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22577_ net211 _02131_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27104_ clknet_leaf_21_clk_sys _00721_ net610 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.a\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_24316_ _03087_ _03672_ _03669_ _03110_ VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__o2bb2a_1
X_21528_ net122 _01089_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25296_ _04631_ _04641_ _03829_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_133_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27035_ clknet_leaf_8_clk_sys _00652_ net595 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_24247_ _03603_ _03570_ _03601_ _03602_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__a22o_1
X_21459_ _01023_ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14000_ _05683_ _06211_ _06212_ _05894_ net1030 VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__o32a_1
XFILLER_0_181_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24178_ _03478_ _03533_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__nand2_1
Xoutput7 net7 VGND VGND VPWR VPWR ready sky130_fd_sc_hd__buf_2
X_23129_ top0.svm0.delta\[10\] _02620_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15951_ _07907_ _07908_ _07906_ VGND VGND VPWR VPWR _08046_ sky130_fd_sc_hd__o21ai_1
X_14902_ _07071_ VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__clkbuf_1
X_18670_ _10646_ _10647_ VGND VGND VPWR VPWR _10648_ sky130_fd_sc_hd__and2b_1
X_15882_ _07976_ _07977_ VGND VGND VPWR VPWR _07978_ sky130_fd_sc_hd__or2b_1
X_17621_ _09604_ _09607_ VGND VGND VPWR VPWR _09608_ sky130_fd_sc_hd__xnor2_2
X_14833_ _07020_ _07031_ VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__xnor2_1
X_26819_ clknet_leaf_48_clk_sys _00436_ net676 VGND VGND VPWR VPWR top0.svm0.state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14764_ _06960_ _06965_ VGND VGND VPWR VPWR _06966_ sky130_fd_sc_hd__xnor2_1
X_17552_ _09349_ _09538_ VGND VGND VPWR VPWR _09539_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13715_ _05918_ _05927_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__xnor2_2
X_16503_ _08588_ _08590_ VGND VGND VPWR VPWR _08591_ sky130_fd_sc_hd__xnor2_1
X_17483_ net398 net350 VGND VGND VPWR VPWR _09470_ sky130_fd_sc_hd__nand2_1
X_14695_ _06879_ _06898_ VGND VGND VPWR VPWR _06899_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19222_ net76 _11160_ VGND VGND VPWR VPWR _11171_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13646_ _05809_ _05852_ _05850_ _05854_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__o211a_1
X_16434_ _08429_ _08440_ _08522_ VGND VGND VPWR VPWR _08523_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16365_ _08446_ _08454_ VGND VGND VPWR VPWR _08455_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19153_ top0.kid\[11\] _11097_ _11099_ top0.kpd\[11\] VGND VGND VPWR VPWR _11112_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13577_ net66 net63 _05619_ _05666_ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__nand4_2
XFILLER_0_13_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18104_ _10077_ _10087_ VGND VGND VPWR VPWR _10088_ sky130_fd_sc_hd__xnor2_2
X_15316_ _07408_ _07409_ _07414_ VGND VGND VPWR VPWR _07415_ sky130_fd_sc_hd__o21ba_1
X_16296_ _08384_ _08386_ VGND VGND VPWR VPWR _08387_ sky130_fd_sc_hd__xnor2_1
X_19084_ _10384_ net308 _09965_ VGND VGND VPWR VPWR _11056_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18035_ _10016_ _10019_ VGND VGND VPWR VPWR _10020_ sky130_fd_sc_hd__xnor2_2
X_15247_ _07304_ _07319_ _07342_ VGND VGND VPWR VPWR _07346_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15178_ _07275_ _07276_ VGND VGND VPWR VPWR _07277_ sky130_fd_sc_hd__xnor2_1
X_14129_ _06304_ _06305_ _06340_ VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout309 net310 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__clkbuf_4
X_19986_ _11837_ _11838_ _11853_ VGND VGND VPWR VPWR _11854_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18937_ _10910_ _10911_ VGND VGND VPWR VPWR _10912_ sky130_fd_sc_hd__or2b_1
XFILLER_0_158_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18868_ _10787_ _10806_ _10842_ VGND VGND VPWR VPWR _10843_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17819_ _09804_ _09805_ VGND VGND VPWR VPWR _09806_ sky130_fd_sc_hd__and2b_1
X_18799_ _10773_ _10774_ VGND VGND VPWR VPWR _10775_ sky130_fd_sc_hd__xor2_2
XFILLER_0_55_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20830_ _12223_ _12226_ _12217_ _12211_ _12210_ VGND VGND VPWR VPWR _12679_ sky130_fd_sc_hd__a311o_1
XFILLER_0_89_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20761_ net263 _12337_ VGND VGND VPWR VPWR _12610_ sky130_fd_sc_hd__xor2_4
XFILLER_0_9_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22500_ _01213_ net107 _02020_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__or3_1
XFILLER_0_130_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23480_ net999 top0.matmul0.sin\[9\] _02904_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20692_ _12460_ _12461_ _12540_ VGND VGND VPWR VPWR _12541_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22431_ _01896_ _01988_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25150_ _04428_ _04430_ _04497_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__o21a_1
X_22362_ _01917_ _01920_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24101_ _03207_ _03208_ _03015_ _03016_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__o22a_1
XFILLER_0_143_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21313_ net1021 _13154_ VGND VGND VPWR VPWR _13155_ sky130_fd_sc_hd__nor2_1
X_25081_ _03280_ _04190_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22293_ net87 _01852_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24032_ _02994_ _02996_ _03088_ _03089_ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__o22a_2
X_21244_ _12660_ _12575_ _13087_ _12546_ VGND VGND VPWR VPWR _13088_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_13_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21175_ net246 _12982_ VGND VGND VPWR VPWR _13019_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20126_ _11975_ _11979_ _11980_ _11982_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__o211a_1
X_25983_ _05187_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24934_ _04276_ _04284_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__xnor2_2
X_20057_ top0.cordic0.slte0.opA\[8\] _11907_ _11919_ VGND VGND VPWR VPWR _11920_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_197_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24865_ _04215_ _04216_ _04069_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23816_ _03119_ _03172_ _03173_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__a21o_1
X_26604_ clknet_leaf_51_clk_sys _00227_ net670 VGND VGND VPWR VPWR top0.pid_q.curr_int\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_200_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24796_ _04035_ _04142_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26535_ clknet_leaf_60_clk_sys _00158_ net652 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_23747_ _03088_ _03089_ _03103_ _03104_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__o22a_2
XFILLER_0_23_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20959_ _12737_ VGND VGND VPWR VPWR _12807_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13500_ _05710_ _05712_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__xnor2_1
X_14480_ _06673_ VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__inv_2
X_26466_ clknet_leaf_17_clk_sys _00000_ net611 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.state\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_95_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23678_ net568 top0.matmul0.matmul_stage_inst.b\[4\] top0.matmul0.matmul_stage_inst.a\[4\]
+ net564 VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__a22o_2
XFILLER_0_95_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25417_ _04661_ _04760_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__nor2_1
X_13431_ _05582_ _05592_ _05584_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22629_ _02094_ _02124_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__or2b_1
X_26397_ clknet_leaf_79_clk_sys _00038_ net632 VGND VGND VPWR VPWR top0.kpd\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16150_ _08236_ _08242_ _07710_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__o21a_1
X_25348_ _04561_ _04630_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__nand2_1
X_13362_ _05571_ _05572_ _05574_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15101_ _07198_ _07199_ VGND VGND VPWR VPWR _07200_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16081_ _08049_ _08173_ VGND VGND VPWR VPWR _08174_ sky130_fd_sc_hd__xnor2_2
X_25279_ _04619_ _04624_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__xor2_2
X_13293_ _05503_ _05505_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__xnor2_1
X_27018_ clknet_leaf_16_clk_sys _00635_ net613 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_15032_ net971 _07140_ _07144_ top0.pid_d.curr_int\[2\] VGND VGND VPWR VPWR _00119_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19840_ _11717_ VGND VGND VPWR VPWR _11718_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19771_ net259 VGND VGND VPWR VPWR _11653_ sky130_fd_sc_hd__inv_2
X_16983_ top0.currT_r\[11\] _09033_ VGND VGND VPWR VPWR _09038_ sky130_fd_sc_hd__nand2_1
X_18722_ _10697_ _10698_ VGND VGND VPWR VPWR _10699_ sky130_fd_sc_hd__xor2_1
X_15934_ net461 net516 VGND VGND VPWR VPWR _08029_ sky130_fd_sc_hd__nand2_1
X_18653_ _10543_ _10547_ _10630_ VGND VGND VPWR VPWR _10631_ sky130_fd_sc_hd__o21a_1
XFILLER_0_189_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15865_ _07959_ _07960_ VGND VGND VPWR VPWR _07961_ sky130_fd_sc_hd__or2b_1
X_17604_ _09588_ _09589_ _09590_ VGND VGND VPWR VPWR _09591_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_192_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14816_ net21 _06824_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__nand2_1
X_18584_ net397 net393 _09967_ VGND VGND VPWR VPWR _10563_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15796_ _07812_ _07891_ VGND VGND VPWR VPWR _07893_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17535_ net422 net343 VGND VGND VPWR VPWR _09522_ sky130_fd_sc_hd__nand2_1
X_14747_ _06913_ _06937_ _06948_ VGND VGND VPWR VPWR _06949_ sky130_fd_sc_hd__o21a_2
XFILLER_0_15_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14678_ _06832_ _06212_ _06880_ net25 VGND VGND VPWR VPWR _06882_ sky130_fd_sc_hd__o22a_1
X_17466_ _09427_ _09438_ VGND VGND VPWR VPWR _09453_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19205_ _11154_ _11145_ top0.pid_d.prev_error\[3\] VGND VGND VPWR VPWR _11155_ sky130_fd_sc_hd__o21ba_1
X_16417_ _08500_ _08505_ VGND VGND VPWR VPWR _08506_ sky130_fd_sc_hd__xnor2_1
X_13629_ _05839_ _05840_ _05841_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__a21oi_1
X_17397_ _09380_ _09383_ VGND VGND VPWR VPWR _09384_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19136_ net421 _11096_ _11103_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__a21o_1
XFILLER_0_171_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16348_ _08365_ _08366_ _08437_ VGND VGND VPWR VPWR _08438_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_54_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16279_ _08262_ _08264_ _08263_ VGND VGND VPWR VPWR _08370_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19067_ _11016_ _11038_ VGND VGND VPWR VPWR _11039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18018_ _09925_ _09927_ _10002_ VGND VGND VPWR VPWR _10003_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout106 top0.cordic0.vec\[1\]\[12\] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout117 top0.cordic0.vec\[1\]\[10\] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_1
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout128 net129 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_4
Xfanout139 top0.cordic0.vec\[1\]\[5\] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__buf_4
X_19969_ _11822_ _11829_ top0.cordic0.slte0.opA\[2\] VGND VGND VPWR VPWR _11838_ sky130_fd_sc_hd__a21boi_1
X_22980_ _06277_ _02488_ net172 VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21931_ _01483_ _01492_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24650_ _03864_ _03865_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__nor2_1
X_21862_ _01399_ _01390_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23601_ _02967_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20813_ _12575_ _12578_ _12606_ _12647_ VGND VGND VPWR VPWR _12662_ sky130_fd_sc_hd__a211o_1
X_24581_ _03826_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21793_ _01262_ _01354_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_132_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26320_ spi0.data_packed\[58\] spi0.data_packed\[59\] net698 VGND VGND VPWR VPWR
+ _05392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23532_ top0.a_in_matmul\[6\] top0.matmul0.a\[6\] _02926_ VGND VGND VPWR VPWR _02932_
+ sky130_fd_sc_hd__mux2_1
X_20744_ _12590_ _12591_ _12592_ VGND VGND VPWR VPWR _12593_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26251_ _05357_ VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23463_ net1003 top0.matmul0.sin\[1\] _05461_ VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__mux2_1
X_20675_ net263 _11689_ _12499_ _12523_ _12493_ VGND VGND VPWR VPWR _12524_ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25202_ net1017 _04182_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22414_ net86 net80 _01923_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26182_ spi0.data_packed\[8\] spi0.data_packed\[9\] _05310_ net18 VGND VGND VPWR
+ VPWR _05318_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23394_ _11714_ _02650_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__or2_1
X_25133_ _03343_ _04272_ _04420_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22345_ net78 _01903_ _01900_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25064_ _03355_ _04252_ _04131_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__and3_1
X_22276_ _01113_ _01412_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__nand2_1
X_24015_ _03308_ _03311_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__xnor2_2
Xhold160 top0.pid_q.prev_error\[4\] VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__dlygate4sd3_1
X_21227_ _12620_ _12627_ VGND VGND VPWR VPWR _13071_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold171 top0.matmul0.matmul_stage_inst.b\[2\] VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 top0.svm0.tA\[12\] VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 _00312_ VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__dlygate4sd3_1
X_21158_ _13001_ _13002_ VGND VGND VPWR VPWR _13003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout640 net645 VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__clkbuf_4
Xfanout651 net653 VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__clkbuf_4
Xfanout662 net663 VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__clkbuf_4
X_20109_ _11965_ _11966_ VGND VGND VPWR VPWR _11967_ sky130_fd_sc_hd__or2_1
X_13980_ _06192_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_176_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout673 net674 VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__clkbuf_2
X_25966_ net998 _05174_ _05165_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__mux2_1
X_21089_ _12892_ _12934_ VGND VGND VPWR VPWR _12935_ sky130_fd_sc_hd__xnor2_1
Xfanout684 net685 VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__clkbuf_4
Xfanout695 net696 VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24917_ _04262_ _04267_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__xnor2_4
X_25897_ _05102_ _05104_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__and2b_1
X_15650_ _07745_ _07747_ VGND VGND VPWR VPWR _07748_ sky130_fd_sc_hd__xor2_1
X_24848_ _03254_ _03280_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14601_ _06802_ _06803_ _06804_ _06805_ VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__o211a_1
X_15581_ _07281_ VGND VGND VPWR VPWR _07680_ sky130_fd_sc_hd__inv_2
X_24779_ _03017_ _03185_ _04131_ _03047_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__o22a_1
XFILLER_0_197_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14532_ _06737_ _06738_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__nor2_2
X_17320_ _09310_ _09306_ _09311_ VGND VGND VPWR VPWR _09312_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26518_ clknet_leaf_67_clk_sys _00141_ net659 VGND VGND VPWR VPWR top0.pid_q.out\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_154_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14463_ _06662_ _06663_ _06666_ _06560_ _06670_ VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__o221a_2
X_17251_ top0.matmul0.matmul_stage_inst.mult1\[0\] top0.matmul0.matmul_stage_inst.mult2\[0\]
+ VGND VGND VPWR VPWR _09253_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26449_ clknet_leaf_55_clk_sys _00090_ net667 VGND VGND VPWR VPWR top0.kiq\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_187_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13414_ _05621_ _05622_ _05626_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__a21oi_1
X_16202_ _08288_ _08290_ _08292_ net473 _08293_ VGND VGND VPWR VPWR _08294_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17182_ top0.pid_q.prev_int\[7\] VGND VGND VPWR VPWR _09193_ sky130_fd_sc_hd__inv_2
X_14394_ _06560_ _06602_ VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16133_ _08140_ _08147_ _08137_ VGND VGND VPWR VPWR _08226_ sky130_fd_sc_hd__a21o_1
X_13345_ _05529_ _05557_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16064_ net545 _08085_ _08086_ net548 _08157_ VGND VGND VPWR VPWR _08158_ sky130_fd_sc_hd__a32o_1
X_13276_ _05488_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__buf_2
X_15015_ spi0.data_packed\[13\] top0.periodTop\[13\] _07125_ VGND VGND VPWR VPWR _07133_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_102_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19823_ _11560_ _11557_ _11701_ VGND VGND VPWR VPWR _11702_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19754_ _11635_ _11636_ _11632_ VGND VGND VPWR VPWR _11637_ sky130_fd_sc_hd__mux2_1
X_16966_ net552 _09021_ _09022_ VGND VGND VPWR VPWR _09023_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18705_ _10682_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__clkbuf_1
X_15917_ _07932_ _07942_ _08011_ VGND VGND VPWR VPWR _08012_ sky130_fd_sc_hd__o21a_2
X_19685_ net286 VGND VGND VPWR VPWR _11571_ sky130_fd_sc_hd__inv_2
X_16897_ top0.currT_r\[5\] _08946_ VGND VGND VPWR VPWR _08958_ sky130_fd_sc_hd__or2_1
XFILLER_0_188_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18636_ net377 net316 VGND VGND VPWR VPWR _10614_ sky130_fd_sc_hd__nand2_1
X_15848_ _07932_ _07943_ VGND VGND VPWR VPWR _07944_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_91_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18567_ net362 _10545_ VGND VGND VPWR VPWR _10546_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_111_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15779_ _07873_ _07875_ VGND VGND VPWR VPWR _07876_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17518_ _09418_ _09421_ VGND VGND VPWR VPWR _09505_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18498_ _10471_ _10476_ VGND VGND VPWR VPWR _10478_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17449_ _09356_ _09354_ _09428_ VGND VGND VPWR VPWR _09436_ sky130_fd_sc_hd__o21ba_1
X_20460_ net295 net278 VGND VGND VPWR VPWR _12309_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_51_clk_sys clknet_3_6__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_51_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_19119_ _11078_ _11079_ _11081_ _11090_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__a31o_1
XFILLER_0_162_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20391_ _12236_ _12239_ VGND VGND VPWR VPWR _12240_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22130_ _01225_ _01686_ _01691_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_120_Left_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22061_ _01552_ _01549_ _01553_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21012_ _12849_ _12857_ VGND VGND VPWR VPWR _12859_ sky130_fd_sc_hd__nor2_1
XFILLER_0_199_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25820_ _05043_ _05044_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25751_ net770 _04925_ _04996_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__a21o_1
X_22963_ _02466_ _02468_ _02473_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__a21o_1
X_24702_ _03934_ _04054_ _04055_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__a21oi_2
X_21914_ net166 _01462_ _01475_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25682_ top0.matmul0.sin\[10\] top0.matmul0.sin\[11\] _04942_ VGND VGND VPWR VPWR
+ _04951_ sky130_fd_sc_hd__or3_1
X_22894_ _02347_ top0.svm0.tC\[2\] _02411_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24633_ _03985_ _03986_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__xnor2_1
X_21845_ _01318_ _01365_ _01406_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_38_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24564_ _03916_ _03917_ _03918_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__a21oi_1
X_21776_ net147 net141 VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_33_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26303_ _05383_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__clkbuf_1
X_23515_ top0.cordic0.cos\[12\] top0.matmul0.cos\[12\] _02915_ VGND VGND VPWR VPWR
+ _02923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20727_ _12503_ _12512_ VGND VGND VPWR VPWR _12576_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27283_ clknet_3_0__leaf_clk_mosi _00897_ VGND VGND VPWR VPWR spi0.data_packed\[69\]
+ sky130_fd_sc_hd__dfxtp_1
X_24495_ _03663_ _03751_ _03850_ _03676_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26234_ spi0.data_packed\[15\] spi0.data_packed\[16\] net695 VGND VGND VPWR VPWR
+ _05349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23446_ _02877_ _02881_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20658_ _12156_ _12506_ _11438_ VGND VGND VPWR VPWR _12507_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26165_ spi0.data_packed\[6\] _05304_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23377_ _02810_ _02818_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20589_ net240 _12437_ VGND VGND VPWR VPWR _12438_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25116_ _04461_ _04464_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22328_ _01868_ _01870_ _01867_ VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26096_ _05426_ _05013_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__and2_1
XFILLER_0_182_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25047_ _04395_ _04392_ _04396_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__o21bai_1
X_22259_ _01758_ _01763_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16820_ net550 _08886_ VGND VGND VPWR VPWR _08887_ sky130_fd_sc_hd__and2_1
X_26998_ clknet_leaf_23_clk_sys _00615_ net625 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout470 top0.pid_q.mult0.b\[6\] VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__buf_4
Xfanout481 net482 VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__buf_2
X_16751_ _08526_ _08833_ _08834_ _08312_ VGND VGND VPWR VPWR _08835_ sky130_fd_sc_hd__o22a_1
Xfanout492 top0.pid_q.mult0.b\[1\] VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__buf_4
X_13963_ _06170_ _06175_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__xor2_1
X_25949_ net921 _05028_ _05153_ _05161_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15702_ top0.pid_q.out\[1\] _07700_ _07799_ _07710_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__o211a_1
X_19470_ _10754_ _11341_ _11363_ _11292_ _11365_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__a221o_1
X_16682_ _08765_ _08766_ net498 VGND VGND VPWR VPWR _08767_ sky130_fd_sc_hd__or3b_1
X_13894_ _06106_ _05567_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__nor2_1
X_18421_ _10266_ _10268_ _10401_ VGND VGND VPWR VPWR _10402_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_185_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15633_ _07725_ _07730_ VGND VGND VPWR VPWR _07731_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18352_ net434 _10248_ _10249_ _10333_ net436 VGND VGND VPWR VPWR _10334_ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15564_ _07563_ _07661_ _07662_ VGND VGND VPWR VPWR _07663_ sky130_fd_sc_hd__o21a_2
XFILLER_0_83_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17303_ _09297_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__clkbuf_1
X_14515_ _05579_ _06640_ _06720_ net28 _06721_ VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18283_ _10263_ _10264_ VGND VGND VPWR VPWR _10265_ sky130_fd_sc_hd__xor2_2
X_15495_ _07586_ _07587_ _07593_ VGND VGND VPWR VPWR _07594_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_127_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17234_ top0.pid_q.prev_int\[13\] _09231_ _09238_ VGND VGND VPWR VPWR _09239_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14446_ _06574_ _06579_ _06653_ VGND VGND VPWR VPWR _06654_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_36_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14377_ _06584_ _06585_ VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_181_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17165_ top0.pid_q.prev_int\[5\] _09172_ _09177_ VGND VGND VPWR VPWR _09178_ sky130_fd_sc_hd__o21ai_1
X_13328_ net51 VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__inv_2
X_16116_ _08109_ _08111_ _08208_ VGND VGND VPWR VPWR _08209_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17096_ net842 _09115_ _09124_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13259_ _05468_ _05471_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__nor2_4
X_16047_ net502 VGND VGND VPWR VPWR _08141_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_clk_sys clk_sys VGND VGND VPWR VPWR clknet_0_clk_sys sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19806_ _11430_ _11686_ VGND VGND VPWR VPWR _11687_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17998_ _09981_ _09982_ VGND VGND VPWR VPWR _09983_ sky130_fd_sc_hd__and2_1
XFILLER_0_159_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19737_ _11604_ _11609_ _11611_ _11620_ VGND VGND VPWR VPWR _11621_ sky130_fd_sc_hd__o211ai_4
X_16949_ _09005_ _09006_ VGND VGND VPWR VPWR _09007_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19668_ net199 net84 VGND VGND VPWR VPWR _11555_ sky130_fd_sc_hd__and2b_1
XFILLER_0_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18619_ top0.pid_d.out\[9\] top0.pid_d.curr_int\[9\] VGND VGND VPWR VPWR _10597_
+ sky130_fd_sc_hd__xnor2_1
X_19599_ top0.cordic0.slte0.opA\[7\] _11487_ top0.cordic0.slte0.opB\[7\] VGND VGND
+ VPWR VPWR _11488_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_94_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21630_ _01064_ _01191_ VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__xor2_1
XFILLER_0_177_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21561_ net151 net145 VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__and2_2
XFILLER_0_157_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23300_ _02744_ _02746_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__xnor2_1
X_20512_ _12268_ _12270_ _12275_ VGND VGND VPWR VPWR _12361_ sky130_fd_sc_hd__o21a_1
XFILLER_0_166_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24280_ _03630_ _03632_ VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__or2_1
X_21492_ _12968_ _01038_ _01054_ _01055_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_160_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23231_ _01320_ _02669_ _02659_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__or3b_1
XFILLER_0_166_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20443_ _12286_ _12288_ _12291_ VGND VGND VPWR VPWR _12292_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23162_ _02641_ _06275_ _02645_ net830 VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20374_ _11438_ _12220_ _12221_ _12222_ VGND VGND VPWR VPWR _12223_ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22113_ _01674_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__inv_2
X_23093_ top0.svm0.rising net9 _02305_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22044_ _01362_ _01335_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__or2_1
X_26921_ clknet_leaf_0_clk_sys _00538_ net578 VGND VGND VPWR VPWR top0.matmul0.sin\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_11_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26852_ clknet_leaf_47_clk_sys _00469_ net676 VGND VGND VPWR VPWR top0.svm0.delta\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25803_ _05030_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23995_ _03351_ _03352_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__xnor2_2
X_26783_ clknet_leaf_109_clk_sys _00400_ net579 VGND VGND VPWR VPWR top0.cordic0.sin\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_177_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_170_Right_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22946_ top0.svm0.delta\[3\] VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__inv_2
X_25734_ net72 _04951_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22877_ top0.svm0.tB\[9\] _02394_ _02395_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_195_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25665_ net779 _04904_ _04936_ _04938_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24616_ _03967_ _03968_ _03969_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__nand3_1
X_21828_ net153 _01281_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_149_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25596_ net846 _00000_ _04888_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__o21a_1
XFILLER_0_167_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24547_ _02985_ _02987_ _03029_ _03030_ VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21759_ net147 _01177_ net162 VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14300_ _06501_ _06509_ VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_163_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15280_ _07344_ _07345_ _07346_ _07347_ VGND VGND VPWR VPWR _07379_ sky130_fd_sc_hd__a211o_1
X_24478_ _03821_ _03832_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__nand2_1
X_27266_ clknet_3_6__leaf_clk_mosi _00880_ VGND VGND VPWR VPWR spi0.data_packed\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14231_ _06333_ _06441_ _06331_ VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__mux2_1
X_23429_ _02855_ _02856_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__or2_1
X_26217_ _05340_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__clkbuf_1
X_27197_ clknet_leaf_57_clk_sys _00811_ net664 VGND VGND VPWR VPWR top0.currT_r\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_117_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14162_ _06179_ _06254_ VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26148_ _05291_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14093_ _06233_ _06236_ _06221_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__o21bai_1
X_18970_ _10942_ _10943_ VGND VGND VPWR VPWR _10944_ sky130_fd_sc_hd__xor2_2
X_26079_ _05261_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__clkbuf_1
X_17921_ _09903_ _09906_ VGND VGND VPWR VPWR _09907_ sky130_fd_sc_hd__xnor2_2
X_17852_ _09833_ _09838_ VGND VGND VPWR VPWR _09839_ sky130_fd_sc_hd__xnor2_1
X_16803_ top0.kiq\[11\] _05448_ _08866_ VGND VGND VPWR VPWR _08875_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17783_ _09674_ _09768_ _09769_ VGND VGND VPWR VPWR _09770_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_191_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14995_ _07122_ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__clkbuf_1
X_19522_ _11409_ _11410_ _11411_ VGND VGND VPWR VPWR _11412_ sky130_fd_sc_hd__and3_1
X_16734_ _08764_ _08762_ _08767_ VGND VGND VPWR VPWR _08818_ sky130_fd_sc_hd__a21bo_1
X_13946_ _05734_ _05740_ _06158_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__o21a_1
X_19453_ _10590_ _11341_ _11350_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__a21o_1
XFILLER_0_198_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16665_ _08707_ _08714_ _08713_ VGND VGND VPWR VPWR _08750_ sky130_fd_sc_hd__a21o_1
X_13877_ net47 net43 _05585_ _05587_ _05774_ VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__a41o_1
XFILLER_0_9_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18404_ net348 _10384_ net344 VGND VGND VPWR VPWR _10385_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15616_ _07593_ _07546_ _07547_ _07713_ VGND VGND VPWR VPWR _07714_ sky130_fd_sc_hd__a31o_1
XFILLER_0_202_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19384_ _11289_ VGND VGND VPWR VPWR _11290_ sky130_fd_sc_hd__clkbuf_4
X_16596_ _08599_ _08678_ VGND VGND VPWR VPWR _08683_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18335_ _10306_ _10316_ VGND VGND VPWR VPWR _10317_ sky130_fd_sc_hd__xnor2_1
X_15547_ _07565_ _07566_ _07645_ VGND VGND VPWR VPWR _07646_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18266_ _10246_ _10247_ VGND VGND VPWR VPWR _10248_ sky130_fd_sc_hd__nand2_1
X_15478_ net538 net454 VGND VGND VPWR VPWR _07577_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17217_ top0.pid_q.curr_int\[11\] top0.pid_q.prev_int\[11\] VGND VGND VPWR VPWR _09224_
+ sky130_fd_sc_hd__and2_1
X_14429_ _06437_ _06590_ VGND VGND VPWR VPWR _06637_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18197_ _10174_ _10179_ VGND VGND VPWR VPWR _10180_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17148_ top0.pid_q.prev_int\[3\] VGND VGND VPWR VPWR _09163_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout8 _05444_ VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__buf_4
XFILLER_0_188_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17079_ _09113_ VGND VGND VPWR VPWR _09114_ sky130_fd_sc_hd__buf_2
XFILLER_0_200_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20090_ _11940_ _11941_ top0.cordic0.slte0.opA\[11\] VGND VGND VPWR VPWR _11950_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22800_ _02314_ _02316_ _02318_ _02319_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__or4b_1
XFILLER_0_58_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23780_ _03075_ _03082_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20992_ _12126_ _12778_ VGND VGND VPWR VPWR _12839_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22731_ _12963_ _02279_ _02280_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25450_ _04723_ _04724_ _04792_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22662_ _02159_ _02199_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24401_ _03757_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__clkbuf_1
X_21613_ net131 _01078_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__xnor2_4
X_25381_ _04723_ _04724_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_164_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22593_ top0.cordic0.vec\[1\]\[13\] _01980_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24332_ _03015_ _03016_ _03150_ _03151_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__o22a_1
X_27120_ clknet_leaf_33_clk_sys _00734_ net665 VGND VGND VPWR VPWR top0.c_out_calc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21544_ net155 _01105_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27051_ clknet_leaf_22_clk_sys _00668_ net607 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.d\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24263_ _03442_ _03436_ _03445_ VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__o21a_1
XFILLER_0_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21475_ _01025_ _01039_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__xor2_2
X_26002_ _05202_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23214_ net279 net272 net266 net260 net198 net191 VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__mux4_1
X_20426_ net276 _12108_ _12272_ _12273_ _12274_ VGND VGND VPWR VPWR _12275_ sky130_fd_sc_hd__a221o_2
X_24194_ _03185_ _03114_ _03550_ _03551_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_31_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23145_ _02598_ _02632_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20357_ net229 net221 VGND VGND VPWR VPWR _12206_ sky130_fd_sc_hd__xor2_2
XFILLER_0_101_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23076_ _05607_ top0.svm0.counter\[1\] _02574_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__or3_1
X_20288_ _12135_ _12136_ VGND VGND VPWR VPWR _12137_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22027_ _01568_ _01588_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__xnor2_1
X_26904_ clknet_leaf_4_clk_sys _00521_ net580 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold20 top0.cordic0.sin\[9\] VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 top0.cordic0.cos\[4\] VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 top0.matmul0.matmul_stage_inst.d\[13\] VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__dlygate4sd3_1
X_26835_ clknet_leaf_40_clk_sys _00452_ net682 VGND VGND VPWR VPWR top0.svm0.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold53 top0.matmul0.matmul_stage_inst.d\[10\] VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 top0.matmul0.matmul_stage_inst.b\[6\] VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold75 top0.kpq\[7\] VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13800_ _05586_ _06011_ _06010_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__or3_1
Xhold86 top0.matmul0.matmul_stage_inst.b\[13\] VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 top0.svm0.tB\[9\] VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__dlygate4sd3_1
X_14780_ _06972_ _06980_ VGND VGND VPWR VPWR _06981_ sky130_fd_sc_hd__xnor2_1
X_26766_ clknet_leaf_4_clk_sys _00383_ net580 VGND VGND VPWR VPWR top0.cordic0.cos\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_23978_ _03004_ _03005_ _03022_ _03023_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13731_ _05897_ _05892_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25717_ top0.matmul0.sin\[6\] _04975_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22929_ top0.svm0.counter\[1\] top0.svm0.delta\[1\] VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26697_ clknet_leaf_63_clk_sys _00314_ net647 VGND VGND VPWR VPWR top0.pid_d.prev_error\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16450_ _08537_ _08538_ VGND VGND VPWR VPWR _08539_ sky130_fd_sc_hd__or2b_1
X_13662_ _05863_ _05874_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__nor2_1
X_25648_ net822 _04904_ _04922_ _04924_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15401_ _07491_ _07492_ _07496_ _07499_ VGND VGND VPWR VPWR _07500_ sky130_fd_sc_hd__or4_1
X_13593_ _05805_ net61 _05621_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__and3_1
X_16381_ _08468_ _08469_ _08470_ VGND VGND VPWR VPWR _08471_ sky130_fd_sc_hd__a21o_1
X_25579_ top0.matmul0.a\[12\] top0.matmul0.matmul_stage_inst.e\[12\] _04867_ VGND
+ VGND VPWR VPWR _04877_ sky130_fd_sc_hd__mux2_1
X_18120_ _10103_ _10010_ _10011_ VGND VGND VPWR VPWR _10104_ sky130_fd_sc_hd__o21ai_1
X_15332_ _07418_ _07423_ VGND VGND VPWR VPWR _07431_ sky130_fd_sc_hd__xor2_1
X_18051_ _10024_ _10035_ VGND VGND VPWR VPWR _10036_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27249_ clknet_3_2__leaf_clk_mosi _00863_ VGND VGND VPWR VPWR spi0.data_packed\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_15263_ _07307_ _07361_ VGND VGND VPWR VPWR _07362_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17002_ top0.currT_r\[12\] _09039_ top0.matmul0.beta_pass\[12\] VGND VGND VPWR VPWR
+ _09056_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_50_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14214_ _06421_ _06424_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__xor2_2
XFILLER_0_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15194_ _07286_ _07292_ VGND VGND VPWR VPWR _07293_ sky130_fd_sc_hd__xnor2_4
XANTENNA_6 _05444_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_98_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_98_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_151_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14145_ _06346_ _06356_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14076_ _06286_ _06287_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__nand2_2
X_18953_ _10903_ _10926_ VGND VGND VPWR VPWR _10927_ sky130_fd_sc_hd__and2b_1
X_17904_ _09826_ _09890_ VGND VGND VPWR VPWR _09891_ sky130_fd_sc_hd__xnor2_1
X_18884_ _09863_ _10858_ _09356_ VGND VGND VPWR VPWR _10859_ sky130_fd_sc_hd__a21oi_1
X_17835_ _09817_ _09819_ VGND VGND VPWR VPWR _09822_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17766_ _09751_ _09752_ _09724_ VGND VGND VPWR VPWR _09753_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14978_ _07111_ VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19505_ top0.pid_d.curr_int\[14\] _11289_ _11341_ _11031_ _11396_ VGND VGND VPWR
+ VPWR _00340_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16717_ _08750_ _08800_ VGND VGND VPWR VPWR _08801_ sky130_fd_sc_hd__nand2_1
X_13929_ _06140_ _06141_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17697_ _09662_ _09683_ VGND VGND VPWR VPWR _09684_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19436_ _11334_ _11330_ _10427_ VGND VGND VPWR VPWR _11335_ sky130_fd_sc_hd__o21a_1
X_16648_ _08670_ _08668_ _08733_ VGND VGND VPWR VPWR _08734_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_201_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19367_ top0.pid_d.prev_error\[0\] _11285_ _11288_ net940 VGND VGND VPWR VPWR _00310_
+ sky130_fd_sc_hd__a22o_1
X_16579_ _08664_ _08665_ VGND VGND VPWR VPWR _08666_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18318_ _10183_ _10198_ _10197_ VGND VGND VPWR VPWR _10300_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_143_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19298_ _11236_ _11239_ VGND VGND VPWR VPWR _11240_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_199_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18249_ _10225_ _10231_ VGND VGND VPWR VPWR _10232_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_199_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21260_ _13098_ _13102_ _13053_ VGND VGND VPWR VPWR _13104_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_13_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20211_ _12056_ _12057_ _12058_ _12059_ VGND VGND VPWR VPWR _12060_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_163_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21191_ _12924_ _12140_ _13034_ VGND VGND VPWR VPWR _13035_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_40_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20142_ _11993_ _11996_ _11997_ VGND VGND VPWR VPWR _11998_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24950_ _04285_ _04300_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__xnor2_2
X_20073_ top0.cordic0.slte0.opA\[10\] _11785_ VGND VGND VPWR VPWR _11935_ sky130_fd_sc_hd__nor2_1
X_23901_ _03257_ _03258_ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24881_ _04217_ _04232_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26620_ clknet_leaf_28_clk_sys _00237_ net622 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_23832_ _03186_ _03189_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_170_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23763_ _03063_ _03064_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__or2_1
X_26551_ clknet_leaf_52_clk_sys _00174_ net671 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_20975_ _12072_ _12819_ _12821_ VGND VGND VPWR VPWR _12822_ sky130_fd_sc_hd__o21ai_1
X_25502_ top0.matmul0.matmul_stage_inst.mult1\[7\] _04328_ _04829_ VGND VGND VPWR
+ VPWR _04837_ sky130_fd_sc_hd__mux2_1
X_22714_ _02258_ _02263_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__or2_1
X_23694_ _03048_ _03051_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__xnor2_4
X_26482_ clknet_leaf_89_clk_sys _00113_ net604 VGND VGND VPWR VPWR top0.periodTop\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25433_ _04561_ _04736_ _04775_ _04371_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22645_ _02196_ _02197_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25364_ _04663_ _04708_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22576_ _02130_ _02003_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__or2b_1
XFILLER_0_8_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27103_ clknet_leaf_20_clk_sys _00720_ net609 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.a\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_24315_ _03110_ _03665_ _03669_ VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21527_ net132 net127 VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__nor2b_2
X_25295_ _04562_ _04640_ _04558_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__and3b_1
XFILLER_0_35_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24246_ _03600_ _03601_ _03602_ _03603_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__a211o_1
X_27034_ clknet_leaf_15_clk_sys _00651_ net614 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_16_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21458_ _00964_ _00966_ _01018_ _01011_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_181_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20409_ net289 _12047_ _12251_ _12257_ VGND VGND VPWR VPWR _12258_ sky130_fd_sc_hd__o31a_1
XFILLER_0_31_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24177_ _03478_ _03489_ _03533_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__or3_1
X_21389_ _00954_ _00956_ VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23128_ _02596_ _02619_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__nand2_1
X_23059_ _05541_ _02558_ _02559_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__o21a_1
X_15950_ _08041_ _08044_ VGND VGND VPWR VPWR _08045_ sky130_fd_sc_hd__xnor2_2
X_14901_ spi0.data_packed\[58\] top0.kpq\[10\] _07064_ VGND VGND VPWR VPWR _07071_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15881_ _07965_ _07975_ VGND VGND VPWR VPWR _07977_ sky130_fd_sc_hd__nand2_1
X_17620_ _09605_ _09606_ VGND VGND VPWR VPWR _09607_ sky130_fd_sc_hd__xor2_1
X_14832_ net21 _07030_ VGND VGND VPWR VPWR _07031_ sky130_fd_sc_hd__nand2_1
X_26818_ clknet_leaf_47_clk_sys _00435_ net676 VGND VGND VPWR VPWR top0.svm0.out_valid
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_144_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17551_ _09344_ _09389_ VGND VGND VPWR VPWR _09538_ sky130_fd_sc_hd__xor2_1
X_14763_ _06963_ _06964_ VGND VGND VPWR VPWR _06965_ sky130_fd_sc_hd__xnor2_1
X_26749_ clknet_leaf_92_clk_sys _00366_ net599 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_59_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16502_ _08312_ _08589_ VGND VGND VPWR VPWR _08590_ sky130_fd_sc_hd__xnor2_2
X_13714_ _05913_ _05919_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17482_ net403 net343 VGND VGND VPWR VPWR _09469_ sky130_fd_sc_hd__nand2_1
X_14694_ _06896_ _06897_ VGND VGND VPWR VPWR _06898_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19221_ net439 _11168_ _11169_ VGND VGND VPWR VPWR _11170_ sky130_fd_sc_hd__and3_1
X_16433_ _08429_ _08440_ _08427_ VGND VGND VPWR VPWR _08522_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_39_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13645_ _05799_ _05856_ _05857_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__a21o_1
XFILLER_0_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19152_ net383 _11095_ _11111_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__a21o_1
X_16364_ _08451_ _08453_ VGND VGND VPWR VPWR _08454_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13576_ _05710_ _05712_ _05676_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__o21a_1
X_18103_ _10085_ _10086_ VGND VGND VPWR VPWR _10087_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15315_ _07410_ _07413_ VGND VGND VPWR VPWR _07414_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_87_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19083_ _10790_ net314 net311 _11053_ VGND VGND VPWR VPWR _11055_ sky130_fd_sc_hd__a211o_1
X_16295_ _08283_ _08302_ _08385_ VGND VGND VPWR VPWR _08386_ sky130_fd_sc_hd__o21ai_2
X_18034_ _10017_ _10018_ VGND VGND VPWR VPWR _10019_ sky130_fd_sc_hd__xnor2_1
X_15246_ _07335_ _07336_ VGND VGND VPWR VPWR _07345_ sky130_fd_sc_hd__xor2_2
XFILLER_0_169_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15177_ net493 net508 VGND VGND VPWR VPWR _07276_ sky130_fd_sc_hd__and2_1
X_14128_ _06319_ _06339_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__xnor2_1
X_19985_ _11851_ _11836_ VGND VGND VPWR VPWR _11853_ sky130_fd_sc_hd__nor2_1
X_14059_ _06260_ _06267_ _06270_ _06271_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__a211o_1
X_18936_ top0.pid_d.out\[12\] top0.pid_d.curr_int\[12\] VGND VGND VPWR VPWR _10911_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_24_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_176_Left_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18867_ _10718_ _10716_ _10787_ _10806_ VGND VGND VPWR VPWR _10842_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17818_ _09789_ _09790_ _09803_ VGND VGND VPWR VPWR _09805_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18798_ net374 net314 VGND VGND VPWR VPWR _10774_ sky130_fd_sc_hd__nand2_1
X_17749_ _09734_ _09735_ _09503_ VGND VGND VPWR VPWR _09736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20760_ _12553_ _12608_ VGND VGND VPWR VPWR _12609_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_43_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19419_ _11318_ _11319_ VGND VGND VPWR VPWR _11321_ sky130_fd_sc_hd__nand2_1
XFILLER_0_175_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20691_ _12476_ _12486_ _12488_ VGND VGND VPWR VPWR _12540_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_185_Left_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22430_ _01942_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22361_ _01259_ _01919_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__xor2_1
XFILLER_0_190_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24100_ _03045_ _03046_ _03057_ _03058_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21312_ _13014_ _13153_ VGND VGND VPWR VPWR _13154_ sky130_fd_sc_hd__and2_1
X_25080_ _03900_ _03200_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22292_ net95 net91 VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__or2_2
XFILLER_0_41_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24031_ _02976_ _02977_ _03076_ _03077_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__o22a_2
XFILLER_0_4_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21243_ _12606_ _13086_ _12578_ VGND VGND VPWR VPWR _13087_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21174_ _12987_ _12992_ _13017_ VGND VGND VPWR VPWR _13018_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_194_Left_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20125_ net176 _11981_ net212 VGND VGND VPWR VPWR _11982_ sky130_fd_sc_hd__a21o_1
X_25982_ net1004 _05186_ _05165_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24933_ _04278_ _04283_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__xnor2_1
X_20056_ top0.cordic0.slte0.opA\[8\] _11907_ _11911_ VGND VGND VPWR VPWR _11919_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_175_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24864_ _04071_ _04076_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_46_clk_sys clknet_3_7__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_46_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_26603_ clknet_leaf_54_clk_sys _00226_ net670 VGND VGND VPWR VPWR top0.pid_q.curr_int\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_23815_ _03126_ _03127_ _03125_ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__o21a_1
XFILLER_0_197_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24795_ _04032_ _04144_ _04147_ _04145_ VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__a211o_1
XFILLER_0_185_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26534_ clknet_leaf_61_clk_sys _00157_ net652 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_23746_ net566 net558 top0.matmul0.matmul_stage_inst.e\[12\] VGND VGND VPWR VPWR
+ _03104_ sky130_fd_sc_hd__o21a_2
X_20958_ _12804_ _12805_ VGND VGND VPWR VPWR _12806_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26465_ clknet_leaf_14_clk_sys net563 net617 VGND VGND VPWR VPWR top0.matmul0.done_pass
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_177_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23677_ _03003_ _03034_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__xnor2_4
X_20889_ _12736_ _12737_ VGND VGND VPWR VPWR _12738_ sky130_fd_sc_hd__nor2_2
X_25416_ _04664_ _04756_ _04757_ _04663_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__a2bb2o_1
X_13430_ net65 net63 _05642_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22628_ net211 _02180_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26396_ clknet_leaf_85_clk_sys _00037_ net640 VGND VGND VPWR VPWR top0.kpd\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13361_ _05573_ _05567_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__nor2_1
X_25347_ _03326_ _04630_ _04371_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__o21ai_1
X_22559_ net89 _02031_ _02112_ net79 _02113_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15100_ net522 net475 VGND VGND VPWR VPWR _07199_ sky130_fd_sc_hd__nand2_1
X_13292_ _05504_ _05493_ _05494_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__nor3_1
X_16080_ _08167_ _08172_ VGND VGND VPWR VPWR _08173_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25278_ _04620_ _04623_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27017_ clknet_leaf_16_clk_sys _00634_ net611 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_15031_ top0.pid_d.prev_int\[1\] _07140_ _07144_ top0.pid_d.curr_int\[1\] VGND VGND
+ VPWR VPWR _00118_ sky130_fd_sc_hd__a22o_1
X_24229_ _03563_ _03585_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19770_ _11646_ _11647_ _11652_ net266 VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__o22a_1
X_16982_ net452 _08890_ _09037_ _08930_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__o211a_1
X_18721_ net389 net308 VGND VGND VPWR VPWR _10698_ sky130_fd_sc_hd__nand2_1
X_15933_ net458 net1028 VGND VGND VPWR VPWR _08028_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18652_ _10543_ _10547_ _10541_ VGND VGND VPWR VPWR _10630_ sky130_fd_sc_hd__a21o_1
X_15864_ _07947_ _07958_ VGND VGND VPWR VPWR _07960_ sky130_fd_sc_hd__nand2_1
X_17603_ _09574_ _09579_ VGND VGND VPWR VPWR _09590_ sky130_fd_sc_hd__nor2_1
X_14815_ _05666_ _06867_ net26 VGND VGND VPWR VPWR _07015_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18583_ _10445_ _10462_ _10461_ VGND VGND VPWR VPWR _10562_ sky130_fd_sc_hd__a21oi_2
X_15795_ _07812_ _07891_ VGND VGND VPWR VPWR _07892_ sky130_fd_sc_hd__nor2_1
XFILLER_0_192_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17534_ _09342_ _09520_ VGND VGND VPWR VPWR _09521_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14746_ _06913_ _06937_ _06900_ VGND VGND VPWR VPWR _06948_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_80_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17465_ _09373_ _09442_ _09451_ _09437_ VGND VGND VPWR VPWR _09452_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_74_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14677_ _05640_ _06212_ _06880_ _06832_ net25 VGND VGND VPWR VPWR _06881_ sky130_fd_sc_hd__o32a_1
XFILLER_0_58_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19204_ top0.pid_d.curr_error\[3\] VGND VGND VPWR VPWR _11154_ sky130_fd_sc_hd__inv_2
X_16416_ _08501_ _08504_ VGND VGND VPWR VPWR _08505_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13628_ _05839_ _05840_ net50 _05496_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17396_ _09381_ _09382_ VGND VGND VPWR VPWR _09383_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19135_ top0.kid\[2\] _11098_ _11100_ top0.kpd\[2\] VGND VGND VPWR VPWR _11103_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16347_ _08365_ _08366_ _08367_ VGND VGND VPWR VPWR _08437_ sky130_fd_sc_hd__o21a_1
XFILLER_0_137_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13559_ _05685_ _05691_ _05771_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__o21a_2
XFILLER_0_202_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19066_ _11017_ _11021_ VGND VGND VPWR VPWR _11038_ sky130_fd_sc_hd__nor2_1
X_16278_ _08365_ _08368_ VGND VGND VPWR VPWR _08369_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18017_ _09925_ _09927_ _09923_ VGND VGND VPWR VPWR _10002_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_164_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15229_ _07304_ _07319_ VGND VGND VPWR VPWR _07328_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout107 net108 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout118 net120 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__buf_4
Xfanout129 top0.cordic0.vec\[1\]\[7\] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__buf_4
XFILLER_0_201_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19968_ _11822_ _11829_ VGND VGND VPWR VPWR _11837_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18919_ _10813_ _10814_ _10893_ VGND VGND VPWR VPWR _10894_ sky130_fd_sc_hd__a21oi_1
X_19899_ _11761_ _11762_ _11515_ VGND VGND VPWR VPWR _11773_ sky130_fd_sc_hd__o21ai_1
X_21930_ _01486_ _01491_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21861_ _01399_ _01390_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23600_ top0.matmul0.alpha_pass\[7\] _09290_ net561 VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__mux2_1
X_20812_ _12648_ _12649_ _12660_ VGND VGND VPWR VPWR _12661_ sky130_fd_sc_hd__a21o_1
XFILLER_0_194_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24580_ _03161_ _03908_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__nor2_1
X_21792_ _01265_ _01264_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_194_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20743_ net305 _12491_ VGND VGND VPWR VPWR _12592_ sky130_fd_sc_hd__nand2_1
X_23531_ _02931_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26250_ spi0.data_packed\[23\] spi0.data_packed\[24\] net698 VGND VGND VPWR VPWR
+ _05357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23462_ _02895_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20674_ _12521_ _12522_ net263 VGND VGND VPWR VPWR _12523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25201_ _03280_ _04272_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__nor2_1
X_22413_ _01962_ _01970_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23393_ _11632_ net216 _11715_ _02657_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__o22a_1
X_26181_ _05317_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25132_ _04476_ _04479_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22344_ _01066_ net91 VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25063_ _03355_ _04252_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22275_ net143 _01412_ _01833_ _01834_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__o211a_1
X_24014_ _03359_ _03362_ _03371_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__a21o_1
Xhold150 top0.matmul0.matmul_stage_inst.d\[9\] VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__dlygate4sd3_1
X_21226_ _12627_ _13068_ _12620_ VGND VGND VPWR VPWR _13070_ sky130_fd_sc_hd__mux2_1
Xhold161 top0.svm0.tC\[6\] VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 top0.pid_d.prev_error\[3\] VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 top0.svm0.tA\[4\] VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 top0.svm0.tA\[5\] VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__dlygate4sd3_1
X_21157_ net230 _12925_ _12851_ net225 VGND VGND VPWR VPWR _13002_ sky130_fd_sc_hd__o2bb2a_1
Xfanout630 net2 VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__clkbuf_4
X_20108_ top0.cordic0.slte0.opA\[13\] _11957_ VGND VGND VPWR VPWR _11966_ sky130_fd_sc_hd__and2_1
Xfanout641 net645 VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__clkbuf_4
Xfanout652 net653 VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__buf_2
X_25965_ top0.matmul0.beta_pass\[1\] _05169_ _05173_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__a21o_1
Xfanout663 net687 VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__clkbuf_4
X_21088_ _12897_ _12933_ VGND VGND VPWR VPWR _12934_ sky130_fd_sc_hd__xnor2_1
Xfanout674 net675 VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__clkbuf_2
Xfanout685 net686 VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__buf_2
XFILLER_0_176_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24916_ _04264_ _04266_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__xnor2_2
X_20039_ _11518_ _11877_ VGND VGND VPWR VPWR _11903_ sky130_fd_sc_hd__or2_1
Xfanout696 net700 VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__buf_2
X_25896_ _05104_ _05102_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__or2b_1
XFILLER_0_38_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24847_ _03325_ _03900_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__nor2_2
XFILLER_0_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14600_ _06697_ _06792_ _06745_ _06740_ VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__or4b_1
X_15580_ _07590_ _07678_ _07281_ VGND VGND VPWR VPWR _07679_ sky130_fd_sc_hd__mux2_1
X_24778_ _03743_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_185_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14531_ _06727_ _06735_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__nor2_1
XFILLER_0_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26517_ clknet_leaf_68_clk_sys _00140_ net659 VGND VGND VPWR VPWR top0.pid_q.out\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_23729_ _03035_ _03086_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__xor2_4
XFILLER_0_200_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17250_ _09252_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14462_ _06667_ _06668_ _06669_ VGND VGND VPWR VPWR _06670_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26448_ clknet_leaf_60_clk_sys _00089_ net651 VGND VGND VPWR VPWR top0.kiq\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16201_ _07493_ _08170_ net468 VGND VGND VPWR VPWR _08293_ sky130_fd_sc_hd__a21oi_1
X_13413_ _05625_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17181_ _09191_ VGND VGND VPWR VPWR _09192_ sky130_fd_sc_hd__buf_2
X_14393_ _06594_ _06601_ VGND VGND VPWR VPWR _06602_ sky130_fd_sc_hd__xnor2_1
X_26379_ clknet_leaf_43_clk_sys _00020_ net682 VGND VGND VPWR VPWR top0.svm0.tC\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16132_ _08217_ _08224_ VGND VGND VPWR VPWR _08225_ sky130_fd_sc_hd__xor2_2
X_13344_ _05548_ _05556_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16063_ _08088_ _08156_ VGND VGND VPWR VPWR _08157_ sky130_fd_sc_hd__xnor2_1
X_13275_ top0.matmul0.alpha_pass\[1\] _05435_ _05474_ VGND VGND VPWR VPWR _05488_
+ sky130_fd_sc_hd__nand3_2
X_15014_ _07132_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_184_Right_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19822_ _11448_ _11558_ net82 VGND VGND VPWR VPWR _11701_ sky130_fd_sc_hd__o21a_1
X_16965_ _09019_ _09020_ VGND VGND VPWR VPWR _09022_ sky130_fd_sc_hd__or2_1
X_19753_ net128 net123 net111 net107 net199 net187 VGND VGND VPWR VPWR _11636_ sky130_fd_sc_hd__mux4_1
XFILLER_0_194_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15916_ _07932_ _07942_ _07937_ VGND VGND VPWR VPWR _08011_ sky130_fd_sc_hd__a21bo_1
X_18704_ _05449_ _10681_ VGND VGND VPWR VPWR _10682_ sky130_fd_sc_hd__and2_1
X_19684_ _11550_ _11569_ _11570_ VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__a21oi_1
X_16896_ top0.currT_r\[5\] _08946_ top0.matmul0.beta_pass\[5\] VGND VGND VPWR VPWR
+ _08957_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_189_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18635_ net377 net364 _10611_ _10612_ _09364_ VGND VGND VPWR VPWR _10613_ sky130_fd_sc_hd__a32o_1
X_15847_ _07937_ _07942_ VGND VGND VPWR VPWR _07943_ sky130_fd_sc_hd__xor2_1
XFILLER_0_189_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18566_ net334 net338 VGND VGND VPWR VPWR _10545_ sky130_fd_sc_hd__xor2_4
XFILLER_0_115_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15778_ net443 _07874_ VGND VGND VPWR VPWR _07875_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17517_ _09492_ _09503_ VGND VGND VPWR VPWR _09504_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14729_ net31 _05626_ _06929_ _06930_ _06931_ VGND VGND VPWR VPWR _06932_ sky130_fd_sc_hd__a311o_1
XFILLER_0_75_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18497_ _10471_ _10476_ VGND VGND VPWR VPWR _10477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17448_ net398 _09395_ _09434_ net400 VGND VGND VPWR VPWR _09435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17379_ _09364_ _09365_ VGND VGND VPWR VPWR _09366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19118_ top0.pid_d.out\[15\] _09339_ _11087_ _11089_ net1019 VGND VGND VPWR VPWR
+ _11090_ sky130_fd_sc_hd__o221a_1
XFILLER_0_43_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20390_ _12237_ _12238_ VGND VGND VPWR VPWR _12239_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19049_ _11017_ _11021_ VGND VGND VPWR VPWR _11022_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22060_ _01549_ _01553_ _01552_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21011_ _12849_ _12857_ VGND VGND VPWR VPWR _12858_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25750_ net70 top0.matmul0.cos\[3\] _05458_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__and3_1
X_22962_ _02466_ _02468_ _02331_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__o21a_1
X_24701_ _03937_ _03938_ _03944_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__and3_1
X_21913_ _01457_ _01461_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__nand2_1
X_25681_ net825 _04904_ _04936_ _04950_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__a22o_1
X_22893_ _02352_ top0.svm0.tC\[1\] top0.svm0.tC\[2\] _02347_ _02410_ VGND VGND VPWR
+ VPWR _02411_ sky130_fd_sc_hd__a221o_1
X_24632_ _02985_ _02987_ _03150_ _03151_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__o22a_1
XFILLER_0_195_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21844_ _01376_ _01404_ _01405_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24563_ _03794_ _03789_ _03788_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_33_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21775_ _01331_ _01336_ _01332_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26302_ spi0.data_packed\[49\] spi0.data_packed\[50\] net697 VGND VGND VPWR VPWR
+ _05383_ sky130_fd_sc_hd__mux2_1
X_20726_ _12549_ _12566_ _12571_ _12573_ _12574_ VGND VGND VPWR VPWR _12575_ sky130_fd_sc_hd__a221o_2
X_23514_ _02922_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__clkbuf_1
X_27282_ clknet_3_3__leaf_clk_mosi _00896_ VGND VGND VPWR VPWR spi0.data_packed\[68\]
+ sky130_fd_sc_hd__dfxtp_1
X_24494_ _03663_ _03849_ _03751_ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26233_ _05348_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20657_ net270 net287 VGND VGND VPWR VPWR _12506_ sky130_fd_sc_hd__or2b_1
XFILLER_0_74_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23445_ _02878_ _02880_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23376_ _02815_ _02817_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__nand2_1
X_26164_ net18 _05303_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20588_ net264 net253 VGND VGND VPWR VPWR _12437_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25115_ _04386_ _04463_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__xnor2_1
X_22327_ _01742_ _01745_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__xor2_1
XFILLER_0_104_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26095_ _05273_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25046_ _04303_ _04393_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__nor2_1
X_22258_ _01755_ _01815_ _01817_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_40_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21209_ _13044_ _13052_ VGND VGND VPWR VPWR _13053_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22189_ _01089_ _01456_ _01708_ _01144_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__o2bb2a_1
X_26997_ clknet_leaf_24_clk_sys _00614_ net625 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout460 top0.pid_q.mult0.b\[9\] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__buf_4
Xfanout471 top0.pid_q.mult0.b\[5\] VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__clkbuf_4
X_16750_ _08526_ _08753_ VGND VGND VPWR VPWR _08834_ sky130_fd_sc_hd__nor2_1
Xfanout482 net483 VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__clkbuf_2
X_13962_ _06171_ _06172_ _06174_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__o21bai_1
X_25948_ _05154_ _05157_ _05160_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__mux2_1
Xfanout493 net495 VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__clkbuf_4
X_15701_ net549 _07795_ _07798_ net544 _07705_ VGND VGND VPWR VPWR _07799_ sky130_fd_sc_hd__a221o_1
XFILLER_0_198_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16681_ net449 _08696_ VGND VGND VPWR VPWR _08766_ sky130_fd_sc_hd__and2_1
X_13893_ net30 VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__inv_2
X_25879_ _05094_ _05097_ _05088_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__mux2_1
X_18420_ _10266_ _10268_ _10256_ VGND VGND VPWR VPWR _10401_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_115_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15632_ _07726_ _07729_ VGND VGND VPWR VPWR _07730_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18351_ _10252_ _10332_ VGND VGND VPWR VPWR _10333_ sky130_fd_sc_hd__xnor2_1
X_15563_ _07563_ _07661_ _07549_ VGND VGND VPWR VPWR _07662_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17302_ top0.matmul0.beta_pass\[8\] _09296_ net562 VGND VGND VPWR VPWR _09297_ sky130_fd_sc_hd__mux2_1
X_14514_ _05579_ _06585_ net23 VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18282_ net411 net310 VGND VGND VPWR VPWR _10264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15494_ _07589_ _07592_ VGND VGND VPWR VPWR _07593_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17233_ top0.pid_q.prev_int\[13\] _09231_ top0.pid_q.curr_int\[13\] VGND VGND VPWR
+ VPWR _09238_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14445_ _06574_ _06579_ _06576_ VGND VGND VPWR VPWR _06653_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17164_ top0.pid_q.prev_int\[5\] _09172_ top0.pid_q.curr_int\[5\] VGND VGND VPWR
+ VPWR _09177_ sky130_fd_sc_hd__a21o_1
X_14376_ net30 _05588_ VGND VGND VPWR VPWR _06585_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16115_ _08109_ _08111_ _08110_ VGND VGND VPWR VPWR _08208_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13327_ _05536_ _05538_ _05539_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__nor3_1
XFILLER_0_12_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17095_ top0.pid_q.curr_error\[6\] _00011_ _09117_ VGND VGND VPWR VPWR _09124_ sky130_fd_sc_hd__and3_1
XFILLER_0_161_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16046_ _08040_ _08138_ _08139_ VGND VGND VPWR VPWR _08140_ sky130_fd_sc_hd__o21a_1
XFILLER_0_177_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13258_ top0.matmul0.beta_pass\[5\] _05466_ _05470_ _05464_ top0.c_out_calc\[5\]
+ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__a32o_1
XFILLER_0_86_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13189_ top0.matmul0.matmul_stage_inst.start VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19805_ _11684_ _11685_ VGND VGND VPWR VPWR _11686_ sky130_fd_sc_hd__nor2_1
X_17997_ top0.pid_d.out\[1\] top0.pid_d.curr_int\[1\] VGND VGND VPWR VPWR _09982_
+ sky130_fd_sc_hd__or2_1
X_16948_ top0.pid_q.prev_error\[9\] top0.pid_q.curr_error\[9\] VGND VGND VPWR VPWR
+ _09006_ sky130_fd_sc_hd__xnor2_1
X_19736_ _11619_ VGND VGND VPWR VPWR _11620_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16879_ _08941_ VGND VGND VPWR VPWR _08942_ sky130_fd_sc_hd__inv_2
X_19667_ net111 net108 net199 VGND VGND VPWR VPWR _11554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18618_ _10594_ _10514_ _10595_ VGND VGND VPWR VPWR _10596_ sky130_fd_sc_hd__a21o_1
X_19598_ top0.cordic0.slte0.opB\[6\] top0.cordic0.slte0.opA\[6\] VGND VGND VPWR VPWR
+ _11487_ sky130_fd_sc_hd__and2b_1
XFILLER_0_176_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18549_ _10526_ _10527_ VGND VGND VPWR VPWR _10528_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21560_ net122 VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20511_ _12268_ _12270_ _12275_ VGND VGND VPWR VPWR _12360_ sky130_fd_sc_hd__or3_2
XFILLER_0_129_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21491_ _01024_ _01049_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23230_ _02679_ _01320_ _02659_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__or3b_1
XFILLER_0_71_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20442_ _12059_ net281 _12057_ _12290_ VGND VGND VPWR VPWR _12291_ sky130_fd_sc_hd__and4b_1
XFILLER_0_160_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23161_ _02644_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20373_ net283 _12127_ _12128_ VGND VGND VPWR VPWR _12222_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22112_ _01406_ _01318_ _01608_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__and3_1
X_23092_ _02548_ _02549_ _02556_ _02563_ _02592_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_3_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22043_ _01599_ _01604_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__or2_1
X_26920_ clknet_leaf_0_clk_sys _00537_ net578 VGND VGND VPWR VPWR top0.matmul0.sin\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_26851_ clknet_leaf_47_clk_sys _00468_ net676 VGND VGND VPWR VPWR top0.svm0.delta\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25802_ _02282_ _12014_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__nor2_1
XFILLER_0_177_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26782_ clknet_leaf_110_clk_sys _00399_ net579 VGND VGND VPWR VPWR top0.cordic0.sin\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_23994_ _03336_ _03339_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25733_ net891 _04890_ _04913_ _04986_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22945_ top0.svm0.delta\[4\] VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25664_ top0.matmul0.sin\[7\] _04937_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__xor2_1
X_22876_ top0.svm0.tB\[9\] _02394_ _02360_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__o21a_1
XFILLER_0_167_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24615_ _03907_ _03913_ _03905_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__a21o_1
X_21827_ _01386_ _01388_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__nor2b_1
X_25595_ _04886_ top0.matmul0.cos\[1\] _04878_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__or3_1
XFILLER_0_39_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24546_ _03765_ _03900_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__nor2_1
X_21758_ _01319_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_202_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20709_ net292 net278 net261 VGND VGND VPWR VPWR _12558_ sky130_fd_sc_hd__and3_1
X_27265_ clknet_3_6__leaf_clk_mosi _00879_ VGND VGND VPWR VPWR spi0.data_packed\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_24477_ _03821_ _03832_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21689_ _01130_ _01249_ _01162_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__a21o_1
X_14230_ _06046_ _06426_ VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26216_ spi0.data_packed\[6\] spi0.data_packed\[7\] net694 VGND VGND VPWR VPWR _05340_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23428_ net215 _11760_ _02712_ _11730_ VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__a22o_1
X_27196_ clknet_leaf_57_clk_sys _00810_ net664 VGND VGND VPWR VPWR top0.currT_r\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_184_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14161_ _06266_ VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26147_ _05290_ top0.cordic0.slte0.opB\[4\] _12006_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23359_ _02800_ _02791_ _02801_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__a21oi_1
X_14092_ _06233_ _06236_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__nand2_1
X_26078_ top0.a_in_matmul\[11\] _05260_ _05230_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25029_ _04287_ _04299_ _04378_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__o21a_1
X_17920_ _09904_ _09905_ VGND VGND VPWR VPWR _09906_ sky130_fd_sc_hd__xnor2_1
X_17851_ _09834_ _09837_ VGND VGND VPWR VPWR _09838_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16802_ net512 _08855_ _08858_ net796 _08874_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__a221o_1
X_17782_ _09677_ _09680_ VGND VGND VPWR VPWR _09769_ sky130_fd_sc_hd__nand2_1
X_14994_ spi0.data_packed\[3\] top0.periodTop\[3\] _07108_ VGND VGND VPWR VPWR _07122_
+ sky130_fd_sc_hd__mux2_1
Xfanout290 net293 VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkbuf_4
X_16733_ net498 _08816_ VGND VGND VPWR VPWR _08817_ sky130_fd_sc_hd__nand2_1
X_19521_ net183 net189 VGND VGND VPWR VPWR _11411_ sky130_fd_sc_hd__nor2_1
X_13945_ _05734_ _05740_ _05730_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_159_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_94_clk_sys clknet_3_0__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_94_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_19452_ top0.pid_d.curr_int\[8\] _11289_ _11292_ _11349_ VGND VGND VPWR VPWR _11350_
+ sky130_fd_sc_hd__a22o_1
X_16664_ _08717_ _08722_ _08748_ VGND VGND VPWR VPWR _08749_ sky130_fd_sc_hd__a21o_1
X_13876_ _05765_ _05766_ net42 _05472_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18403_ net368 VGND VGND VPWR VPWR _10384_ sky130_fd_sc_hd__inv_2
X_15615_ _07585_ _07683_ VGND VGND VPWR VPWR _07713_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19383_ top0.pid_d.state\[0\] top0.pid_d.state\[3\] net433 _05441_ VGND VGND VPWR
+ VPWR _11289_ sky130_fd_sc_hd__o31a_4
X_16595_ _08601_ _08678_ VGND VGND VPWR VPWR _08682_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18334_ _10308_ _10315_ VGND VGND VPWR VPWR _10316_ sky130_fd_sc_hd__xnor2_2
X_15546_ _07565_ _07566_ _07567_ VGND VGND VPWR VPWR _07645_ sky130_fd_sc_hd__o21a_1
XFILLER_0_189_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_7_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18265_ top0.pid_d.out\[5\] top0.pid_d.curr_int\[5\] VGND VGND VPWR VPWR _10247_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15477_ net535 net457 VGND VGND VPWR VPWR _07576_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17216_ top0.pid_q.curr_int\[11\] top0.pid_q.prev_int\[11\] VGND VGND VPWR VPWR _09223_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14428_ _06629_ _06635_ VGND VGND VPWR VPWR _06636_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_181_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18196_ _10175_ _10178_ VGND VGND VPWR VPWR _10179_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17147_ top0.pid_q.curr_int\[3\] _09141_ _09162_ _09136_ VGND VGND VPWR VPWR _00216_
+ sky130_fd_sc_hd__a22o_1
X_14359_ net39 _05605_ VGND VGND VPWR VPWR _06568_ sky130_fd_sc_hd__nand2_2
XFILLER_0_188_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout9 _11651_ VGND VGND VPWR VPWR net1020 sky130_fd_sc_hd__buf_4
XFILLER_0_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17078_ _00008_ _08855_ VGND VGND VPWR VPWR _09113_ sky130_fd_sc_hd__or2_1
X_16029_ _08042_ _08043_ _08122_ VGND VGND VPWR VPWR _08123_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19719_ _11584_ _11588_ _11603_ VGND VGND VPWR VPWR _11604_ sky130_fd_sc_hd__o21bai_2
X_20991_ _12776_ _12837_ VGND VGND VPWR VPWR _12838_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22730_ top0.cordic0.sin\[12\] _12004_ _12036_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22661_ _02159_ _02199_ _02154_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__a21o_1
XFILLER_0_177_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24400_ top0.matmul0.matmul_stage_inst.mult2\[1\] _03756_ _03642_ VGND VGND VPWR
+ VPWR _03757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21612_ _01083_ _01173_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__xnor2_4
X_25380_ _04288_ _04182_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22592_ net95 _01980_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24331_ _03572_ _03687_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__nand2_2
XFILLER_0_168_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21543_ net133 VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27050_ clknet_leaf_22_clk_sys _00667_ net607 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.d\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_24262_ _03439_ _03440_ _03619_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__o21a_1
X_21474_ _12968_ _01037_ _01038_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__and3_1
X_26001_ top0.b_in_matmul\[9\] _05201_ _05196_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__mux2_1
X_20425_ net281 net274 VGND VGND VPWR VPWR _12274_ sky130_fd_sc_hd__nor2_1
X_23213_ net254 net250 net244 net243 net198 net192 VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__mux4_2
XFILLER_0_160_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24193_ _03542_ _03543_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23144_ top0.svm0.delta\[13\] _02628_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__or2_1
X_20356_ _12198_ _12200_ _12203_ VGND VGND VPWR VPWR _12205_ sky130_fd_sc_hd__nand3_1
XFILLER_0_141_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23075_ top0.svm0.counter\[0\] _05805_ _02574_ _02575_ VGND VGND VPWR VPWR _02576_
+ sky130_fd_sc_hd__or4_1
X_20287_ net234 net226 VGND VGND VPWR VPWR _12136_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22026_ _01574_ _01576_ _01577_ _01587_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__o31a_1
X_26903_ clknet_leaf_4_clk_sys _00520_ net580 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold10 top0.kpq\[12\] VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 top0.cordic0.sin\[1\] VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 top0.cordic0.cos\[0\] VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__dlygate4sd3_1
X_26834_ clknet_leaf_43_clk_sys _00451_ net682 VGND VGND VPWR VPWR top0.svm0.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold43 top0.c_out_calc\[5\] VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold54 top0.periodTop\[14\] VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 top0.pid_d.curr_error\[14\] VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 top0.svm0.tB\[7\] VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 top0.kpq\[2\] VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26765_ clknet_leaf_87_clk_sys _00382_ net642 VGND VGND VPWR VPWR top0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold98 top0.c_out_calc\[2\] VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__dlygate4sd3_1
X_23977_ _03330_ _03334_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_187_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13730_ _05936_ _05941_ _05942_ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__a21o_1
X_25716_ net73 _04926_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__nand2_1
X_22928_ top0.svm0.delta\[2\] VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__inv_2
X_26696_ clknet_leaf_64_clk_sys _00313_ net656 VGND VGND VPWR VPWR top0.pid_d.prev_error\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13661_ _05865_ _05868_ _05873_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__a21oi_2
X_25647_ net72 _04923_ _04890_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__a21oi_1
X_22859_ _02321_ _02373_ _02378_ _02315_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15400_ _07497_ _07498_ _07440_ VGND VGND VPWR VPWR _07499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16380_ _08383_ _08381_ VGND VGND VPWR VPWR _08470_ sky130_fd_sc_hd__nor2_1
X_13592_ net65 VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__inv_2
X_25578_ _04876_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15331_ _07427_ _07429_ VGND VGND VPWR VPWR _07430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24529_ _02979_ _02980_ _03069_ _03071_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__o22a_2
XFILLER_0_136_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18050_ _10029_ _10034_ VGND VGND VPWR VPWR _10035_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27248_ clknet_3_2__leaf_clk_mosi _00862_ VGND VGND VPWR VPWR spi0.data_packed\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_15262_ _07305_ _07306_ VGND VGND VPWR VPWR _07361_ sky130_fd_sc_hd__xor2_1
XFILLER_0_108_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17001_ _09053_ _09054_ VGND VGND VPWR VPWR _09055_ sky130_fd_sc_hd__xnor2_1
X_14213_ _06422_ _06423_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__xor2_1
XFILLER_0_112_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27179_ clknet_leaf_57_clk_sys _00793_ net643 VGND VGND VPWR VPWR top0.periodTop_r\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_15193_ _07288_ _07291_ VGND VGND VPWR VPWR _07292_ sky130_fd_sc_hd__xnor2_2
XANTENNA_7 net1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14144_ _06348_ _06355_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__xor2_2
XFILLER_0_120_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_89_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14075_ net48 _05605_ _06184_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__a21o_1
X_18952_ _10923_ _10925_ _10904_ VGND VGND VPWR VPWR _10926_ sky130_fd_sc_hd__a21o_1
X_17903_ _09883_ _09889_ VGND VGND VPWR VPWR _09890_ sky130_fd_sc_hd__xnor2_1
X_18883_ _09395_ _10781_ VGND VGND VPWR VPWR _10858_ sky130_fd_sc_hd__nand2_1
X_17834_ _09747_ _09750_ _09753_ _09820_ VGND VGND VPWR VPWR _09821_ sky130_fd_sc_hd__o31a_1
XFILLER_0_83_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14977_ spi0.data_packed\[30\] top0.kiq\[14\] _07108_ VGND VGND VPWR VPWR _07111_
+ sky130_fd_sc_hd__mux2_1
X_17765_ _09716_ _09717_ _09738_ _09743_ VGND VGND VPWR VPWR _09752_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19504_ _11261_ _11395_ _11388_ VGND VGND VPWR VPWR _11396_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13928_ net48 _05639_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__nand2_2
X_16716_ _08757_ _08754_ _08776_ VGND VGND VPWR VPWR _08800_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17696_ _09669_ _09682_ VGND VGND VPWR VPWR _09683_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16647_ _08670_ _08668_ _08671_ VGND VGND VPWR VPWR _08733_ sky130_fd_sc_hd__a21bo_1
X_19435_ top0.pid_d.prev_int\[6\] VGND VGND VPWR VPWR _11334_ sky130_fd_sc_hd__inv_2
XFILLER_0_202_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13859_ _06022_ _06070_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16578_ _08312_ _08663_ VGND VGND VPWR VPWR _08665_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19366_ _11287_ VGND VGND VPWR VPWR _11288_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18317_ _10286_ _10298_ VGND VGND VPWR VPWR _10299_ sky130_fd_sc_hd__xnor2_1
X_15529_ _07624_ _07627_ VGND VGND VPWR VPWR _07628_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19297_ _11227_ _11237_ _11238_ VGND VGND VPWR VPWR _11239_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18248_ _10141_ _10230_ VGND VGND VPWR VPWR _10231_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18179_ _10154_ VGND VGND VPWR VPWR _10162_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20210_ net290 net296 VGND VGND VPWR VPWR _12059_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_25_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21190_ net230 _12819_ net226 VGND VGND VPWR VPWR _13034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20141_ _11433_ net180 VGND VGND VPWR VPWR _11997_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20072_ net1014 _11933_ net177 VGND VGND VPWR VPWR _11934_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23900_ _03065_ _03072_ VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__xnor2_2
X_24880_ _04226_ _04231_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__xnor2_1
X_23831_ _03187_ _03188_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_197_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26550_ clknet_leaf_50_clk_sys _00173_ net675 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_178_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23762_ _03088_ _03089_ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__or2_4
XFILLER_0_170_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20974_ net222 net213 _12820_ VGND VGND VPWR VPWR _12821_ sky130_fd_sc_hd__or3_1
X_25501_ _04836_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22713_ _02186_ _02263_ _02172_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__o21a_1
X_26481_ clknet_leaf_89_clk_sys _00112_ net603 VGND VGND VPWR VPWR top0.periodTop\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_23693_ _03049_ _03050_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25432_ _03363_ _04437_ _04736_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22644_ _02194_ _02195_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__nand2_1
XFILLER_0_192_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25363_ _04702_ _04707_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22575_ _02128_ _02129_ _02083_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__mux2_1
X_27102_ clknet_leaf_20_clk_sys _00719_ net610 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.a\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24314_ _03665_ _03666_ _03668_ _03670_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21526_ net159 net139 VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__xor2_4
X_25294_ _03112_ _04174_ _04561_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__or3b_1
XFILLER_0_69_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_42_clk_sys clknet_3_7__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_42_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_27033_ clknet_leaf_18_clk_sys _00650_ net614 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_24245_ _03555_ _03557_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__and2_1
X_21457_ _00964_ _01020_ _01021_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__o21ai_2
X_20408_ net269 _12254_ _12256_ _11571_ _12050_ VGND VGND VPWR VPWR _12257_ sky130_fd_sc_hd__a221o_2
X_24176_ _03478_ _03489_ _03533_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__o21a_1
X_21388_ _13159_ _13184_ _00955_ VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__a21o_2
X_23127_ top0.svm0.delta\[7\] top0.svm0.delta\[8\] top0.svm0.delta\[9\] _02612_ VGND
+ VGND VPWR VPWR _02619_ sky130_fd_sc_hd__or4_1
X_20339_ _12164_ _12176_ _12178_ VGND VGND VPWR VPWR _12188_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23058_ net52 top0.svm0.counter\[5\] _02557_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__or3_1
X_14900_ _07070_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__clkbuf_1
X_22009_ net163 _01266_ net136 VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__or3_1
X_15880_ _07965_ _07975_ VGND VGND VPWR VPWR _07976_ sky130_fd_sc_hd__nor2_1
X_14831_ _07029_ _06867_ _06975_ VGND VGND VPWR VPWR _07030_ sky130_fd_sc_hd__mux2_1
X_26817_ clknet_leaf_60_clk_sys net773 net652 VGND VGND VPWR VPWR top0.pid_q.prev_int\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17550_ _09528_ _09536_ VGND VGND VPWR VPWR _09537_ sky130_fd_sc_hd__xor2_2
X_14762_ net34 _06867_ VGND VGND VPWR VPWR _06964_ sky130_fd_sc_hd__nand2_1
X_26748_ clknet_leaf_97_clk_sys _00365_ net588 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_16501_ _08453_ _08525_ _08526_ VGND VGND VPWR VPWR _08589_ sky130_fd_sc_hd__o21ba_1
X_13713_ _05886_ _05925_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17481_ net408 net340 VGND VGND VPWR VPWR _09468_ sky130_fd_sc_hd__and2_1
X_14693_ _06893_ _06895_ VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26679_ clknet_leaf_64_clk_sys _00296_ net656 VGND VGND VPWR VPWR top0.pid_d.curr_error\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_169_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16432_ _08507_ _08520_ VGND VGND VPWR VPWR _08521_ sky130_fd_sc_hd__xnor2_2
X_19220_ _11166_ _11167_ VGND VGND VPWR VPWR _11169_ sky130_fd_sc_hd__or2_1
X_13644_ _05716_ _05798_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19151_ top0.kid\[10\] _11097_ _11099_ top0.kpd\[10\] VGND VGND VPWR VPWR _11111_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16363_ _08452_ VGND VGND VPWR VPWR _08453_ sky130_fd_sc_hd__buf_2
XFILLER_0_27_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13575_ _05786_ _05787_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18102_ _10079_ _10084_ VGND VGND VPWR VPWR _10086_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15314_ _07411_ _07412_ VGND VGND VPWR VPWR _07413_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19082_ net311 net370 _11004_ _11053_ net365 VGND VGND VPWR VPWR _11054_ sky130_fd_sc_hd__o32a_1
XFILLER_0_87_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16294_ _08283_ _08302_ _08285_ VGND VGND VPWR VPWR _08385_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_13_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18033_ net332 net393 VGND VGND VPWR VPWR _10018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15245_ _07304_ _07319_ VGND VGND VPWR VPWR _07344_ sky130_fd_sc_hd__xor2_2
XFILLER_0_151_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_97_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15176_ net514 net485 VGND VGND VPWR VPWR _07275_ sky130_fd_sc_hd__nand2_1
X_14127_ _06328_ _06338_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19984_ _11851_ _11836_ VGND VGND VPWR VPWR _11852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14058_ _06263_ _06269_ _06258_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__and3b_1
X_18935_ top0.pid_d.out\[12\] top0.pid_d.curr_int\[12\] VGND VGND VPWR VPWR _10910_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_94_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18866_ _10751_ _10840_ _10752_ VGND VGND VPWR VPWR _10841_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17817_ _09789_ _09790_ _09803_ VGND VGND VPWR VPWR _09804_ sky130_fd_sc_hd__and3_1
XFILLER_0_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18797_ net377 net311 VGND VGND VPWR VPWR _10773_ sky130_fd_sc_hd__nand2_1
X_17748_ _09508_ _09509_ VGND VGND VPWR VPWR _09735_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17679_ net322 net420 VGND VGND VPWR VPWR _09666_ sky130_fd_sc_hd__and2_1
X_19418_ _11318_ _11319_ VGND VGND VPWR VPWR _11320_ sky130_fd_sc_hd__or2_1
X_20690_ _12446_ _12455_ _12537_ _12538_ VGND VGND VPWR VPWR _12539_ sky130_fd_sc_hd__a31o_1
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19349_ _05443_ _11120_ _11276_ VGND VGND VPWR VPWR _11280_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22360_ _01143_ _01918_ net134 VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_198_Right_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21311_ _13144_ _13152_ _13142_ VGND VGND VPWR VPWR _13153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22291_ net99 _01820_ _01849_ _01850_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24030_ _02985_ _02987_ _03063_ _03064_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__o22a_1
X_21242_ _12583_ _12605_ _13085_ VGND VGND VPWR VPWR _13086_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_5_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold310 top0.cordic0.sin\[3\] VGND VGND VPWR VPWR net1010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21173_ _12987_ _12992_ _12980_ VGND VGND VPWR VPWR _13017_ sky130_fd_sc_hd__o21a_1
XFILLER_0_159_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20124_ _11936_ _11978_ VGND VGND VPWR VPWR _11981_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25981_ top0.matmul0.beta_pass\[5\] _05169_ _05185_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__a21o_1
X_24932_ _04279_ _04282_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__xnor2_2
X_20055_ _11915_ _11917_ _11426_ VGND VGND VPWR VPWR _11918_ sky130_fd_sc_hd__o21a_1
X_24863_ _04071_ _04076_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26602_ clknet_leaf_51_clk_sys _00225_ net670 VGND VGND VPWR VPWR top0.pid_q.curr_int\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_198_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23814_ _03125_ _03126_ _03127_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__or3_1
X_24794_ _04035_ _04143_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26533_ clknet_leaf_61_clk_sys _00156_ net651 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_23745_ net571 net575 top0.matmul0.matmul_stage_inst.f\[12\] VGND VGND VPWR VPWR
+ _03103_ sky130_fd_sc_hd__o21a_2
XFILLER_0_200_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20957_ _12677_ _12728_ _12727_ VGND VGND VPWR VPWR _12805_ sky130_fd_sc_hd__a21o_1
XFILLER_0_191_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26464_ clknet_leaf_17_clk_sys net567 net612 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23676_ _03014_ _03033_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20888_ _12730_ _12735_ VGND VGND VPWR VPWR _12737_ sky130_fd_sc_hd__and2_1
XFILLER_0_165_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25415_ _04663_ _04757_ _04758_ _04661_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__o211a_1
X_22627_ _02175_ _02176_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__or2_2
X_26395_ clknet_leaf_85_clk_sys _00036_ net640 VGND VGND VPWR VPWR top0.kpd\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25346_ _04626_ _04636_ _04635_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__a21o_1
X_13360_ net46 VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__inv_2
X_22558_ net107 net100 _01924_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_165_Right_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21509_ net126 VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__inv_2
X_25277_ _04621_ _04622_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__xor2_1
X_13291_ net40 VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__inv_1
XFILLER_0_51_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22489_ _02007_ _02045_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__xnor2_1
X_27016_ clknet_leaf_16_clk_sys _00633_ net613 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_122_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15030_ net968 _07140_ _07144_ top0.pid_d.curr_int\[0\] VGND VGND VPWR VPWR _00117_
+ sky130_fd_sc_hd__a22o_1
X_24228_ _03563_ _03585_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24159_ _03468_ _03470_ _03483_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_20_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16981_ net552 _09029_ _09036_ top0.pid_q.state\[3\] _08881_ VGND VGND VPWR VPWR
+ _09037_ sky130_fd_sc_hd__a221o_1
X_18720_ _10695_ _10696_ VGND VGND VPWR VPWR _10697_ sky130_fd_sc_hd__xor2_1
X_15932_ net467 net1029 VGND VGND VPWR VPWR _08027_ sky130_fd_sc_hd__nand2_2
XFILLER_0_155_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18651_ _10610_ _10628_ VGND VGND VPWR VPWR _10629_ sky130_fd_sc_hd__xor2_2
X_15863_ _07947_ _07958_ VGND VGND VPWR VPWR _07959_ sky130_fd_sc_hd__nor2_1
XFILLER_0_188_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14814_ net21 _06824_ VGND VGND VPWR VPWR _07014_ sky130_fd_sc_hd__and2_1
X_17602_ net425 _09584_ _09582_ VGND VGND VPWR VPWR _09589_ sky130_fd_sc_hd__a21o_1
X_18582_ _10464_ _10488_ _10560_ VGND VGND VPWR VPWR _10561_ sky130_fd_sc_hd__a21o_1
X_15794_ _07882_ _07890_ VGND VGND VPWR VPWR _07891_ sky130_fd_sc_hd__xnor2_1
X_14745_ _06942_ _06946_ VGND VGND VPWR VPWR _06947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17533_ _09340_ _09341_ VGND VGND VPWR VPWR _09520_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17464_ _09427_ _09440_ _09439_ VGND VGND VPWR VPWR _09451_ sky130_fd_sc_hd__o21a_1
X_14676_ _05626_ _06832_ VGND VGND VPWR VPWR _06880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16415_ _08502_ _08503_ VGND VGND VPWR VPWR _08504_ sky130_fd_sc_hd__xnor2_1
X_19203_ _11125_ _11149_ _11152_ _11153_ _07800_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__o311a_1
XFILLER_0_200_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13627_ net43 _05484_ _05486_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17395_ net333 net422 VGND VGND VPWR VPWR _09382_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16346_ _08356_ _08358_ _08435_ VGND VGND VPWR VPWR _08436_ sky130_fd_sc_hd__a21oi_2
X_19134_ net424 _11096_ _11102_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__a21o_1
X_13558_ _05685_ _05691_ _05681_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19065_ _10992_ VGND VGND VPWR VPWR _11037_ sky130_fd_sc_hd__inv_2
X_16277_ _08366_ _08367_ VGND VGND VPWR VPWR _08368_ sky130_fd_sc_hd__xnor2_1
X_13489_ _05477_ _05480_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18016_ _09990_ _10000_ VGND VGND VPWR VPWR _10001_ sky130_fd_sc_hd__xnor2_2
X_15228_ net522 _07244_ _07325_ _07326_ _07324_ VGND VGND VPWR VPWR _07327_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15159_ net517 net485 _07256_ _07257_ VGND VGND VPWR VPWR _07258_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout108 top0.cordic0.vec\[1\]\[12\] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_4
X_19967_ _11410_ _11511_ _11833_ _11835_ _11827_ VGND VGND VPWR VPWR _11836_ sky130_fd_sc_hd__a311o_2
Xfanout119 net120 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_4
X_18918_ _10813_ _10814_ _10809_ VGND VGND VPWR VPWR _10893_ sky130_fd_sc_hd__o21a_1
X_19898_ net228 _11764_ VGND VGND VPWR VPWR _11772_ sky130_fd_sc_hd__nand2_1
X_18849_ _10824_ VGND VGND VPWR VPWR _10825_ sky130_fd_sc_hd__inv_2
XFILLER_0_179_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21860_ _01408_ _01409_ _01419_ _01420_ _01421_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20811_ _11608_ net254 _12559_ _12659_ VGND VGND VPWR VPWR _12660_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_78_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21791_ _01352_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23530_ top0.a_in_matmul\[5\] top0.matmul0.a\[5\] _02926_ VGND VGND VPWR VPWR _02931_
+ sky130_fd_sc_hd__mux2_1
X_20742_ net295 _12553_ _11437_ VGND VGND VPWR VPWR _12591_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23461_ top0.cordic0.sin\[0\] top0.matmul0.sin\[0\] _05461_ VGND VGND VPWR VPWR _02895_
+ sky130_fd_sc_hd__mux2_1
X_20673_ _11689_ _12499_ _12490_ VGND VGND VPWR VPWR _12522_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_190_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25200_ _03343_ _03936_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22412_ _01966_ _01969_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26180_ _05316_ top0.cordic0.slte0.opB\[11\] _12003_ VGND VGND VPWR VPWR _05317_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23392_ _01213_ _02831_ _02832_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25131_ _04477_ _04478_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22343_ _01643_ net91 _01845_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__o21ai_1
X_25062_ _04252_ _03305_ _03829_ _04258_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__and4_2
XFILLER_0_131_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22274_ net143 net126 _01113_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__or3b_1
X_24013_ _03248_ _03323_ _03365_ _03368_ _03370_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__a311o_2
Xhold140 top0.c_out_calc\[10\] VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__dlygate4sd3_1
X_21225_ _12622_ _13068_ _12627_ VGND VGND VPWR VPWR _13069_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold151 top0.svm0.tC\[13\] VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 top0.matmul0.matmul_stage_inst.b\[0\] VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 top0.pid_q.prev_error\[13\] VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 top0.pid_d.prev_error\[5\] VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 top0.periodTop\[12\] VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__dlygate4sd3_1
X_21156_ net223 net219 VGND VGND VPWR VPWR _13001_ sky130_fd_sc_hd__nand2_2
Xfanout620 net629 VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__clkbuf_2
Xfanout631 net635 VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__clkbuf_4
Xfanout642 net645 VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__clkbuf_4
X_20107_ top0.cordic0.slte0.opA\[13\] _11957_ _11960_ VGND VGND VPWR VPWR _11965_
+ sky130_fd_sc_hd__o21ba_1
Xfanout653 net654 VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__buf_2
X_21087_ _12899_ _12932_ VGND VGND VPWR VPWR _12933_ sky130_fd_sc_hd__xnor2_2
X_25964_ top0.pid_q.out\[1\] _12032_ _05014_ spi0.data_packed\[49\] VGND VGND VPWR
+ VPWR _05173_ sky130_fd_sc_hd__a22o_1
Xfanout664 net666 VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__buf_4
Xfanout675 net687 VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__clkbuf_4
Xfanout686 net687 VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__clkbuf_4
X_24915_ _04206_ _04208_ _04265_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__o21a_1
X_20038_ _11612_ _11518_ VGND VGND VPWR VPWR _11902_ sky130_fd_sc_hd__nand2_1
Xfanout697 net700 VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_198_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25895_ top0.matmul0.alpha_pass\[10\] net429 _05110_ _05111_ VGND VGND VPWR VPWR
+ _05112_ sky130_fd_sc_hd__o31a_1
X_24846_ _04094_ _04196_ _04197_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_73_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24777_ _03830_ _04129_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__nor2_1
X_21989_ _01312_ _01550_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__or2b_1
XFILLER_0_200_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14530_ _06736_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__inv_2
X_26516_ clknet_leaf_66_clk_sys _00139_ net659 VGND VGND VPWR VPWR top0.pid_q.out\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_23728_ _03053_ _03083_ _03084_ _03085_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__o22a_2
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14461_ _06596_ _06664_ _06594_ VGND VGND VPWR VPWR _06669_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26447_ clknet_leaf_59_clk_sys _00088_ net644 VGND VGND VPWR VPWR top0.kiq\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23659_ _03015_ _03016_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__nor2_4
XFILLER_0_126_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16200_ net500 _08169_ _08291_ VGND VGND VPWR VPWR _08292_ sky130_fd_sc_hd__o21ai_1
X_13412_ _05624_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17180_ net543 _05441_ _09134_ VGND VGND VPWR VPWR _09191_ sky130_fd_sc_hd__and3_1
X_14392_ _06598_ _06600_ VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__xnor2_1
X_26378_ clknet_leaf_40_clk_sys _00019_ net682 VGND VGND VPWR VPWR top0.svm0.tC\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16131_ _08219_ _08223_ VGND VGND VPWR VPWR _08224_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25329_ _04621_ _04622_ _04620_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__o21ba_1
X_13343_ _05553_ _05555_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16062_ _08153_ _08155_ VGND VGND VPWR VPWR _08156_ sky130_fd_sc_hd__xnor2_1
X_13274_ net38 _05484_ _05486_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__and3_1
X_15013_ spi0.data_packed\[12\] top0.periodTop\[12\] _07125_ VGND VGND VPWR VPWR _07132_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19821_ _11676_ _11677_ _11692_ VGND VGND VPWR VPWR _11700_ sky130_fd_sc_hd__or3_1
XFILLER_0_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19752_ net120 net116 net103 net98 net200 net187 VGND VGND VPWR VPWR _11635_ sky130_fd_sc_hd__mux4_1
X_16964_ _09019_ _09020_ VGND VGND VPWR VPWR _09021_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_16_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18703_ top0.pid_d.out\[9\] _10680_ _07141_ VGND VGND VPWR VPWR _10681_ sky130_fd_sc_hd__mux2_1
X_15915_ _08001_ _08009_ VGND VGND VPWR VPWR _08010_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19683_ net291 _11435_ _11568_ VGND VGND VPWR VPWR _11570_ sky130_fd_sc_hd__and3_1
X_16895_ net473 _08890_ _08956_ _08930_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__o211a_1
XFILLER_0_194_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18634_ _09706_ net377 VGND VGND VPWR VPWR _10612_ sky130_fd_sc_hd__nor2_1
X_15846_ _07938_ _07941_ VGND VGND VPWR VPWR _07942_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_189_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_201_Right_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18565_ net331 net368 VGND VGND VPWR VPWR _10544_ sky130_fd_sc_hd__nand2_1
X_15777_ net506 net483 VGND VGND VPWR VPWR _07874_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17516_ net395 _09496_ _09497_ _09495_ _09502_ VGND VGND VPWR VPWR _09503_ sky130_fd_sc_hd__o221a_2
X_14728_ _06892_ _06887_ VGND VGND VPWR VPWR _06931_ sky130_fd_sc_hd__and2b_1
XFILLER_0_185_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18496_ _10472_ _10475_ VGND VGND VPWR VPWR _10476_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14659_ _06861_ _06862_ VGND VGND VPWR VPWR _06863_ sky130_fd_sc_hd__nand2_2
X_17447_ _09431_ _09432_ _09433_ VGND VGND VPWR VPWR _09434_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_200_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_25_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17378_ net410 net405 VGND VGND VPWR VPWR _09365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19117_ net435 _11029_ _11077_ _11088_ VGND VGND VPWR VPWR _11089_ sky130_fd_sc_hd__a31o_1
X_16329_ _08417_ _08418_ VGND VGND VPWR VPWR _08419_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19048_ net374 _11019_ _11020_ VGND VGND VPWR VPWR _11021_ sky130_fd_sc_hd__o21ai_2
Xclkbuf_leaf_89_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_89_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21010_ _12851_ _12856_ VGND VGND VPWR VPWR _12857_ sky130_fd_sc_hd__xor2_2
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_34_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22961_ _02472_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24700_ _03944_ _03939_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__or2b_1
X_21912_ _01462_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__inv_2
X_25680_ top0.matmul0.sin\[11\] _04949_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__xor2_1
X_22892_ _02352_ top0.svm0.tC\[1\] top0.svm0.tC\[0\] _02298_ VGND VGND VPWR VPWR _02410_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24631_ _02994_ _02996_ _03029_ _03030_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__o22a_1
X_21843_ _01397_ _01403_ _01389_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24562_ _03767_ _03772_ _03763_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__a21o_1
X_21774_ net152 _01325_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_43_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26301_ _05382_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__clkbuf_1
X_23513_ top0.cordic0.cos\[11\] top0.matmul0.cos\[11\] _02915_ VGND VGND VPWR VPWR
+ _02922_ sky130_fd_sc_hd__mux2_1
X_20725_ net306 _12571_ VGND VGND VPWR VPWR _12574_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27281_ clknet_3_0__leaf_clk_mosi _00895_ VGND VGND VPWR VPWR spi0.data_packed\[67\]
+ sky130_fd_sc_hd__dfxtp_1
X_24493_ _03752_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26232_ net19 spi0.data_packed\[15\] net695 VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__mux2_1
X_23444_ _11519_ _02879_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__or2_1
X_20656_ net298 _12504_ VGND VGND VPWR VPWR _12505_ sky130_fd_sc_hd__or2_1
XFILLER_0_191_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26163_ spi0.data_packed\[5\] _05299_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23375_ net120 _02799_ _02816_ _02785_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_162_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20587_ net270 net258 net245 VGND VGND VPWR VPWR _12436_ sky130_fd_sc_hd__and3_1
X_25114_ _04387_ _04389_ _04462_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__o21a_1
X_22326_ _01873_ _01883_ _01884_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__a21boi_4
X_26094_ top0.a_in_matmul\[15\] _05272_ _05164_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25045_ _04382_ _04303_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22257_ _01755_ _01815_ _01816_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_52_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21208_ _13049_ _13051_ VGND VGND VPWR VPWR _13052_ sky130_fd_sc_hd__nand2_1
X_22188_ net131 _01144_ _01708_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21139_ _12134_ _12983_ net267 VGND VGND VPWR VPWR _12984_ sky130_fd_sc_hd__mux2_1
X_26996_ clknet_leaf_24_clk_sys _00613_ net625 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[12\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout450 net451 VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkbuf_2
Xfanout461 net463 VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__buf_4
Xfanout472 top0.pid_q.mult0.b\[5\] VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__buf_2
X_13961_ _05786_ _05787_ _06173_ _06171_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__o211a_1
X_25947_ net428 _05158_ _05159_ top0.matmul0.alpha_pass\[14\] VGND VGND VPWR VPWR
+ _05160_ sky130_fd_sc_hd__a22oi_1
Xfanout483 top0.pid_q.mult0.b\[3\] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__buf_4
Xfanout494 net496 VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__dlymetal6s2s_1
X_15700_ _07796_ _07797_ VGND VGND VPWR VPWR _07798_ sky130_fd_sc_hd__xnor2_1
X_16680_ net449 _08696_ VGND VGND VPWR VPWR _08765_ sky130_fd_sc_hd__nor2_1
X_13892_ net1030 _05893_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__nand2_1
X_25878_ top0.matmul0.beta_pass\[8\] _05095_ _05096_ net1024 VGND VGND VPWR VPWR _05097_
+ sky130_fd_sc_hd__a22o_1
Xmax_cap8 _03432_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_159_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24829_ _03313_ _03720_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__nand2_2
XFILLER_0_159_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15631_ _07727_ _07728_ VGND VGND VPWR VPWR _07729_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_61_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18350_ _10330_ _10331_ VGND VGND VPWR VPWR _10332_ sky130_fd_sc_hd__or2_1
X_15562_ _07288_ _07286_ VGND VGND VPWR VPWR _07661_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14513_ _05586_ _06640_ net23 VGND VGND VPWR VPWR _06720_ sky130_fd_sc_hd__o21a_1
X_17301_ _09294_ _09295_ VGND VGND VPWR VPWR _09296_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18281_ _10261_ _10262_ VGND VGND VPWR VPWR _10263_ sky130_fd_sc_hd__xor2_2
X_15493_ _07590_ _07591_ _07281_ VGND VGND VPWR VPWR _07592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14444_ _06636_ _06651_ VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__xnor2_4
X_17232_ top0.pid_q.curr_int\[14\] _09236_ VGND VGND VPWR VPWR _09237_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout90 net93 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_4
X_17163_ _00007_ _09134_ VGND VGND VPWR VPWR _09176_ sky130_fd_sc_hd__nand2_1
X_14375_ net33 _05551_ VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16114_ _08100_ _08102_ _08206_ VGND VGND VPWR VPWR _08207_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13326_ net1024 _05466_ _05467_ _05464_ top0.c_out_calc\[8\] VGND VGND VPWR VPWR
+ _05539_ sky130_fd_sc_hd__a32o_2
XFILLER_0_161_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17094_ net849 _09115_ _09123_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_90_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_90_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_70_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16045_ _08039_ _08059_ VGND VGND VPWR VPWR _08139_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13257_ _05469_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__buf_6
XFILLER_0_150_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19804_ _11680_ _11683_ VGND VGND VPWR VPWR _11685_ sky130_fd_sc_hd__and2_1
XFILLER_0_202_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17996_ top0.pid_d.out\[0\] top0.pid_d.curr_int\[0\] top0.pid_d.curr_int\[1\] top0.pid_d.out\[1\]
+ VGND VGND VPWR VPWR _09981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19735_ _11616_ _11618_ VGND VGND VPWR VPWR _11619_ sky130_fd_sc_hd__xor2_4
X_16947_ _09003_ _08990_ _09004_ VGND VGND VPWR VPWR _09005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19666_ net94 net88 net200 VGND VGND VPWR VPWR _11553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16878_ _08939_ _08940_ VGND VGND VPWR VPWR _08941_ sky130_fd_sc_hd__xnor2_1
X_18617_ _10594_ _10514_ top0.pid_d.out\[8\] VGND VGND VPWR VPWR _10595_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_56_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15829_ _07921_ _07923_ VGND VGND VPWR VPWR _07925_ sky130_fd_sc_hd__nor2_1
X_19597_ _11485_ top0.cordic0.slte0.opA\[8\] VGND VGND VPWR VPWR _11486_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18548_ net396 net309 VGND VGND VPWR VPWR _10527_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18479_ _10383_ _10387_ _10457_ _10458_ net341 VGND VGND VPWR VPWR _10459_ sky130_fd_sc_hd__a32o_1
XFILLER_0_173_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20510_ _12325_ _12357_ _12358_ VGND VGND VPWR VPWR _12359_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21490_ _01024_ _01049_ _01022_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__or3b_1
XFILLER_0_15_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20441_ net275 _12284_ _12289_ VGND VGND VPWR VPWR _12290_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_43_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23160_ _02643_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__buf_6
XFILLER_0_166_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20372_ _11437_ _12131_ VGND VGND VPWR VPWR _12221_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22111_ _01640_ _01660_ _01653_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__and3b_1
XFILLER_0_101_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23091_ _02573_ _02587_ _02589_ _02591_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22042_ _01213_ _01286_ _01287_ _01600_ _01603_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__a221oi_2
X_26850_ clknet_leaf_46_clk_sys _00467_ net681 VGND VGND VPWR VPWR top0.svm0.delta\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_103_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25801_ _05028_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__buf_2
X_26781_ clknet_leaf_109_clk_sys _00398_ net579 VGND VGND VPWR VPWR top0.cordic0.sin\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_23993_ _03337_ _03338_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__nand2_1
X_25732_ top0.matmul0.sin\[11\] _04985_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__xnor2_1
X_22944_ _02457_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25663_ _04884_ _04931_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__and2_1
X_22875_ _02367_ top0.svm0.tB\[8\] _02393_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24614_ _03907_ _03913_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__or2_1
X_21826_ _01379_ _01383_ _01387_ _01385_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__a31o_1
XFILLER_0_167_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25594_ net759 _00000_ _04882_ _04887_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__o22a_1
XFILLER_0_183_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24545_ _03152_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__buf_4
X_21757_ net163 VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20708_ net285 _12552_ _12555_ _12278_ _12556_ VGND VGND VPWR VPWR _12557_ sky130_fd_sc_hd__a311o_1
X_27264_ clknet_3_6__leaf_clk_mosi _00878_ VGND VGND VPWR VPWR spi0.data_packed\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_24476_ _03824_ _03831_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_164_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21688_ _01130_ _01162_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__and2_1
XFILLER_0_191_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26215_ _05339_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23427_ net98 _02863_ _02864_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__a21bo_1
X_27195_ clknet_leaf_56_clk_sys _00809_ net666 VGND VGND VPWR VPWR top0.currT_r\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_20639_ _12463_ _12475_ VGND VGND VPWR VPWR _12488_ sky130_fd_sc_hd__nor2_1
XFILLER_0_190_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14160_ _06256_ _06266_ _06371_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26146_ spi0.data_packed\[2\] _05289_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__xor2_1
X_23358_ _02800_ _02791_ _01408_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__o21a_1
X_22309_ _01796_ _01801_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__nand2_1
X_14091_ _06295_ _06302_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__xnor2_4
X_26077_ top0.matmul0.alpha_pass\[11\] _05237_ _05259_ VGND VGND VPWR VPWR _05260_
+ sky130_fd_sc_hd__a21o_1
X_23289_ _11784_ _02735_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__nor2_1
X_25028_ _04287_ _04299_ _04285_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__a21bo_1
X_17850_ _09835_ _09836_ VGND VGND VPWR VPWR _09837_ sky130_fd_sc_hd__xnor2_1
X_16801_ top0.kiq\[10\] _08863_ _08866_ VGND VGND VPWR VPWR _08874_ sky130_fd_sc_hd__and3_1
X_17781_ _09677_ _09680_ VGND VGND VPWR VPWR _09768_ sky130_fd_sc_hd__nor2_1
X_26979_ clknet_leaf_29_clk_sys _00596_ net624 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_14993_ _07121_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__clkbuf_1
Xfanout280 net284 VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkbuf_4
Xfanout291 net292 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__buf_4
X_19520_ net201 VGND VGND VPWR VPWR _11410_ sky130_fd_sc_hd__inv_2
X_16732_ _08812_ _08815_ VGND VGND VPWR VPWR _08816_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13944_ _05779_ _05781_ _06156_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_37_clk_sys clknet_3_7__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_37_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_163_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19451_ net441 _11347_ _11348_ _11200_ VGND VGND VPWR VPWR _11349_ sky130_fd_sc_hd__a31o_1
XFILLER_0_186_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13875_ _05765_ _05766_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__and2_1
X_16663_ _08717_ _08722_ _08716_ VGND VGND VPWR VPWR _08748_ sky130_fd_sc_hd__o21a_1
XFILLER_0_201_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18402_ _10271_ _10273_ _10382_ VGND VGND VPWR VPWR _10383_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_57_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15614_ _07616_ _07711_ _07695_ VGND VGND VPWR VPWR _07712_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19382_ top0.pid_d.prev_error\[15\] _11284_ _11287_ net722 VGND VGND VPWR VPWR _00325_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16594_ top0.pid_q.out\[12\] _07705_ _08627_ net544 _08680_ VGND VGND VPWR VPWR _08681_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18333_ _10229_ _10314_ VGND VGND VPWR VPWR _10315_ sky130_fd_sc_hd__xnor2_1
X_15545_ _07576_ _07577_ _07643_ VGND VGND VPWR VPWR _07644_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18264_ top0.pid_d.curr_int\[4\] _10159_ _10245_ VGND VGND VPWR VPWR _10246_ sky130_fd_sc_hd__o21ai_2
X_15476_ _07569_ _07574_ VGND VGND VPWR VPWR _07575_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14427_ _06632_ _06634_ VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__xor2_2
XFILLER_0_182_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17215_ _08685_ VGND VGND VPWR VPWR _09222_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18195_ _10176_ _10177_ VGND VGND VPWR VPWR _10178_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14358_ _06495_ _06497_ _06566_ VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__o21a_1
X_17146_ net543 _07991_ _09161_ VGND VGND VPWR VPWR _09162_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13309_ net47 _05520_ _05521_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__and3_1
X_17077_ net885 _09100_ _09102_ _09090_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__a22o_1
X_14289_ _06495_ _06498_ VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__xor2_4
XFILLER_0_150_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16028_ _08042_ _08043_ _08041_ VGND VGND VPWR VPWR _08122_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_108_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17979_ net314 VGND VGND VPWR VPWR _09965_ sky130_fd_sc_hd__inv_2
X_19718_ _11585_ _11586_ _11587_ _11571_ VGND VGND VPWR VPWR _11603_ sky130_fd_sc_hd__o31a_1
X_20990_ net267 _12135_ VGND VGND VPWR VPWR _12837_ sky130_fd_sc_hd__or2_1
XFILLER_0_196_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19649_ net133 net128 net123 net121 net199 net193 VGND VGND VPWR VPWR _11537_ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22660_ net720 _12813_ _02212_ _12742_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21611_ _01073_ _01077_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22591_ net79 _02144_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24330_ _03162_ _03163_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__or2_2
XFILLER_0_47_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21542_ _01078_ _01103_ net158 VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_117_Left_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24261_ _03439_ _03440_ _03438_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21473_ _01033_ _01036_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26000_ top0.matmul0.beta_pass\[9\] _05169_ _05200_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__a21o_1
X_23212_ net237 net233 net228 net223 net204 net196 VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__mux4_2
X_20424_ net275 net289 VGND VGND VPWR VPWR _12273_ sky130_fd_sc_hd__or2b_1
X_24192_ _03542_ _03543_ VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23143_ _02631_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__clkbuf_1
X_20355_ _12198_ _12200_ _12203_ VGND VGND VPWR VPWR _12204_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23074_ net63 top0.svm0.counter\[1\] VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__xor2_1
XFILLER_0_144_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20286_ net238 _12134_ VGND VGND VPWR VPWR _12135_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_105_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22025_ net153 _01299_ _01578_ _01581_ _01586_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__o311a_1
X_26902_ clknet_leaf_4_clk_sys _00519_ net585 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold11 top0.matmul0.matmul_stage_inst.b\[15\] VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold22 top0.pid_d.curr_error\[15\] VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__dlygate4sd3_1
X_26833_ clknet_leaf_42_clk_sys _00450_ net684 VGND VGND VPWR VPWR top0.svm0.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold33 top0.cordic0.sin\[11\] VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 state\[1\] VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 top0.matmul0.matmul_stage_inst.d\[6\] VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 _00324_ VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 top0.svm0.tA\[13\] VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 top0.svm0.tA\[7\] VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__dlygate4sd3_1
X_23976_ _03332_ _03333_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__xor2_1
X_26764_ clknet_leaf_87_clk_sys _00381_ net642 VGND VGND VPWR VPWR top0.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold99 top0.matmul0.matmul_stage_inst.c\[5\] VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22927_ _02442_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__clkbuf_1
X_25715_ net866 _04964_ _04936_ _04974_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26695_ clknet_leaf_71_clk_sys net893 net657 VGND VGND VPWR VPWR top0.pid_d.prev_error\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13660_ _05865_ _05868_ _05872_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__o21a_1
X_22858_ net168 _02376_ _02377_ _02314_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__a211o_1
XFILLER_0_168_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25646_ net69 top0.matmul0.sin\[4\] VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21809_ _01331_ _01332_ _01301_ net162 _01370_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__o221ai_1
X_13591_ _05626_ _05639_ _05622_ net66 VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__o22a_1
X_25577_ top0.matmul0.a\[11\] top0.matmul0.matmul_stage_inst.e\[11\] _04867_ VGND
+ VGND VPWR VPWR _04876_ sky130_fd_sc_hd__mux2_1
X_22789_ _02310_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15330_ _07390_ _07428_ VGND VGND VPWR VPWR _07429_ sky130_fd_sc_hd__xnor2_1
X_24528_ _03024_ _03025_ _03054_ _03055_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__o22a_2
XFILLER_0_54_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15261_ _07358_ _07359_ VGND VGND VPWR VPWR _07360_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_151_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24459_ _03783_ _03814_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__xor2_1
X_27247_ clknet_3_2__leaf_clk_mosi _00861_ VGND VGND VPWR VPWR spi0.data_packed\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_14212_ _05688_ _05543_ _05545_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__or3_2
X_17000_ top0.pid_q.prev_error\[13\] top0.pid_q.curr_error\[13\] VGND VGND VPWR VPWR
+ _09054_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15192_ _07289_ _07290_ VGND VGND VPWR VPWR _07291_ sky130_fd_sc_hd__xor2_4
X_27178_ clknet_leaf_88_clk_sys _00792_ net642 VGND VGND VPWR VPWR top0.periodTop_r\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_8 _09593_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14143_ _06191_ _06193_ _06349_ _06354_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__a31o_1
X_26129_ spi0.data_packed\[24\] _05281_ _05282_ net948 VGND VGND VPWR VPWR _00805_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14074_ net48 _05604_ _06184_ _05624_ net51 VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__a32o_1
X_18951_ _10828_ _10924_ VGND VGND VPWR VPWR _10925_ sky130_fd_sc_hd__or2_1
X_17902_ _09885_ _09888_ VGND VGND VPWR VPWR _09889_ sky130_fd_sc_hd__xor2_1
X_18882_ _10850_ _10856_ VGND VGND VPWR VPWR _10857_ sky130_fd_sc_hd__xnor2_1
X_17833_ _09817_ _09819_ _09718_ _09740_ VGND VGND VPWR VPWR _09820_ sky130_fd_sc_hd__o22a_1
XFILLER_0_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17764_ _09743_ VGND VGND VPWR VPWR _09751_ sky130_fd_sc_hd__inv_2
X_14976_ _07110_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19503_ net441 _11394_ VGND VGND VPWR VPWR _11395_ sky130_fd_sc_hd__nand2_1
X_16715_ _08747_ _08782_ _08798_ VGND VGND VPWR VPWR _08799_ sky130_fd_sc_hd__a21oi_1
X_13927_ net1025 _05624_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_199_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17695_ _09674_ _09681_ VGND VGND VPWR VPWR _09682_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19434_ top0.pid_d.curr_int\[6\] _11290_ _11293_ _11333_ VGND VGND VPWR VPWR _00332_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_179_Right_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16646_ _08728_ _08731_ VGND VGND VPWR VPWR _08732_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13858_ _05992_ _05993_ _06022_ _06070_ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_187_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19365_ _11286_ VGND VGND VPWR VPWR _11287_ sky130_fd_sc_hd__buf_2
XFILLER_0_186_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16577_ _08312_ _08663_ VGND VGND VPWR VPWR _08664_ sky130_fd_sc_hd__nand2_1
X_13789_ _06000_ _06001_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18316_ _10287_ _10297_ VGND VGND VPWR VPWR _10298_ sky130_fd_sc_hd__xor2_1
XFILLER_0_139_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15528_ _07625_ _07626_ VGND VGND VPWR VPWR _07627_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19296_ top0.pid_d.prev_error\[11\] top0.pid_d.curr_error\[11\] VGND VGND VPWR VPWR
+ _11238_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18247_ _10227_ _10229_ VGND VGND VPWR VPWR _10230_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15459_ net489 net508 VGND VGND VPWR VPWR _07558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18178_ _10159_ _10160_ VGND VGND VPWR VPWR _10161_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17129_ top0.pid_q.curr_int\[1\] _09141_ _09146_ _09136_ VGND VGND VPWR VPWR _00214_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20140_ _11994_ _11995_ net212 _11519_ VGND VGND VPWR VPWR _11996_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_111_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20071_ _11931_ _11932_ VGND VGND VPWR VPWR _11933_ sky130_fd_sc_hd__and2b_1
XFILLER_0_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23830_ _03045_ _03046_ _03018_ _03019_ VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__o22a_1
XFILLER_0_174_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23761_ _03115_ _03118_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_196_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20973_ net236 _11739_ VGND VGND VPWR VPWR _12820_ sky130_fd_sc_hd__nor2_2
XFILLER_0_135_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25500_ top0.matmul0.matmul_stage_inst.mult1\[6\] _04243_ _04829_ VGND VGND VPWR
+ VPWR _04836_ sky130_fd_sc_hd__mux2_1
X_22712_ _02125_ _02171_ _02173_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__o21a_1
XFILLER_0_178_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26480_ clknet_leaf_11_clk_sys _00111_ net601 VGND VGND VPWR VPWR top0.periodTop\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23692_ _03018_ _03019_ _03027_ _03028_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__o22a_2
XFILLER_0_178_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25431_ _04646_ _04773_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__nand2_1
X_22643_ _02194_ _02195_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25362_ _04664_ _04703_ _04705_ _04706_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22574_ _02007_ _02084_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24313_ _03225_ _03226_ _03669_ _03110_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__a31o_1
X_27101_ clknet_leaf_20_clk_sys _00718_ net609 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.a\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_21525_ _01063_ _01064_ _01068_ _01085_ _01086_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__a221oi_4
X_25293_ _04553_ _04566_ _04565_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27032_ clknet_leaf_15_clk_sys _00649_ net613 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_24244_ _03513_ _03515_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__xor2_1
XFILLER_0_161_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21456_ _00996_ _01012_ _01011_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20407_ _12253_ _12255_ VGND VGND VPWR VPWR _12256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24175_ _03528_ _03530_ _03531_ _03532_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__o22a_2
XFILLER_0_181_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21387_ _13159_ _13184_ _13185_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__o21ba_1
X_23126_ _07117_ _02618_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__nor2_1
X_20338_ _12182_ _12183_ VGND VGND VPWR VPWR _12187_ sky130_fd_sc_hd__nand2_2
X_23057_ top0.svm0.counter\[5\] _02557_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__xnor2_1
X_20269_ net289 _11571_ VGND VGND VPWR VPWR _12118_ sky130_fd_sc_hd__nand2_1
X_22008_ _01319_ net158 _01310_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__or3_1
X_14830_ _06867_ _05726_ _05727_ VGND VGND VPWR VPWR _07029_ sky130_fd_sc_hd__and3b_1
X_26816_ clknet_leaf_60_clk_sys _00433_ net652 VGND VGND VPWR VPWR top0.pid_q.prev_int\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14761_ net33 _06824_ _06961_ _06962_ VGND VGND VPWR VPWR _06963_ sky130_fd_sc_hd__a31o_1
X_26747_ clknet_leaf_92_clk_sys _00364_ net599 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_23959_ _03015_ _03016_ _02989_ _02991_ VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__o22a_2
X_16500_ _08521_ _08530_ _08529_ VGND VGND VPWR VPWR _08588_ sky130_fd_sc_hd__a21o_1
X_13712_ _05901_ _05899_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__xnor2_1
X_14692_ _06893_ _06895_ VGND VGND VPWR VPWR _06896_ sky130_fd_sc_hd__nor2_1
X_17480_ _09458_ _09461_ _09465_ _09466_ VGND VGND VPWR VPWR _09467_ sky130_fd_sc_hd__a22o_1
X_26678_ clknet_leaf_64_clk_sys _00295_ net656 VGND VGND VPWR VPWR top0.pid_d.curr_error\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16431_ _08509_ _08519_ VGND VGND VPWR VPWR _08520_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13643_ _05801_ _05855_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__nand2_1
X_25629_ net72 _04908_ _04890_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19150_ net389 _11096_ _11110_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__a21o_1
X_13574_ _05785_ _05754_ _05755_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__and3_1
X_16362_ net468 net473 net476 _08286_ VGND VGND VPWR VPWR _08452_ sky130_fd_sc_hd__and4_1
XFILLER_0_13_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18101_ _10079_ _10084_ VGND VGND VPWR VPWR _10085_ sky130_fd_sc_hd__nor2_1
X_15313_ net533 net487 VGND VGND VPWR VPWR _07412_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16293_ _08142_ _08383_ VGND VGND VPWR VPWR _08384_ sky130_fd_sc_hd__xnor2_1
X_19081_ net370 net308 VGND VGND VPWR VPWR _11053_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18032_ net1022 net398 VGND VGND VPWR VPWR _10017_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15244_ _07328_ _07334_ _07337_ _07342_ VGND VGND VPWR VPWR _07343_ sky130_fd_sc_hd__or4b_1
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15175_ net489 net511 VGND VGND VPWR VPWR _07274_ sky130_fd_sc_hd__and2_2
XFILLER_0_23_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14126_ _06331_ _06337_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__xor2_2
XFILLER_0_162_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19983_ top0.cordic0.slte0.opA\[3\] VGND VGND VPWR VPWR _11851_ sky130_fd_sc_hd__inv_2
XFILLER_0_197_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14057_ _06133_ _06269_ _06258_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__and3b_1
XFILLER_0_120_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18934_ _10841_ _10905_ _10906_ _10908_ VGND VGND VPWR VPWR _10909_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18865_ _10606_ _10683_ _10677_ VGND VGND VPWR VPWR _10840_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17816_ _09795_ _09802_ VGND VGND VPWR VPWR _09803_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18796_ _10770_ _10771_ net362 VGND VGND VPWR VPWR _10772_ sky130_fd_sc_hd__o21ai_4
X_17747_ _09506_ _09728_ _09730_ _09510_ VGND VGND VPWR VPWR _09734_ sky130_fd_sc_hd__a2bb2o_1
X_14959_ _07101_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__clkbuf_1
X_17678_ net322 net420 VGND VGND VPWR VPWR _09665_ sky130_fd_sc_hd__nor2_1
X_19417_ top0.pid_d.curr_int\[4\] top0.pid_d.prev_int\[4\] VGND VGND VPWR VPWR _11319_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_187_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16629_ _08713_ _08714_ VGND VGND VPWR VPWR _08715_ sky130_fd_sc_hd__or2b_1
XFILLER_0_159_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19348_ _11180_ _11181_ _11279_ _11273_ top0.pid_d.curr_error\[6\] VGND VGND VPWR
+ VPWR _00300_ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19279_ _11221_ _11222_ VGND VGND VPWR VPWR _11223_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21310_ _13104_ _13105_ _13145_ VGND VGND VPWR VPWR _13152_ sky130_fd_sc_hd__mux2_1
X_22290_ net78 net99 VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21241_ _12609_ _13080_ _13081_ _13083_ _13084_ VGND VGND VPWR VPWR _13085_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold300 top0.cordic0.sin\[7\] VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 spi0.data_packed\[43\] VGND VGND VPWR VPWR net1011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21172_ _12998_ _13005_ _13004_ VGND VGND VPWR VPWR _13016_ sky130_fd_sc_hd__a21oi_2
X_20123_ _11428_ _11947_ _11978_ _11976_ VGND VGND VPWR VPWR _11980_ sky130_fd_sc_hd__a211o_1
XFILLER_0_111_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25980_ top0.pid_q.out\[5\] _12032_ _05014_ spi0.data_packed\[53\] VGND VGND VPWR
+ VPWR _05185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24931_ _04280_ _04281_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__xnor2_1
X_20054_ _11410_ _11916_ VGND VGND VPWR VPWR _11917_ sky130_fd_sc_hd__nor2_1
X_24862_ _04104_ _04120_ _04213_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__a21oi_1
X_26601_ clknet_leaf_68_clk_sys _00224_ net659 VGND VGND VPWR VPWR top0.pid_q.curr_int\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_139_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23813_ _03014_ _03033_ _03003_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__a21o_1
XFILLER_0_169_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24793_ _04035_ _04142_ _04144_ _04032_ _04145_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__o221ai_2
X_23744_ _03063_ _03064_ _03090_ _03091_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__o22a_2
XFILLER_0_75_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26532_ clknet_leaf_61_clk_sys _00155_ net651 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_20956_ _12746_ _12803_ VGND VGND VPWR VPWR _12804_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23675_ _03021_ _03032_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__xnor2_2
X_26463_ clknet_leaf_16_clk_sys net560 net611 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20887_ _12730_ _12735_ VGND VGND VPWR VPWR _12736_ sky130_fd_sc_hd__nor2_2
XFILLER_0_95_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25414_ _04664_ _04755_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22626_ net724 _12004_ _12740_ _02179_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__a31o_1
X_26394_ clknet_leaf_86_clk_sys _00035_ net640 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfstp_2
XFILLER_0_64_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25345_ _04683_ _04689_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22557_ net107 net101 VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21508_ net124 net118 _01069_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__a21o_1
X_25276_ _03280_ _04182_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__nor2_1
X_13290_ net38 _05489_ _05491_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__and3_1
X_22488_ _02009_ _02044_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__xnor2_1
X_27015_ clknet_leaf_24_clk_sys _00632_ net626 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_24227_ _03464_ _03545_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__xor2_2
XFILLER_0_146_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21439_ _12180_ _12238_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24158_ _03513_ _03515_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__or2_2
X_23109_ _02458_ _02598_ _02604_ _02606_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24089_ _03436_ _03446_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__xnor2_4
X_16980_ _09033_ _09035_ VGND VGND VPWR VPWR _09036_ sky130_fd_sc_hd__xnor2_2
X_15931_ _08017_ _08025_ VGND VGND VPWR VPWR _08026_ sky130_fd_sc_hd__xnor2_1
X_18650_ _10626_ _10627_ VGND VGND VPWR VPWR _10628_ sky130_fd_sc_hd__nor2_1
X_15862_ _07952_ _07957_ VGND VGND VPWR VPWR _07958_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17601_ net425 _09582_ _09584_ _09586_ _09587_ VGND VGND VPWR VPWR _09588_ sky130_fd_sc_hd__a311o_1
X_14813_ _07009_ _07010_ _07012_ VGND VGND VPWR VPWR _07013_ sky130_fd_sc_hd__o21a_1
XFILLER_0_153_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18581_ _10464_ _10488_ _10487_ VGND VGND VPWR VPWR _10560_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_118_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15793_ _07888_ _07889_ VGND VGND VPWR VPWR _07890_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17532_ net415 net412 _09354_ VGND VGND VPWR VPWR _09519_ sky130_fd_sc_hd__and3_1
X_14744_ _06910_ _06943_ VGND VGND VPWR VPWR _06946_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17463_ _09376_ _09379_ _09384_ VGND VGND VPWR VPWR _09450_ sky130_fd_sc_hd__o21ai_1
X_14675_ _06873_ _06878_ VGND VGND VPWR VPWR _06879_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19202_ net346 _11094_ VGND VGND VPWR VPWR _11153_ sky130_fd_sc_hd__or2_1
X_16414_ net516 net445 VGND VGND VPWR VPWR _08503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13626_ net47 _05489_ _05491_ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__and3_1
X_17394_ net330 net427 VGND VGND VPWR VPWR _09381_ sky130_fd_sc_hd__nand2_1
X_19133_ top0.kid\[1\] _11098_ _11100_ top0.kpd\[1\] VGND VGND VPWR VPWR _11102_ sky130_fd_sc_hd__a22o_1
X_16345_ _08356_ _08358_ _08357_ VGND VGND VPWR VPWR _08435_ sky130_fd_sc_hd__o21a_1
X_13557_ _05760_ _05769_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_183_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19064_ top0.pid_d.out\[14\] _09339_ _11036_ _10067_ VGND VGND VPWR VPWR _00259_
+ sky130_fd_sc_hd__o211a_1
X_13488_ _05477_ _05480_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__nor2_1
X_16276_ net458 net507 VGND VGND VPWR VPWR _08367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18015_ _09998_ _09999_ VGND VGND VPWR VPWR _10000_ sky130_fd_sc_hd__and2b_1
XFILLER_0_180_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15227_ _07304_ _07319_ _07243_ _07241_ VGND VGND VPWR VPWR _07326_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15158_ _07204_ _07205_ VGND VGND VPWR VPWR _07257_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14109_ net24 _05489_ _05491_ net1030 VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__and4b_1
XFILLER_0_22_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19966_ _11517_ _11834_ net181 VGND VGND VPWR VPWR _11835_ sky130_fd_sc_hd__a21o_1
Xfanout109 net110 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_4
X_15089_ net535 net462 VGND VGND VPWR VPWR _07188_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18917_ _10847_ _10891_ VGND VGND VPWR VPWR _10892_ sky130_fd_sc_hd__xnor2_1
X_19897_ _11742_ _11753_ _11765_ _11770_ VGND VGND VPWR VPWR _11771_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18848_ _10821_ _10822_ _10823_ VGND VGND VPWR VPWR _10824_ sky130_fd_sc_hd__nand3_2
XFILLER_0_59_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18779_ top0.pid_d.curr_int\[9\] VGND VGND VPWR VPWR _10756_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20810_ _11571_ _12656_ _12658_ VGND VGND VPWR VPWR _12659_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_85_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_85_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21790_ _01350_ _01351_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__xor2_1
XFILLER_0_166_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20741_ net301 _11525_ _12551_ VGND VGND VPWR VPWR _12590_ sky130_fd_sc_hd__or3_1
XFILLER_0_147_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23460_ _11651_ net85 _02893_ _02894_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__a211o_1
XFILLER_0_18_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20672_ net249 _12499_ _12490_ VGND VGND VPWR VPWR _12521_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22411_ _01967_ _01968_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23391_ net111 _11784_ _02830_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__or3_1
XFILLER_0_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25130_ _03343_ _04182_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22342_ net97 _01900_ net78 VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_171_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25061_ _04370_ _04373_ _04409_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_143_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22273_ _01135_ _01412_ _01113_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24012_ _03253_ _03369_ _03323_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__a21oi_1
Xhold130 top0.svm0.tA\[0\] VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__dlygate4sd3_1
X_21224_ _12626_ VGND VGND VPWR VPWR _13068_ sky130_fd_sc_hd__inv_2
Xhold141 top0.matmul0.matmul_stage_inst.c\[12\] VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 top0.svm0.tC\[1\] VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 top0.cordic0.cos\[13\] VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 top0.pid_d.prev_error\[10\] VGND VGND VPWR VPWR net874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 top0.pid_q.curr_error\[15\] VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__dlygate4sd3_1
X_21155_ _12921_ _12931_ _12999_ VGND VGND VPWR VPWR _13000_ sky130_fd_sc_hd__a21o_1
Xhold196 top0.svm0.delta\[2\] VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 net630 VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__clkbuf_4
Xfanout621 net624 VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__clkbuf_4
X_20106_ _11964_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__clkbuf_1
Xfanout632 net634 VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__clkbuf_4
X_25963_ _05172_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__clkbuf_1
Xfanout643 net645 VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__clkbuf_2
X_21086_ _12921_ _12931_ VGND VGND VPWR VPWR _12932_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout654 net687 VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__buf_2
Xfanout665 net666 VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__clkbuf_4
Xfanout676 net686 VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__clkbuf_4
X_24914_ _04206_ _04208_ _04203_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__a21o_1
X_20037_ _11632_ top0.cordic0.gm0.iter\[2\] VGND VGND VPWR VPWR _11901_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout687 net2 VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__clkbuf_8
X_25894_ net430 _05438_ _05104_ _05110_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__nand4_1
Xfanout698 net699 VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24845_ _04096_ _04102_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24776_ _03572_ _04040_ _04042_ VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21988_ net127 net124 VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26515_ clknet_leaf_66_clk_sys _00138_ net659 VGND VGND VPWR VPWR top0.pid_q.out\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_23727_ _03042_ _03052_ _03044_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__a21oi_1
X_20939_ _12785_ _12683_ VGND VGND VPWR VPWR _12787_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14460_ _06596_ _06594_ _06664_ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__and3_1
X_26446_ clknet_leaf_59_clk_sys _00087_ net644 VGND VGND VPWR VPWR top0.kiq\[3\] sky130_fd_sc_hd__dfrtp_1
X_23658_ net565 net557 top0.matmul0.matmul_stage_inst.e\[2\] VGND VGND VPWR VPWR _03016_
+ sky130_fd_sc_hd__o21a_4
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13411_ _05608_ _05609_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__nor2_2
XFILLER_0_138_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14391_ _06501_ _06504_ _06599_ VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_3_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22609_ _02153_ _02162_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__xor2_2
XFILLER_0_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23589_ _02961_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26377_ _05420_ VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13342_ _05522_ _05525_ _05554_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__a21o_1
X_16130_ _08220_ _08222_ VGND VGND VPWR VPWR _08223_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_51_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25328_ _04669_ _04672_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13273_ _05485_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__buf_2
X_16061_ _08063_ _08066_ _08154_ VGND VGND VPWR VPWR _08155_ sky130_fd_sc_hd__o21ai_2
X_25259_ _04605_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__clkbuf_1
X_15012_ _07131_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__clkbuf_1
X_19820_ net175 _11689_ _11698_ _11699_ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19751_ _11632_ _11553_ _11633_ net83 VGND VGND VPWR VPWR _11634_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_75_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16963_ top0.pid_q.prev_error\[10\] top0.pid_q.curr_error\[10\] VGND VGND VPWR VPWR
+ _09020_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18702_ net432 _10598_ _10599_ _10679_ net437 VGND VGND VPWR VPWR _10680_ sky130_fd_sc_hd__a32o_1
X_15914_ _08007_ _08008_ VGND VGND VPWR VPWR _08009_ sky130_fd_sc_hd__xnor2_1
X_19682_ net1014 _11568_ net174 VGND VGND VPWR VPWR _11569_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_194_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16894_ net546 _08949_ _08955_ _08882_ VGND VGND VPWR VPWR _08956_ sky130_fd_sc_hd__a211o_1
XFILLER_0_189_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18633_ net381 _10203_ _09364_ VGND VGND VPWR VPWR _10611_ sky130_fd_sc_hd__o21ai_1
X_15845_ _07939_ _07940_ VGND VGND VPWR VPWR _07941_ sky130_fd_sc_hd__xor2_1
XFILLER_0_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18564_ _10465_ _10467_ _10542_ VGND VGND VPWR VPWR _10543_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15776_ _07727_ _07728_ _07872_ VGND VGND VPWR VPWR _07873_ sky130_fd_sc_hd__a21oi_2
X_17515_ net352 _09501_ VGND VGND VPWR VPWR _09502_ sky130_fd_sc_hd__nand2_1
X_14727_ _05629_ _06832_ _05640_ _06320_ VGND VGND VPWR VPWR _06930_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18495_ _10473_ _10474_ VGND VGND VPWR VPWR _10475_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17446_ net396 net391 VGND VGND VPWR VPWR _09433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14658_ _06551_ _06807_ _06819_ _06858_ _06816_ VGND VGND VPWR VPWR _06862_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13609_ _05534_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__buf_6
X_17377_ _09363_ VGND VGND VPWR VPWR _09364_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14589_ _06740_ _06793_ _06794_ VGND VGND VPWR VPWR _06795_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19116_ net432 top0.pid_d.out\[14\] top0.pid_d.curr_int\[14\] _11084_ _07137_ VGND
+ VGND VPWR VPWR _11088_ sky130_fd_sc_hd__a41o_1
XFILLER_0_171_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16328_ net1028 net446 VGND VGND VPWR VPWR _08418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19047_ net309 _10942_ _11018_ _10690_ VGND VGND VPWR VPWR _11020_ sky130_fd_sc_hd__a211o_1
X_16259_ _08255_ _08257_ _08349_ VGND VGND VPWR VPWR _08350_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19949_ top0.cordic0.slte0.opA\[1\] _11818_ _11819_ _11817_ VGND VGND VPWR VPWR _00361_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22960_ _02470_ _02471_ _02331_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21911_ _01472_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__inv_2
X_22891_ top0.svm0.tC\[10\] VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__inv_2
X_24630_ _03765_ _03164_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__nor2_1
X_21842_ _01389_ _01397_ _01403_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__nand3_1
XFILLER_0_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24561_ _03767_ _03772_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__or2_1
XFILLER_0_188_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21773_ _01334_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26300_ spi0.data_packed\[48\] spi0.data_packed\[49\] net697 VGND VGND VPWR VPWR
+ _05382_ sky130_fd_sc_hd__mux2_1
X_20724_ _12572_ _12564_ _12565_ VGND VGND VPWR VPWR _12573_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23512_ _02921_ VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__clkbuf_1
X_24492_ _03663_ _03676_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27280_ clknet_3_1__leaf_clk_mosi _00894_ VGND VGND VPWR VPWR spi0.data_packed\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23443_ _02865_ _02866_ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__nor2_1
X_26231_ _05347_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__clkbuf_1
X_20655_ net270 net280 net287 VGND VGND VPWR VPWR _12504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23374_ net125 _02791_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__xnor2_1
X_26162_ _05302_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__clkbuf_1
X_20586_ _12428_ _12433_ _12434_ VGND VGND VPWR VPWR _12435_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25113_ _04387_ _04389_ _04381_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__a21o_1
X_22325_ _01805_ _01807_ _01873_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26093_ top0.matmul0.alpha_pass\[15\] _05168_ _05271_ VGND VGND VPWR VPWR _05272_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25044_ _04303_ _04393_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__nand2_1
X_22256_ _01113_ _01768_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21207_ _13050_ VGND VGND VPWR VPWR _13051_ sky130_fd_sc_hd__inv_2
XFILLER_0_197_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22187_ _01706_ _01746_ _01747_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_100_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21138_ _11689_ net246 VGND VGND VPWR VPWR _12983_ sky130_fd_sc_hd__nor2_1
X_26995_ clknet_leaf_23_clk_sys _00612_ net625 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout440 top0.pid_d.state\[2\] VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__clkbuf_2
Xfanout451 top0.pid_q.mult0.b\[12\] VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__clkbuf_4
Xfanout462 top0.pid_q.mult0.b\[8\] VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__clkbuf_4
X_13960_ _05795_ _05789_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__or2_1
Xfanout473 net474 VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__clkbuf_4
X_25946_ net428 _05155_ _05158_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__a21o_1
X_21069_ _11672_ net251 VGND VGND VPWR VPWR _12915_ sky130_fd_sc_hd__nor2_1
Xfanout484 net486 VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__buf_2
Xfanout495 net496 VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13891_ net22 _05683_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__nand2_2
X_25877_ top0.matmul0.beta_pass\[8\] _05095_ _05093_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__o21a_1
X_15630_ net505 net492 VGND VGND VPWR VPWR _07728_ sky130_fd_sc_hd__nand2_1
X_24828_ _03564_ _03826_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__nand2_2
XFILLER_0_154_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15561_ _07636_ _07659_ VGND VGND VPWR VPWR _07660_ sky130_fd_sc_hd__xnor2_2
X_24759_ _04021_ _04022_ _04023_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17300_ top0.matmul0.matmul_stage_inst.mult1\[8\] top0.matmul0.matmul_stage_inst.mult2\[8\]
+ VGND VGND VPWR VPWR _09295_ sky130_fd_sc_hd__xor2_1
XFILLER_0_28_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14512_ _06217_ _05579_ _06718_ _06106_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__o22a_1
XFILLER_0_167_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18280_ net402 net314 VGND VGND VPWR VPWR _10262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15492_ _07293_ _07296_ VGND VGND VPWR VPWR _07591_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17231_ net546 _08853_ VGND VGND VPWR VPWR _09236_ sky130_fd_sc_hd__or2_1
XFILLER_0_193_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14443_ _06638_ _06650_ VGND VGND VPWR VPWR _06651_ sky130_fd_sc_hd__xor2_2
X_26429_ clknet_leaf_77_clk_sys _00070_ net631 VGND VGND VPWR VPWR top0.kid\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout80 net81 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_153_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout91 net92 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
X_17162_ top0.pid_q.curr_int\[5\] _09141_ _09175_ _09136_ VGND VGND VPWR VPWR _00218_
+ sky130_fd_sc_hd__a22o_1
X_14374_ _06217_ _05822_ VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__nor2_2
XFILLER_0_182_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16113_ _08100_ _08102_ _08101_ VGND VGND VPWR VPWR _08206_ sky130_fd_sc_hd__o21a_1
X_13325_ _05537_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_33_clk_sys clknet_3_6__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_33_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_17093_ top0.pid_q.curr_error\[5\] _00011_ _09117_ VGND VGND VPWR VPWR _09123_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16044_ _08039_ _08059_ VGND VGND VPWR VPWR _08138_ sky130_fd_sc_hd__nor2_1
X_13256_ net173 top0.svm0.state\[0\] top0.svm0.state\[1\] VGND VGND VPWR VPWR _05469_
+ sky130_fd_sc_hd__nor3b_4
XFILLER_0_161_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19803_ _11680_ _11683_ VGND VGND VPWR VPWR _11684_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17995_ _09980_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16946_ _09003_ _08990_ top0.pid_q.prev_error\[8\] VGND VGND VPWR VPWR _09004_ sky130_fd_sc_hd__o21ba_1
X_19734_ _11512_ _11617_ VGND VGND VPWR VPWR _11618_ sky130_fd_sc_hd__nand2_2
XFILLER_0_159_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19665_ _11544_ _11551_ VGND VGND VPWR VPWR _11552_ sky130_fd_sc_hd__nand2_1
X_16877_ top0.pid_q.prev_error\[4\] top0.pid_q.curr_error\[4\] VGND VGND VPWR VPWR
+ _08940_ sky130_fd_sc_hd__xor2_1
X_18616_ top0.pid_d.curr_int\[8\] VGND VGND VPWR VPWR _10594_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15828_ _07921_ _07923_ VGND VGND VPWR VPWR _07924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19596_ top0.cordic0.slte0.opB\[8\] VGND VGND VPWR VPWR _11485_ sky130_fd_sc_hd__inv_2
X_18547_ _10524_ _10525_ VGND VGND VPWR VPWR _10526_ sky130_fd_sc_hd__xor2_1
X_15759_ _07739_ _07740_ _07741_ VGND VGND VPWR VPWR _07856_ sky130_fd_sc_hd__o21a_1
XFILLER_0_176_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18478_ net344 net348 VGND VGND VPWR VPWR _10458_ sky130_fd_sc_hd__and2_2
XFILLER_0_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17429_ net403 net347 VGND VGND VPWR VPWR _09416_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20440_ _11407_ net301 net275 VGND VGND VPWR VPWR _12289_ sky130_fd_sc_hd__or3_1
XFILLER_0_160_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20371_ _12049_ _12131_ _12127_ _12128_ VGND VGND VPWR VPWR _12220_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_67_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22110_ _01318_ _01669_ _01670_ _01590_ _01671_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__o221a_1
XFILLER_0_43_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23090_ _02541_ _02590_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22041_ _01262_ _01601_ _01602_ net106 net122 VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_11_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25800_ _12009_ _02282_ _12012_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__a21o_2
XFILLER_0_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26780_ clknet_leaf_109_clk_sys _00397_ net579 VGND VGND VPWR VPWR top0.cordic0.sin\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_23992_ _03345_ _03349_ VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_199_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25731_ top0.matmul0.sin\[10\] _04942_ net73 VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__o21ai_1
X_22943_ _02455_ _02456_ _02339_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__mux2_1
X_25662_ _04913_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__clkbuf_4
X_22874_ _02367_ top0.svm0.tB\[8\] _02391_ _02392_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24613_ _03887_ _03895_ _03966_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__o21a_1
X_21825_ net121 _01377_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__nand2_2
X_25593_ _04884_ _04886_ _04846_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24544_ _03879_ _03898_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__xnor2_4
X_21756_ _01285_ _01317_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__xnor2_2
X_20707_ net285 _11608_ VGND VGND VPWR VPWR _12556_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27263_ clknet_3_6__leaf_clk_mosi _00877_ VGND VGND VPWR VPWR spi0.data_packed\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_24475_ _03826_ _03830_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__xnor2_1
X_21687_ _01213_ _01248_ _01163_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__or3b_2
XPHY_EDGE_ROW_199_Left_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26214_ spi0.data_packed\[5\] spi0.data_packed\[6\] net694 VGND VGND VPWR VPWR _05339_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20638_ _12460_ _12461_ _12476_ _12486_ VGND VGND VPWR VPWR _12487_ sky130_fd_sc_hd__a31o_1
X_23426_ net98 _11783_ _02862_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__or3_1
XFILLER_0_191_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27194_ clknet_leaf_56_clk_sys _00808_ net666 VGND VGND VPWR VPWR top0.currT_r\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23357_ _02785_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__inv_2
X_26145_ spi0.data_packed\[0\] spi0.data_packed\[15\] spi0.data_packed\[1\] net19
+ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__a31o_1
XFILLER_0_184_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20569_ _12416_ _12417_ _12408_ VGND VGND VPWR VPWR _12418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22308_ _01796_ _01801_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__nor2_1
X_14090_ _06300_ _06301_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__nor2_2
XFILLER_0_15_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23288_ _11649_ _02735_ _11954_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__a21o_1
X_26076_ top0.pid_d.out\[11\] _05232_ _05233_ spi0.data_packed\[75\] VGND VGND VPWR
+ VPWR _05259_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25027_ _04361_ _04376_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__xnor2_1
X_22239_ _01224_ _01798_ _01799_ net80 VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16800_ net515 _08856_ _08859_ net734 _08873_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__a221o_1
X_17780_ _09761_ _09766_ VGND VGND VPWR VPWR _09767_ sky130_fd_sc_hd__xnor2_2
X_26978_ clknet_leaf_25_clk_sys _00595_ net628 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_14992_ spi0.data_packed\[2\] top0.periodTop\[2\] _07108_ VGND VGND VPWR VPWR _07121_
+ sky130_fd_sc_hd__mux2_1
Xfanout270 top0.cordic0.vec\[0\]\[6\] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_191_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout281 net284 VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__clkbuf_2
X_16731_ _08654_ _08813_ _08814_ net459 VGND VGND VPWR VPWR _08815_ sky130_fd_sc_hd__a2bb2o_1
Xfanout292 net293 VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__buf_4
X_13943_ _05779_ _05781_ _05777_ VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__a21bo_1
X_25929_ _05437_ _05140_ _05138_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_202_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19450_ _11345_ _11346_ VGND VGND VPWR VPWR _11348_ sky130_fd_sc_hd__or2_1
X_16662_ _08692_ _08725_ _08726_ VGND VGND VPWR VPWR _08747_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13874_ _05763_ _05768_ _05760_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_198_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18401_ _10271_ _10273_ _10272_ VGND VGND VPWR VPWR _10382_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15613_ _07694_ VGND VGND VPWR VPWR _07711_ sky130_fd_sc_hd__inv_2
X_19381_ top0.pid_d.prev_error\[14\] _11284_ _11287_ net765 VGND VGND VPWR VPWR _00324_
+ sky130_fd_sc_hd__a22o_1
X_16593_ net549 net13 _08679_ VGND VGND VPWR VPWR _08680_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18332_ _10310_ _10313_ net416 VGND VGND VPWR VPWR _10314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15544_ _07576_ _07577_ _07578_ VGND VGND VPWR VPWR _07643_ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18263_ top0.pid_d.curr_int\[4\] _10159_ top0.pid_d.out\[4\] VGND VGND VPWR VPWR
+ _10245_ sky130_fd_sc_hd__a21o_1
X_15475_ _07572_ _07573_ VGND VGND VPWR VPWR _07574_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_189_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17214_ top0.pid_q.curr_int\[11\] _09141_ _09220_ _09136_ _09221_ VGND VGND VPWR
+ VPWR _00224_ sky130_fd_sc_hd__a221o_1
X_14426_ _06587_ _06589_ _06633_ VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18194_ net325 net394 VGND VGND VPWR VPWR _10177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17145_ net553 _09159_ _09160_ net548 _08928_ VGND VGND VPWR VPWR _09161_ sky130_fd_sc_hd__a32o_1
X_14357_ _06495_ _06497_ _06496_ VGND VGND VPWR VPWR _06566_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_4_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13308_ _05476_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__buf_2
X_17076_ net865 _09100_ _09102_ _09070_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__a22o_1
X_14288_ _06496_ _06497_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16027_ _08106_ _08120_ VGND VGND VPWR VPWR _08121_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13239_ _05455_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17978_ _09861_ _09962_ _09963_ VGND VGND VPWR VPWR _09964_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16929_ top0.pid_q.curr_error\[7\] VGND VGND VPWR VPWR _08988_ sky130_fd_sc_hd__inv_2
X_19717_ _11600_ _11601_ VGND VGND VPWR VPWR _11602_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19648_ net116 net111 net108 net103 net199 net193 VGND VGND VPWR VPWR _11536_ sky130_fd_sc_hd__mux4_1
XFILLER_0_189_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19579_ _11464_ _11465_ _11466_ _11467_ VGND VGND VPWR VPWR _11468_ sky130_fd_sc_hd__or4_1
XFILLER_0_172_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21610_ _01130_ _01171_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22590_ _02112_ _01924_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21541_ _01102_ net139 VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24260_ _03539_ _03615_ _03617_ _03449_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_44_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21472_ _01033_ _01036_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__or2_1
X_23211_ _01320_ net1013 _02660_ _02662_ VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__a31o_1
X_20423_ net304 net299 VGND VGND VPWR VPWR _12272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24191_ top0.matmul0.matmul_stage_inst.f\[0\] _03146_ _03148_ top0.matmul0.matmul_stage_inst.e\[0\]
+ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__a22o_4
XFILLER_0_44_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23142_ _02629_ _02630_ top0.svm0.delta\[13\] VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__mux2_1
X_20354_ _11672_ _12126_ _12201_ _12202_ _12043_ VGND VGND VPWR VPWR _12203_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23073_ net61 top0.svm0.counter\[2\] VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20285_ net252 net246 VGND VGND VPWR VPWR _12134_ sky130_fd_sc_hd__nor2b_2
X_22024_ _01281_ _01582_ _01583_ net145 _01585_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__a2111o_1
X_26901_ clknet_leaf_108_clk_sys _00518_ net585 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold12 top0.cordic0.sin\[3\] VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__dlygate4sd3_1
X_26832_ clknet_leaf_42_clk_sys _00449_ net684 VGND VGND VPWR VPWR top0.svm0.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold23 _00325_ VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 top0.kpq\[9\] VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 top0.cordic0.sin\[0\] VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 top0.cordic0.cos\[2\] VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 top0.matmul0.matmul_stage_inst.a\[5\] VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 top0.matmul0.matmul_stage_inst.b\[14\] VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__dlygate4sd3_1
X_26763_ clknet_leaf_87_clk_sys _00380_ net645 VGND VGND VPWR VPWR top0.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23975_ _03267_ _03268_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__xnor2_1
Xhold89 top0.kpq\[3\] VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__dlygate4sd3_1
X_25714_ top0.matmul0.sin\[5\] _04973_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22926_ _02438_ _02441_ _02352_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26694_ clknet_leaf_71_clk_sys _00311_ net657 VGND VGND VPWR VPWR top0.pid_d.prev_error\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25645_ _04920_ _04921_ net69 VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__o21ai_1
X_22857_ top0.svm0.tA\[14\] _02375_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21808_ _01368_ _01369_ _01267_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13590_ _05647_ _05802_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25576_ _04875_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__clkbuf_1
X_22788_ _05719_ _05717_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24527_ _03199_ _03880_ _03881_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__o21ai_4
X_21739_ _01300_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15260_ net1026 net487 VGND VGND VPWR VPWR _07359_ sky130_fd_sc_hd__nand2_1
X_27246_ clknet_3_0__leaf_clk_mosi _00860_ VGND VGND VPWR VPWR spi0.data_packed\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24458_ _03797_ _03813_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__xnor2_2
X_14211_ _05504_ _05538_ _05539_ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__nor3_1
XFILLER_0_136_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23409_ net216 _02663_ _11730_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15191_ net540 net454 VGND VGND VPWR VPWR _07290_ sky130_fd_sc_hd__nand2_2
X_27177_ clknet_leaf_88_clk_sys _00791_ net643 VGND VGND VPWR VPWR top0.periodTop_r\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_24389_ _03160_ _03165_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_9 net1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14142_ _06135_ _06350_ _06352_ _06353_ net60 VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__o221a_1
X_26128_ spi0.data_packed\[23\] _05281_ _05282_ net962 VGND VGND VPWR VPWR _00804_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14073_ _06281_ _06284_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__xnor2_4
X_18950_ _10751_ _10840_ _10829_ _10752_ VGND VGND VPWR VPWR _10924_ sky130_fd_sc_hd__o211a_1
X_26059_ _05246_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__clkbuf_1
X_17901_ _09807_ _09886_ _09887_ VGND VGND VPWR VPWR _09888_ sky130_fd_sc_hd__o21a_1
X_18881_ _10854_ _10855_ VGND VGND VPWR VPWR _10856_ sky130_fd_sc_hd__xnor2_1
X_17832_ _09686_ _09818_ _09714_ VGND VGND VPWR VPWR _09819_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17763_ _09515_ _09749_ _09742_ VGND VGND VPWR VPWR _09750_ sky130_fd_sc_hd__o21a_1
X_14975_ spi0.data_packed\[29\] top0.kiq\[13\] _07108_ VGND VGND VPWR VPWR _07110_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16714_ _08747_ _08782_ _08746_ VGND VGND VPWR VPWR _08798_ sky130_fd_sc_hd__o21a_1
X_19502_ _11390_ _11393_ VGND VGND VPWR VPWR _11394_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13926_ net51 _05602_ _05603_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__and3_2
X_17694_ _09677_ _09680_ VGND VGND VPWR VPWR _09681_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19433_ net431 _10423_ _11332_ net442 _11179_ VGND VGND VPWR VPWR _11333_ sky130_fd_sc_hd__a221o_1
X_16645_ _08664_ _08730_ VGND VGND VPWR VPWR _08731_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13857_ _06036_ _06038_ _06066_ _06067_ _06069_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19364_ _11284_ _00006_ VGND VGND VPWR VPWR _11286_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_202_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16576_ _08526_ _08584_ _08534_ VGND VGND VPWR VPWR _08663_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_201_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13788_ _05974_ _05975_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18315_ _10291_ _10296_ VGND VGND VPWR VPWR _10297_ sky130_fd_sc_hd__xnor2_2
X_15527_ net470 net520 VGND VGND VPWR VPWR _07626_ sky130_fd_sc_hd__nand2_1
X_19295_ top0.pid_d.prev_error\[11\] top0.pid_d.curr_error\[11\] VGND VGND VPWR VPWR
+ _11237_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18246_ net421 _10228_ net416 net411 VGND VGND VPWR VPWR _10229_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_199_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15458_ net485 net511 VGND VGND VPWR VPWR _07557_ sky130_fd_sc_hd__nand2_2
XFILLER_0_154_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14409_ net44 _05666_ VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__nand2_2
XFILLER_0_128_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18177_ top0.pid_d.out\[4\] top0.pid_d.curr_int\[4\] VGND VGND VPWR VPWR _10160_
+ sky130_fd_sc_hd__xnor2_1
X_15389_ _07482_ _07486_ _07487_ VGND VGND VPWR VPWR _07488_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_163_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17128_ net543 _07795_ _09145_ VGND VGND VPWR VPWR _09146_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17059_ top0.pid_q.curr_error\[5\] _09100_ _09102_ _08949_ VGND VGND VPWR VPWR _00186_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20070_ _11930_ _11924_ _11925_ VGND VGND VPWR VPWR _11932_ sky130_fd_sc_hd__or3_1
XFILLER_0_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23760_ _03116_ _03117_ VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_135_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20972_ _11726_ net230 VGND VGND VPWR VPWR _12819_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22711_ _02260_ _02261_ _02182_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__mux2_1
X_23691_ _03024_ _03025_ _03015_ _03016_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__o22a_2
XFILLER_0_95_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25430_ _04516_ _04770_ _04772_ _04406_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22642_ net79 _01248_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25361_ _04612_ _04704_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22573_ _02045_ _02085_ _02007_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27100_ clknet_leaf_16_clk_sys _00717_ net611 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.a\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_24312_ _03130_ _03135_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21524_ _01063_ _01064_ _01067_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__nor3_1
X_25292_ _04626_ _04637_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_173_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27031_ clknet_leaf_15_clk_sys _00648_ net614 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24243_ _03558_ _03570_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21455_ _00988_ _01012_ _01019_ _00966_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_69_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20406_ net277 net271 VGND VGND VPWR VPWR _12255_ sky130_fd_sc_hd__nand2_1
X_24174_ _03409_ _03410_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__nor2_1
X_21386_ _00932_ _00953_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23125_ top0.svm0.delta\[9\] _02617_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__xnor2_1
X_20337_ _12174_ _12179_ _12184_ _12185_ _12161_ VGND VGND VPWR VPWR _12186_ sky130_fd_sc_hd__o311a_1
X_23056_ top0.periodTop_r\[4\] _02539_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__nor2_1
X_20268_ _12115_ _12116_ VGND VGND VPWR VPWR _12117_ sky130_fd_sc_hd__nor2_1
X_22007_ net166 _01512_ _01311_ _01442_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_179_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20199_ net269 net283 VGND VGND VPWR VPWR _12048_ sky130_fd_sc_hd__or2b_1
XFILLER_0_179_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26815_ clknet_leaf_55_clk_sys _00432_ net667 VGND VGND VPWR VPWR top0.pid_q.prev_int\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14760_ _06921_ _06922_ VGND VGND VPWR VPWR _06962_ sky130_fd_sc_hd__nor2_1
X_26746_ clknet_leaf_97_clk_sys _00363_ net588 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23958_ _03313_ _03315_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__nand2_2
X_13711_ _05922_ _05923_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22909_ _02345_ top0.svm0.tC\[11\] _02425_ _02426_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__o22a_1
X_14691_ _06839_ _06844_ _06894_ VGND VGND VPWR VPWR _06895_ sky130_fd_sc_hd__a21o_1
XFILLER_0_169_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26677_ clknet_leaf_64_clk_sys _00294_ net656 VGND VGND VPWR VPWR top0.pid_d.curr_error\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_23889_ _03237_ _03242_ _03246_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16430_ _08513_ _08518_ VGND VGND VPWR VPWR _08519_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13642_ _05803_ _05853_ _05854_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__a21bo_1
X_25628_ net69 top0.matmul0.sin\[1\] VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16361_ net497 _08447_ _08450_ VGND VGND VPWR VPWR _08451_ sky130_fd_sc_hd__nand3_1
XFILLER_0_184_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13573_ _05754_ _05755_ _05785_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__a21oi_1
X_25559_ _04866_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18100_ _10082_ _10083_ VGND VGND VPWR VPWR _10084_ sky130_fd_sc_hd__xor2_1
X_15312_ net527 net495 VGND VGND VPWR VPWR _07411_ sky130_fd_sc_hd__nand2_1
X_19080_ net307 _11051_ VGND VGND VPWR VPWR _11052_ sky130_fd_sc_hd__nand2_1
X_16292_ _08296_ _08300_ _08382_ VGND VGND VPWR VPWR _08383_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18031_ net335 net389 VGND VGND VPWR VPWR _10016_ sky130_fd_sc_hd__nand2_2
XFILLER_0_152_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15243_ _07243_ _07341_ VGND VGND VPWR VPWR _07342_ sky130_fd_sc_hd__xnor2_1
X_27229_ clknet_3_1__leaf_clk_mosi _00843_ VGND VGND VPWR VPWR spi0.data_packed\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_169_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15174_ _07198_ _07199_ _07272_ VGND VGND VPWR VPWR _07273_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_136_Left_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14125_ _06332_ _06334_ _06335_ _06336_ VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__o22a_1
XFILLER_0_127_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19982_ net184 _11844_ _11849_ net181 _11808_ VGND VGND VPWR VPWR _11850_ sky130_fd_sc_hd__a2111oi_1
X_14056_ net65 _06268_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__nand2_1
X_18933_ _10841_ _10905_ _10907_ VGND VGND VPWR VPWR _10908_ sky130_fd_sc_hd__nor3_1
XFILLER_0_24_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18864_ _10832_ _10839_ _07710_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__o21a_1
XFILLER_0_197_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17815_ _09798_ _09801_ VGND VGND VPWR VPWR _09802_ sky130_fd_sc_hd__xnor2_1
X_18795_ _10456_ _10720_ VGND VGND VPWR VPWR _10771_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17746_ _09727_ _09732_ _09492_ VGND VGND VPWR VPWR _09733_ sky130_fd_sc_hd__o21a_1
XFILLER_0_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14958_ spi0.data_packed\[21\] top0.kiq\[5\] _07097_ VGND VGND VPWR VPWR _07101_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_145_Left_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13909_ _05772_ _05783_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__or2_1
XFILLER_0_159_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17677_ _09654_ _09613_ _09610_ VGND VGND VPWR VPWR _09664_ sky130_fd_sc_hd__mux2_1
X_14889_ spi0.data_packed\[52\] top0.kpq\[4\] _07064_ VGND VGND VPWR VPWR _07065_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16628_ _08709_ _08712_ VGND VGND VPWR VPWR _08714_ sky130_fd_sc_hd__nand2_1
X_19416_ top0.pid_d.prev_int\[3\] _11311_ _11317_ VGND VGND VPWR VPWR _11318_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16559_ _08554_ _08555_ _08556_ VGND VGND VPWR VPWR _08646_ sky130_fd_sc_hd__o21a_1
X_19347_ top0.pid_d.curr_error\[5\] _11275_ _11279_ _11171_ VGND VGND VPWR VPWR _00299_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19278_ top0.matmul0.alpha_pass\[10\] _11210_ VGND VGND VPWR VPWR _11222_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18229_ _10210_ _10211_ VGND VGND VPWR VPWR _10212_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_154_Left_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21240_ _12642_ _13081_ _13080_ _12609_ VGND VGND VPWR VPWR _13084_ sky130_fd_sc_hd__a211o_1
XFILLER_0_41_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_81_clk_sys clknet_3_4__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_81_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
Xhold301 top0.cordic0.sin\[8\] VGND VGND VPWR VPWR net1001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21171_ net1021 _13014_ VGND VGND VPWR VPWR _13015_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20122_ net212 _11976_ _11978_ VGND VGND VPWR VPWR _11979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24930_ _03343_ _04190_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__nor2_1
X_20053_ _11902_ _11518_ _11657_ VGND VGND VPWR VPWR _11916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24861_ _04118_ _04119_ _04105_ _04106_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_163_Left_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26600_ clknet_leaf_67_clk_sys _00223_ net661 VGND VGND VPWR VPWR top0.pid_q.curr_int\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_23812_ _03014_ _03033_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__or2_1
X_24792_ _03940_ _03941_ _03830_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__a21o_1
XFILLER_0_197_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26531_ clknet_leaf_61_clk_sys _00154_ net651 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_23743_ _03087_ _03100_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__nand2_1
X_20955_ _12749_ _12802_ VGND VGND VPWR VPWR _12803_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26462_ clknet_leaf_11_clk_sys _00014_ net601 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_23674_ _03026_ _03031_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__xor2_1
XFILLER_0_178_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20886_ _12161_ _12187_ _12194_ _12732_ _12734_ VGND VGND VPWR VPWR _12735_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_177_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25413_ _04664_ _04755_ _04756_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_166_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22625_ _02177_ _02178_ _12740_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__a21oi_1
X_26393_ clknet_leaf_37_clk_sys _00034_ net679 VGND VGND VPWR VPWR top0.svm0.tC\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25344_ _04685_ _04688_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__xor2_1
X_22556_ _02109_ _02110_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_172_Left_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21507_ net115 net97 VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__xnor2_4
X_25275_ _03900_ _04272_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22487_ _02036_ _02043_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_185_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27014_ clknet_leaf_24_clk_sys _00631_ net626 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_24226_ _03565_ _03583_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__xor2_1
XFILLER_0_107_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21438_ _00968_ _00982_ _01003_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24157_ _03509_ _03514_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__xnor2_1
X_21369_ net236 _13001_ _13174_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__o21ai_1
X_23108_ _02596_ _02605_ _02458_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__a21oi_1
X_24088_ _03442_ _03445_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__xor2_2
X_15930_ _08019_ _08024_ VGND VGND VPWR VPWR _08025_ sky130_fd_sc_hd__xnor2_1
X_23039_ net54 net52 net49 _02539_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_181_Left_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15861_ _07954_ _07956_ VGND VGND VPWR VPWR _07957_ sky130_fd_sc_hd__xnor2_1
X_17600_ net345 net426 _09585_ VGND VGND VPWR VPWR _09587_ sky130_fd_sc_hd__a21oi_1
X_14812_ _07010_ _07011_ _06978_ VGND VGND VPWR VPWR _07012_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_157_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18580_ _10536_ _10558_ VGND VGND VPWR VPWR _10559_ sky130_fd_sc_hd__xnor2_4
X_15792_ _07718_ _07776_ _07775_ VGND VGND VPWR VPWR _07889_ sky130_fd_sc_hd__o21ba_1
X_17531_ _09355_ _09395_ VGND VGND VPWR VPWR _09518_ sky130_fd_sc_hd__nor2_4
X_14743_ net807 _06279_ _06945_ _05465_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26729_ clknet_leaf_104_clk_sys _00346_ net576 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_54_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17462_ _09368_ _09446_ _09406_ VGND VGND VPWR VPWR _09449_ sky130_fd_sc_hd__or3b_1
X_14674_ _06876_ _06877_ VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__xor2_1
XFILLER_0_74_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16413_ net447 net1029 VGND VGND VPWR VPWR _08502_ sky130_fd_sc_hd__nand2_1
X_19201_ _11120_ _11150_ _11151_ VGND VGND VPWR VPWR _11152_ sky130_fd_sc_hd__and3_1
X_13625_ _05834_ _05835_ _05837_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__and3_1
X_17393_ net419 net337 VGND VGND VPWR VPWR _09380_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_190_Left_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19132_ top0.pid_d.mult0.a\[0\] _11096_ _11101_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__a21o_1
X_16344_ _08430_ _08433_ VGND VGND VPWR VPWR _08434_ sky130_fd_sc_hd__xnor2_2
X_13556_ _05763_ _05768_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19063_ net435 _11031_ _11035_ net432 _07138_ VGND VGND VPWR VPWR _11036_ sky130_fd_sc_hd__a221o_1
X_16275_ net463 net503 VGND VGND VPWR VPWR _08366_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13487_ _05696_ _05699_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__xor2_2
XFILLER_0_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18014_ _09992_ _09997_ VGND VGND VPWR VPWR _09999_ sky130_fd_sc_hd__nand2_1
X_15226_ _07304_ _07319_ _07324_ VGND VGND VPWR VPWR _07325_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15157_ _07204_ _07205_ VGND VGND VPWR VPWR _07256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14108_ net25 net20 VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__and2_2
XFILLER_0_129_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19965_ net195 net185 net189 net201 VGND VGND VPWR VPWR _11834_ sky130_fd_sc_hd__a31o_1
X_15088_ net537 net460 VGND VGND VPWR VPWR _07187_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14039_ _06242_ _06250_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__nand2_1
X_18916_ _10857_ _10890_ VGND VGND VPWR VPWR _10891_ sky130_fd_sc_hd__xor2_1
X_19896_ net228 _11764_ VGND VGND VPWR VPWR _11770_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18847_ _10738_ _10739_ VGND VGND VPWR VPWR _10823_ sky130_fd_sc_hd__or2_1
X_18778_ top0.pid_d.out\[10\] _07137_ VGND VGND VPWR VPWR _10755_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_28_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_28_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17729_ _09686_ _09714_ _09715_ VGND VGND VPWR VPWR _09716_ sky130_fd_sc_hd__or3_1
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20740_ _12587_ _12588_ VGND VGND VPWR VPWR _12589_ sky130_fd_sc_hd__or2_1
XFILLER_0_187_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20671_ _12480_ _12517_ _12518_ VGND VGND VPWR VPWR _12520_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_86_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22410_ net80 net94 net89 VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__o21a_1
XFILLER_0_174_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23390_ _11650_ _02830_ net1020 VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_169_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22341_ _01643_ net91 VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25060_ _04370_ _04373_ _04368_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22272_ _01819_ _01823_ _01827_ _01831_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__o31a_2
X_24011_ _03056_ _03217_ _03363_ _03324_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__a22o_1
X_21223_ _12643_ _12618_ VGND VGND VPWR VPWR _13067_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold120 top0.pid_q.prev_error\[9\] VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 top0.svm0.tB\[1\] VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 top0.pid_q.prev_error\[6\] VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 top0.svm0.tC\[2\] VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 top0.svm0.tC\[5\] VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__dlygate4sd3_1
X_21154_ _12921_ _12931_ _12899_ VGND VGND VPWR VPWR _12999_ sky130_fd_sc_hd__o21ba_1
Xhold175 _00320_ VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 top0.periodTop\[13\] VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 top0.pid_q.prev_error\[2\] VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 net605 VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__clkbuf_4
Xfanout611 net612 VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__clkbuf_4
X_20105_ _11962_ _11963_ top0.cordic0.slte0.opA\[13\] VGND VGND VPWR VPWR _11964_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout622 net624 VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__buf_2
XFILLER_0_10_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25962_ top0.b_in_matmul\[0\] _05171_ _05165_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__mux2_1
X_21085_ _12927_ _12929_ _12930_ VGND VGND VPWR VPWR _12931_ sky130_fd_sc_hd__a21oi_2
Xfanout633 net634 VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout644 net645 VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__clkbuf_4
Xfanout655 net663 VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__clkbuf_4
X_24913_ _04222_ _04225_ _04263_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__o21a_1
Xfanout666 net669 VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__clkbuf_4
X_20036_ top0.cordic0.slte0.opA\[7\] _11899_ _11900_ _11898_ VGND VGND VPWR VPWR _00367_
+ sky130_fd_sc_hd__a22o_1
Xfanout677 net678 VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__clkbuf_4
X_25893_ top0.matmul0.alpha_pass\[11\] top0.matmul0.beta_pass\[11\] VGND VGND VPWR
+ VPWR _05110_ sky130_fd_sc_hd__xor2_4
Xfanout688 net689 VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__clkbuf_4
Xfanout699 net700 VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__clkbuf_4
X_24844_ _04096_ _04102_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24775_ _03995_ _04126_ _04127_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__a21oi_1
X_21987_ net135 _01338_ _01325_ _01548_ _01330_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__a221o_2
X_26514_ clknet_leaf_65_clk_sys _00137_ net659 VGND VGND VPWR VPWR top0.pid_q.out\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_166_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23726_ _03042_ _03052_ _03075_ _03082_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_194_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20938_ _12785_ _12683_ VGND VGND VPWR VPWR _12786_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26445_ clknet_leaf_87_clk_sys _00086_ net644 VGND VGND VPWR VPWR top0.kiq\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_193_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23657_ net569 net573 top0.matmul0.matmul_stage_inst.f\[2\] VGND VGND VPWR VPWR _03015_
+ sky130_fd_sc_hd__o21a_4
X_20869_ _12711_ _12712_ _12717_ VGND VGND VPWR VPWR _12718_ sky130_fd_sc_hd__a21o_1
XFILLER_0_187_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13410_ _05621_ _05622_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__nor2_1
X_22608_ _02160_ _02161_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14390_ _06501_ _06504_ _06508_ VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__a21boi_1
X_26376_ spi0.opcode\[6\] net963 net696 VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23588_ top0.matmul0.alpha_pass\[1\] _09255_ net560 VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__mux2_1
X_25327_ _04670_ _04671_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__xnor2_1
X_13341_ _05522_ _05525_ net50 net1015 VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__o211a_1
X_22539_ _02077_ _02079_ _02093_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16060_ _08063_ _08066_ _08064_ VGND VGND VPWR VPWR _08154_ sky130_fd_sc_hd__a21o_1
X_25258_ top0.matmul0.matmul_stage_inst.mult2\[11\] _04604_ _03146_ VGND VGND VPWR
+ VPWR _04605_ sky130_fd_sc_hd__mux2_1
X_13272_ top0.matmul0.beta_pass\[0\] _05435_ _05470_ _05464_ top0.c_out_calc\[0\]
+ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_122_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15011_ spi0.data_packed\[11\] top0.periodTop\[11\] _07125_ VGND VGND VPWR VPWR _07131_
+ sky130_fd_sc_hd__mux2_1
X_24209_ _03010_ _03549_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__nand2_1
X_25189_ _04536_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19750_ net201 net194 VGND VGND VPWR VPWR _11633_ sky130_fd_sc_hd__and2b_1
X_16962_ _09017_ _09005_ _09018_ VGND VGND VPWR VPWR _09019_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18701_ _10606_ _10678_ VGND VGND VPWR VPWR _10679_ sky130_fd_sc_hd__xnor2_2
X_15913_ net505 net483 _07972_ VGND VGND VPWR VPWR _08008_ sky130_fd_sc_hd__and3_1
X_16893_ net550 _08953_ _08954_ VGND VGND VPWR VPWR _08955_ sky130_fd_sc_hd__and3_1
X_19681_ _11552_ _11567_ VGND VGND VPWR VPWR _11568_ sky130_fd_sc_hd__xnor2_1
X_15844_ net454 net526 VGND VGND VPWR VPWR _07940_ sky130_fd_sc_hd__nand2_1
X_18632_ _10523_ _10528_ _10609_ _10255_ VGND VGND VPWR VPWR _10610_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_188_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18563_ _10465_ _10467_ _10466_ VGND VGND VPWR VPWR _10542_ sky130_fd_sc_hd__o21a_1
X_15775_ _07727_ _07728_ _07726_ VGND VGND VPWR VPWR _07872_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14726_ _06832_ _05640_ _06323_ _06928_ net25 VGND VGND VPWR VPWR _06929_ sky130_fd_sc_hd__a32o_1
X_17514_ net391 _09395_ _09500_ net395 VGND VGND VPWR VPWR _09501_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18494_ net334 net369 VGND VGND VPWR VPWR _10474_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17445_ net395 net392 VGND VGND VPWR VPWR _09432_ sky130_fd_sc_hd__or2_1
X_14657_ _06819_ _06858_ VGND VGND VPWR VPWR _06861_ sky130_fd_sc_hd__or2_1
XFILLER_0_200_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13608_ _05818_ _05819_ _05820_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17376_ _09362_ VGND VGND VPWR VPWR _09363_ sky130_fd_sc_hd__buf_2
X_14588_ _06742_ _06744_ VGND VGND VPWR VPWR _06794_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16327_ net447 net516 VGND VGND VPWR VPWR _08417_ sky130_fd_sc_hd__nand2_1
X_19115_ top0.pid_d.out\[14\] top0.pid_d.curr_int\[14\] _11082_ _11086_ net432 VGND
+ VGND VPWR VPWR _11087_ sky130_fd_sc_hd__o311a_1
X_13539_ _05708_ _05693_ _05695_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19046_ _10494_ _11018_ VGND VGND VPWR VPWR _11019_ sky130_fd_sc_hd__xnor2_1
X_16258_ _08255_ _08257_ _08256_ VGND VGND VPWR VPWR _08349_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15209_ _07305_ _07306_ _07307_ VGND VGND VPWR VPWR _07308_ sky130_fd_sc_hd__o21a_1
X_16189_ _08275_ _08280_ VGND VGND VPWR VPWR _08281_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19948_ top0.cordic0.slte0.opA\[1\] _11785_ VGND VGND VPWR VPWR _11819_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19879_ _11526_ _11754_ net175 VGND VGND VPWR VPWR _11755_ sky130_fd_sc_hd__o21ai_1
X_21910_ _01464_ _01463_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__xor2_2
X_22890_ top0.svm0.calc_ready _02297_ _02408_ net708 _02309_ VGND VGND VPWR VPWR _00440_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21841_ _01398_ _01399_ _01396_ _01401_ _01402_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_136_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24560_ _03905_ _03914_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_136_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21772_ _01324_ _01326_ _01333_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23511_ net794 top0.matmul0.cos\[10\] _02915_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__mux2_1
X_20723_ net306 _12549_ VGND VGND VPWR VPWR _12572_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24491_ _03663_ _03676_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26230_ spi0.data_packed\[13\] net19 net694 VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23442_ _02657_ net217 _11776_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__mux2_2
XFILLER_0_163_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20654_ _12469_ _12502_ VGND VGND VPWR VPWR _12503_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26161_ _05301_ top0.cordic0.slte0.opB\[7\] _12006_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__mux2_1
X_20585_ _12430_ _12431_ _12432_ VGND VGND VPWR VPWR _12434_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23373_ _02814_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25112_ _04455_ _04460_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22324_ _01806_ _01875_ _01882_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__o21ai_2
X_26092_ top0.pid_d.out\[15\] _12031_ _05013_ spi0.data_packed\[79\] VGND VGND VPWR
+ VPWR _05271_ sky130_fd_sc_hd__a22o_1
X_25043_ _04305_ _04312_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22255_ _01765_ _01770_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21206_ _13045_ _13048_ VGND VGND VPWR VPWR _13050_ sky130_fd_sc_hd__nor2_1
X_22186_ _01711_ _01718_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21137_ _11727_ _12981_ _12893_ VGND VGND VPWR VPWR _12982_ sky130_fd_sc_hd__a21oi_4
X_26994_ clknet_leaf_23_clk_sys _00611_ net625 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout430 top0.matmul0.beta_pass\[10\] VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__buf_2
Xfanout441 top0.pid_d.state\[1\] VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkbuf_4
Xfanout452 net454 VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__clkbuf_4
Xfanout463 top0.pid_q.mult0.b\[8\] VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__clkbuf_2
X_25945_ _05145_ _05146_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__nor2_1
X_21068_ _12910_ _12913_ VGND VGND VPWR VPWR _12914_ sky130_fd_sc_hd__xnor2_2
Xfanout474 top0.pid_q.mult0.b\[5\] VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__buf_2
Xfanout485 net486 VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__clkbuf_2
Xfanout496 top0.pid_q.mult0.b\[0\] VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__buf_4
X_20019_ top0.cordic0.slte0.opA\[5\] _11866_ _11884_ VGND VGND VPWR VPWR _11885_ sky130_fd_sc_hd__a21o_1
X_13890_ _06086_ _06087_ _06100_ _06101_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__or4_4
X_25876_ _05082_ _05083_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__nor2_1
XFILLER_0_198_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24827_ _04172_ _04178_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15560_ _07637_ _07658_ VGND VGND VPWR VPWR _07659_ sky130_fd_sc_hd__xor2_1
X_24758_ _04107_ _04110_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14511_ _06640_ _06212_ _06715_ net25 VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__o22a_1
X_23709_ net572 top0.matmul0.matmul_stage_inst.d\[2\] top0.matmul0.matmul_stage_inst.c\[2\]
+ net556 VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__a22o_2
XFILLER_0_166_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15491_ _07193_ _07191_ VGND VGND VPWR VPWR _07590_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24689_ _03572_ _04042_ _04040_ _03549_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17230_ _08738_ _09192_ _09235_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14442_ _06648_ _06649_ VGND VGND VPWR VPWR _06650_ sky130_fd_sc_hd__or2_2
X_26428_ clknet_leaf_77_clk_sys _00069_ net631 VGND VGND VPWR VPWR top0.kid\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout70 net71 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_182_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout81 top0.cordic0.vec\[1\]\[17\] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_2
Xfanout92 net93 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
X_17161_ net543 _08157_ _09174_ net553 _08955_ VGND VGND VPWR VPWR _09175_ sky130_fd_sc_hd__a221o_1
X_14373_ _06516_ _06527_ VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26359_ _05411_ VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16112_ _08201_ _08204_ VGND VGND VPWR VPWR _08205_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13324_ top0.matmul0.beta_pass\[8\] _05434_ _05469_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17092_ net860 _09115_ _09122_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16043_ _08092_ _08136_ VGND VGND VPWR VPWR _08137_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_51_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13255_ net76 _05466_ _05467_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19802_ net260 _11664_ _11681_ _11682_ VGND VGND VPWR VPWR _11683_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_202_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17994_ net1018 _09979_ VGND VGND VPWR VPWR _09980_ sky130_fd_sc_hd__and2_1
X_19733_ _11581_ _11582_ _11600_ VGND VGND VPWR VPWR _11617_ sky130_fd_sc_hd__or3_1
X_16945_ top0.pid_q.curr_error\[8\] VGND VGND VPWR VPWR _09003_ sky130_fd_sc_hd__inv_2
X_19664_ _11543_ _11531_ _11533_ _11534_ net297 VGND VGND VPWR VPWR _11551_ sky130_fd_sc_hd__a41o_1
X_16876_ _08936_ _08925_ _08938_ VGND VGND VPWR VPWR _08939_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_126_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18615_ _10593_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__clkbuf_1
X_15827_ _07819_ _07824_ _07922_ VGND VGND VPWR VPWR _07923_ sky130_fd_sc_hd__a21o_1
X_19595_ _11455_ _11463_ _11483_ VGND VGND VPWR VPWR _11484_ sky130_fd_sc_hd__a21o_4
XFILLER_0_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18546_ net387 net314 VGND VGND VPWR VPWR _10525_ sky130_fd_sc_hd__nand2_1
X_15758_ _07754_ _07755_ _07854_ VGND VGND VPWR VPWR _07855_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_142_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14709_ _06873_ _06911_ _06877_ VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__o21a_1
X_18477_ net369 _10456_ net341 VGND VGND VPWR VPWR _10457_ sky130_fd_sc_hd__or3b_1
X_15689_ _07671_ _07675_ VGND VGND VPWR VPWR _07787_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17428_ net407 net343 VGND VGND VPWR VPWR _09415_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17359_ net412 net347 VGND VGND VPWR VPWR _09346_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20370_ _12210_ _12211_ _12217_ VGND VGND VPWR VPWR _12219_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_15_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19029_ net360 net316 _10944_ VGND VGND VPWR VPWR _11002_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22040_ _01262_ _01601_ _01151_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23991_ _03346_ _03348_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_177_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25730_ net808 _04964_ _04913_ _04984_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__a22o_1
X_22942_ _02440_ _02454_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25661_ net735 _04904_ _04935_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__a21bo_1
X_22873_ top0.svm0.tB\[7\] _02390_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__and2_1
XFILLER_0_183_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24612_ _03890_ _03891_ _03892_ _03893_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__a211o_1
X_21824_ _01377_ _01384_ _01385_ _01217_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25592_ _04885_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__buf_2
XFILLER_0_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24543_ _03882_ _03897_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__xor2_2
X_21755_ _01289_ _01316_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__xnor2_1
X_20706_ net296 _12553_ _12554_ VGND VGND VPWR VPWR _12555_ sky130_fd_sc_hd__a21oi_1
X_27262_ clknet_3_4__leaf_clk_mosi _00876_ VGND VGND VPWR VPWR spi0.data_packed\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_24474_ _03549_ _03829_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__nand2_2
XFILLER_0_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21686_ net96 net90 VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__nand2_2
X_26213_ _05338_ VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23425_ _11650_ _02862_ _11954_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__a21o_1
X_27193_ clknet_leaf_56_clk_sys _00807_ net668 VGND VGND VPWR VPWR top0.currT_r\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_11_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20637_ _12471_ _12477_ _12484_ _12485_ VGND VGND VPWR VPWR _12486_ sky130_fd_sc_hd__a211o_1
XFILLER_0_18_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26144_ _05288_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__clkbuf_1
X_23356_ _02796_ _02798_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20568_ _12411_ _12414_ VGND VGND VPWR VPWR _12417_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22307_ _01861_ _01866_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__xnor2_4
X_26075_ _05258_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__clkbuf_1
X_23287_ _02725_ _02734_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__xnor2_1
X_20499_ net282 net295 VGND VGND VPWR VPWR _12348_ sky130_fd_sc_hd__and2b_1
X_25026_ _04363_ _04375_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22238_ _01213_ net106 net100 net87 _01762_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__a221o_1
X_22169_ _01160_ _01730_ _01165_ _01247_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_79_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14991_ _07120_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__clkbuf_1
X_26977_ clknet_leaf_25_clk_sys _00594_ net627 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[9\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout260 net261 VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__buf_1
Xfanout271 net272 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_4
Xfanout282 net284 VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__clkbuf_4
X_13942_ _06143_ _06154_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__xnor2_4
X_16730_ _08718_ _08813_ VGND VGND VPWR VPWR _08814_ sky130_fd_sc_hd__nand2_1
X_25928_ net936 _05028_ _05031_ _05142_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__a22o_1
Xfanout293 top0.cordic0.vec\[0\]\[3\] VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16661_ _08312_ _08693_ VGND VGND VPWR VPWR _08746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13873_ _05763_ _05768_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__nor2_1
X_25859_ net11 _05077_ _05079_ _02282_ _12014_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_72_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18400_ _10275_ _10284_ _10283_ VGND VGND VPWR VPWR _10381_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15612_ _07702_ _07709_ _07710_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__o21a_1
X_16592_ _08600_ _08601_ _08678_ VGND VGND VPWR VPWR _08679_ sky130_fd_sc_hd__mux2_1
X_19380_ top0.pid_d.prev_error\[13\] _11284_ _11287_ net910 VGND VGND VPWR VPWR _00323_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_201_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18331_ _10311_ _10210_ _10312_ VGND VGND VPWR VPWR _10313_ sky130_fd_sc_hd__a21boi_1
X_15543_ _07638_ _07641_ VGND VGND VPWR VPWR _07642_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18262_ top0.pid_d.out\[4\] _09339_ _10244_ _10067_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15474_ net540 net538 net454 net457 VGND VGND VPWR VPWR _07573_ sky130_fd_sc_hd__and4_1
XFILLER_0_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14425_ _06025_ net1015 _06320_ _06587_ _06589_ VGND VGND VPWR VPWR _06633_ sky130_fd_sc_hd__a32o_1
XFILLER_0_182_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17213_ _08609_ _09176_ VGND VGND VPWR VPWR _09221_ sky130_fd_sc_hd__nor2_1
X_18193_ net1023 net395 VGND VGND VPWR VPWR _10176_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17144_ _09157_ _09158_ VGND VGND VPWR VPWR _09160_ sky130_fd_sc_hd__or2_1
X_14356_ _06561_ _06564_ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_123_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13307_ _05475_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__buf_2
XFILLER_0_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17075_ _09112_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14287_ net39 _05611_ _05612_ VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16026_ _08108_ _08119_ VGND VGND VPWR VPWR _08120_ sky130_fd_sc_hd__xor2_1
X_13238_ net441 _05449_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17977_ _09874_ _09877_ VGND VGND VPWR VPWR _09963_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19716_ _11581_ _11582_ _11512_ VGND VGND VPWR VPWR _11601_ sky130_fd_sc_hd__o21a_1
X_16928_ _08984_ _08986_ VGND VGND VPWR VPWR _08987_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19647_ net98 net94 net88 net83 net199 net193 VGND VGND VPWR VPWR _11535_ sky130_fd_sc_hd__mux4_2
XFILLER_0_189_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16859_ top0.pid_q.prev_error\[2\] VGND VGND VPWR VPWR _08923_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19578_ top0.cordic0.slte0.opA\[11\] top0.cordic0.slte0.opB\[11\] VGND VGND VPWR
+ VPWR _11467_ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18529_ net434 _10431_ _10432_ _10508_ net436 VGND VGND VPWR VPWR _10509_ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21540_ _01080_ VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__buf_4
XFILLER_0_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21471_ _00978_ _01034_ _01035_ _00975_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23210_ _01320_ _02661_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20422_ _12268_ _12270_ VGND VGND VPWR VPWR _12271_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24190_ _03495_ _03497_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_160_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23141_ _02440_ _02628_ _02596_ VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__o21ai_1
X_20353_ net253 net267 VGND VGND VPWR VPWR _12202_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23072_ _02564_ _02569_ _02572_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__o21a_1
X_20284_ _12127_ _12132_ VGND VGND VPWR VPWR _12133_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22023_ _01356_ _01487_ _01584_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__and3_1
X_26900_ clknet_leaf_108_clk_sys _00517_ net585 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26831_ clknet_leaf_46_clk_sys _00448_ net680 VGND VGND VPWR VPWR top0.svm0.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold13 top0.kpq\[11\] VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 top0.cordic0.sin\[8\] VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 top0.matmul0.matmul_stage_inst.c\[6\] VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 top0.matmul0.matmul_stage_inst.d\[12\] VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26762_ clknet_leaf_93_clk_sys _00379_ net599 VGND VGND VPWR VPWR top0.cordic0.domain\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold57 top0.kpq\[1\] VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__dlygate4sd3_1
X_23974_ _03242_ _03331_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__xnor2_2
Xhold68 top0.matmul0.matmul_stage_inst.a\[1\] VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 top0.matmul0.matmul_stage_inst.c\[7\] VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25713_ _04883_ _04920_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__or2_1
XFILLER_0_202_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22925_ _02440_ _02437_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__nor2_1
X_26693_ clknet_leaf_64_clk_sys _00310_ net658 VGND VGND VPWR VPWR top0.pid_d.prev_error\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_76_clk_sys clknet_3_4__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_76_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_25644_ _04884_ top0.matmul0.sin\[4\] _04914_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__and3_1
XFILLER_0_196_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22856_ top0.svm0.tA\[14\] _02375_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21807_ _01294_ _01269_ net162 VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25575_ top0.matmul0.a\[10\] top0.matmul0.matmul_stage_inst.e\[10\] _04867_ VGND
+ VGND VPWR VPWR _04875_ sky130_fd_sc_hd__mux2_1
X_22787_ top0.svm0.state\[1\] top0.start_svm _02308_ _02309_ VGND VGND VPWR VPWR _00436_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_195_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24526_ _03869_ _03804_ _03809_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__mux2_1
X_21738_ net154 net148 VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27245_ clknet_3_5__leaf_clk_mosi _00859_ VGND VGND VPWR VPWR spi0.data_packed\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_24457_ _03798_ _03812_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21669_ net105 net90 _01230_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_49_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14210_ _05500_ _05531_ _05532_ VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__or3_2
XFILLER_0_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_193_Right_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23408_ _11514_ _02846_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__nand2_1
X_27176_ clknet_leaf_32_clk_sys _00790_ net619 VGND VGND VPWR VPWR top0.periodTop_r\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_15190_ net538 net457 VGND VGND VPWR VPWR _07289_ sky130_fd_sc_hd__nand2_2
X_24388_ _03740_ _03744_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__xor2_2
X_14141_ _06351_ _06193_ _06135_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__o21ai_1
X_26127_ spi0.data_packed\[22\] _05281_ _05282_ net960 VGND VGND VPWR VPWR _00803_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23339_ _02781_ _02782_ _02756_ _02762_ _02763_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_160_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14072_ _06282_ _06283_ VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__xnor2_2
X_26058_ top0.a_in_matmul\[6\] _05245_ _05230_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25009_ _04355_ _04358_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__xnor2_2
X_17900_ _09754_ _09755_ _09775_ VGND VGND VPWR VPWR _09887_ sky130_fd_sc_hd__a21o_1
X_18880_ net389 _10494_ _10810_ VGND VGND VPWR VPWR _10855_ sky130_fd_sc_hd__or3b_2
X_17831_ _09702_ _09705_ _09713_ VGND VGND VPWR VPWR _09818_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_58_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17762_ _09406_ _09368_ _09748_ VGND VGND VPWR VPWR _09749_ sky130_fd_sc_hd__o21a_1
X_14974_ _07109_ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__clkbuf_1
X_19501_ _11384_ _11391_ _11392_ VGND VGND VPWR VPWR _11393_ sky130_fd_sc_hd__a21o_1
X_16713_ _00011_ _07700_ _08791_ _08797_ _07800_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__a32o_1
X_13925_ _06130_ _06137_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__xnor2_2
X_17693_ _09621_ _09678_ _09679_ VGND VGND VPWR VPWR _09680_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_57_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19432_ _11330_ _11331_ VGND VGND VPWR VPWR _11332_ sky130_fd_sc_hd__xnor2_1
X_16644_ _08662_ _08666_ _08729_ VGND VGND VPWR VPWR _08730_ sky130_fd_sc_hd__o21ai_2
X_13856_ _06019_ _06068_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_190_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19363_ _11284_ VGND VGND VPWR VPWR _11285_ sky130_fd_sc_hd__clkbuf_4
X_16575_ _08582_ _08585_ _08661_ VGND VGND VPWR VPWR _08662_ sky130_fd_sc_hd__o21ai_2
X_13787_ net58 _05496_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18314_ _10293_ _10295_ VGND VGND VPWR VPWR _10296_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15526_ net472 net518 VGND VGND VPWR VPWR _07625_ sky130_fd_sc_hd__nand2_1
X_19294_ _11234_ _11235_ VGND VGND VPWR VPWR _11236_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_67_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18245_ net307 _09967_ VGND VGND VPWR VPWR _10228_ sky130_fd_sc_hd__nand2_2
X_15457_ _07267_ _07268_ _07555_ VGND VGND VPWR VPWR _07556_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_155_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14408_ net41 _05619_ VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__nand2_2
XFILLER_0_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_160_Right_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18176_ top0.pid_d.curr_int\[3\] _10069_ _10158_ VGND VGND VPWR VPWR _10159_ sky130_fd_sc_hd__o21a_1
X_15388_ net541 net482 _07475_ VGND VGND VPWR VPWR _07487_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_167_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14339_ _06471_ VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17127_ net553 _09143_ _09144_ net548 _08897_ VGND VGND VPWR VPWR _09145_ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17058_ net929 _09100_ _09102_ _08935_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16009_ _08101_ _08102_ VGND VGND VPWR VPWR _08103_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20971_ _12773_ _12817_ VGND VGND VPWR VPWR _12818_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22710_ _02210_ _02224_ _02183_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__or3b_1
X_23690_ _03047_ _02982_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__nor2_2
XFILLER_0_67_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22641_ _01643_ _02193_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_193_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25360_ _04612_ _04704_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__or2_1
X_22572_ _02094_ _02126_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24311_ _03666_ _03667_ _03087_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_111_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21523_ _01073_ _01077_ _01084_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__a21bo_1
X_25291_ _04635_ _04636_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__or2b_2
XFILLER_0_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27030_ clknet_leaf_27_clk_sys _00647_ net621 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_24242_ _03558_ _03570_ _03582_ _03594_ _03599_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21454_ _01018_ _01012_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20405_ _12253_ VGND VGND VPWR VPWR _12254_ sky130_fd_sc_hd__inv_2
X_24173_ _03411_ _03527_ _03410_ _03414_ _03413_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__a32o_1
X_21385_ _00951_ _00952_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__xor2_1
X_23124_ top0.svm0.delta\[7\] top0.svm0.delta\[8\] _02612_ _02595_ VGND VGND VPWR
+ VPWR _02617_ sky130_fd_sc_hd__o31a_1
X_20336_ _12182_ _12183_ _12181_ VGND VGND VPWR VPWR _12185_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23055_ _02553_ _02554_ _02555_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__a21bo_1
X_20267_ _12083_ _12070_ _12071_ VGND VGND VPWR VPWR _12116_ sky130_fd_sc_hd__and3_1
X_22006_ _01563_ _01567_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__xnor2_1
X_20198_ net299 net296 VGND VGND VPWR VPWR _12047_ sky130_fd_sc_hd__nand2_2
X_26814_ clknet_leaf_51_clk_sys _00431_ net670 VGND VGND VPWR VPWR top0.pid_q.prev_int\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23957_ _03314_ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__clkbuf_4
X_26745_ clknet_leaf_96_clk_sys _00362_ net588 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13710_ _05909_ _05921_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__or2_1
X_22908_ net169 _02409_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__nor2_1
X_14690_ _06839_ _06844_ _06837_ VGND VGND VPWR VPWR _06894_ sky130_fd_sc_hd__o21ba_1
X_26676_ clknet_leaf_81_clk_sys _00293_ net636 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[15\]
+ sky130_fd_sc_hd__dfrtp_2
X_23888_ _03243_ _03244_ _03245_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__o21a_1
XFILLER_0_196_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13641_ _05828_ _05809_ _05851_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__nand3_1
X_22839_ top0.svm0.counter\[4\] _02322_ _02330_ _02333_ _02358_ VGND VGND VPWR VPWR
+ _02359_ sky130_fd_sc_hd__a2111o_1
X_25627_ _04905_ _04906_ net69 VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16360_ net469 _08141_ _08048_ _08449_ VGND VGND VPWR VPWR _08450_ sky130_fd_sc_hd__nand4_1
XFILLER_0_52_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13572_ _05770_ _05784_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__xnor2_2
X_25558_ top0.matmul0.a\[2\] top0.matmul0.matmul_stage_inst.e\[2\] _04856_ VGND VGND
+ VPWR VPWR _04866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15311_ net1026 net491 VGND VGND VPWR VPWR _07410_ sky130_fd_sc_hd__nand2_1
X_24509_ _03207_ _03208_ _03103_ _03104_ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__o22a_2
XFILLER_0_137_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16291_ _08296_ _08300_ _08298_ VGND VGND VPWR VPWR _08382_ sky130_fd_sc_hd__a21o_1
X_25489_ _04830_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18030_ _09910_ _09911_ _10014_ VGND VGND VPWR VPWR _10015_ sky130_fd_sc_hd__a21bo_1
X_15242_ _07339_ _07340_ _07233_ VGND VGND VPWR VPWR _07341_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27228_ clknet_3_4__leaf_clk_mosi _00842_ VGND VGND VPWR VPWR spi0.data_packed\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15173_ _07198_ _07199_ _07197_ VGND VGND VPWR VPWR _07272_ sky130_fd_sc_hd__o21ai_1
X_27159_ clknet_leaf_6_clk_sys _00773_ net594 VGND VGND VPWR VPWR top0.a_in_matmul\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14124_ net22 _06046_ _05496_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__and3_1
X_19981_ _11812_ _11845_ _11846_ _11848_ VGND VGND VPWR VPWR _11849_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14055_ _06135_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__buf_4
XFILLER_0_162_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18932_ _10828_ _10829_ VGND VGND VPWR VPWR _10907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18863_ top0.pid_d.out\[11\] _07138_ _10838_ net432 VGND VGND VPWR VPWR _10839_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17814_ _09671_ _09799_ _09800_ VGND VGND VPWR VPWR _09801_ sky130_fd_sc_hd__a21oi_2
X_18794_ _10458_ _10720_ net341 VGND VGND VPWR VPWR _10770_ sky130_fd_sc_hd__o21a_1
X_17745_ _09729_ _09731_ _09503_ VGND VGND VPWR VPWR _09732_ sky130_fd_sc_hd__mux2_1
X_14957_ _07100_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13908_ _05772_ _05783_ _05770_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__a21o_1
X_17676_ net426 _09609_ _09612_ VGND VGND VPWR VPWR _09663_ sky130_fd_sc_hd__or3_1
X_14888_ _07041_ VGND VGND VPWR VPWR _07064_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19415_ _11315_ _11308_ _11310_ _11316_ VGND VGND VPWR VPWR _11317_ sky130_fd_sc_hd__a31o_1
XFILLER_0_202_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16627_ _08709_ _08712_ VGND VGND VPWR VPWR _08713_ sky130_fd_sc_hd__nor2_1
X_13839_ _06029_ _06026_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__xor2_1
XFILLER_0_175_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19346_ _05439_ _00003_ _11276_ VGND VGND VPWR VPWR _11279_ sky130_fd_sc_hd__and3_1
X_16558_ _08560_ _08565_ _08644_ VGND VGND VPWR VPWR _08645_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15509_ _07298_ _07599_ VGND VGND VPWR VPWR _07608_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19277_ top0.matmul0.alpha_pass\[10\] _11210_ VGND VGND VPWR VPWR _11221_ sky130_fd_sc_hd__or2_1
X_16489_ _08571_ _08576_ VGND VGND VPWR VPWR _08577_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18228_ net410 net313 VGND VGND VPWR VPWR _10211_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_24_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_24_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_5_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18159_ _10141_ _10142_ VGND VGND VPWR VPWR _10143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold302 top0.cordic0.cos\[4\] VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21170_ _12952_ _12960_ _13010_ VGND VGND VPWR VPWR _13014_ sky130_fd_sc_hd__and3b_1
XFILLER_0_68_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20121_ top0.cordic0.slte0.opA\[14\] _11970_ _11977_ VGND VGND VPWR VPWR _11978_
+ sky130_fd_sc_hd__o21a_2
XFILLER_0_1_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20052_ net183 _11513_ _11657_ _11904_ VGND VGND VPWR VPWR _11915_ sky130_fd_sc_hd__a22o_1
X_24860_ _04195_ _04211_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_139_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23811_ _03139_ _03141_ _03167_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__a21oi_2
X_24791_ _04035_ _04142_ _04143_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26530_ clknet_leaf_61_clk_sys _00153_ net651 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_23742_ _03097_ _03099_ _03082_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__mux2_2
X_20954_ _12752_ _12801_ VGND VGND VPWR VPWR _12802_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26461_ clknet_leaf_91_clk_sys net702 net640 VGND VGND VPWR VPWR spi0.cs_sync\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_191_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23673_ _03027_ _03028_ _03029_ _03030_ VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__o22a_1
XFILLER_0_193_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20885_ _12179_ _12733_ _12242_ VGND VGND VPWR VPWR _12734_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25412_ _04701_ _04707_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__nand2_1
X_22624_ net211 _02176_ _02175_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__a21bo_1
X_26392_ clknet_leaf_37_clk_sys _00033_ net679 VGND VGND VPWR VPWR top0.svm0.tC\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25343_ _04633_ _04687_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22555_ _01769_ _01798_ net115 VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__mux2_1
X_21506_ _01064_ _01067_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__nand2_1
X_25274_ net1017 _03936_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22486_ _02041_ _02042_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__and2b_1
XFILLER_0_146_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27013_ clknet_leaf_24_clk_sys _00630_ net626 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_24225_ _03576_ _03577_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21437_ _00967_ _00982_ _00945_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24156_ _03490_ _03498_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__xnor2_1
X_21368_ _13001_ _13174_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23107_ _02440_ _02604_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20319_ _12163_ _12167_ VGND VGND VPWR VPWR _12168_ sky130_fd_sc_hd__xnor2_1
X_24087_ _03333_ _03443_ _03444_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__or3_2
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21299_ _13110_ _13141_ VGND VGND VPWR VPWR _13142_ sky130_fd_sc_hd__xor2_2
XFILLER_0_102_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23038_ net57 _02538_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__or2_1
X_15860_ _07849_ _07851_ _07955_ VGND VGND VPWR VPWR _07956_ sky130_fd_sc_hd__a21oi_2
X_14811_ _06974_ _06977_ _07009_ VGND VGND VPWR VPWR _07011_ sky130_fd_sc_hd__a21o_1
X_15791_ net481 _07886_ _07887_ _07765_ VGND VGND VPWR VPWR _07888_ sky130_fd_sc_hd__o2bb2a_1
X_24989_ _03234_ _03007_ _03765_ _04039_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17530_ _09391_ _09368_ _09405_ _09446_ VGND VGND VPWR VPWR _09517_ sky130_fd_sc_hd__or4b_1
XFILLER_0_54_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14742_ _06910_ _06944_ VGND VGND VPWR VPWR _06945_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_118_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26728_ clknet_leaf_104_clk_sys _00345_ net576 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_93_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14673_ net39 _06268_ VGND VGND VPWR VPWR _06877_ sky130_fd_sc_hd__nand2_1
X_17461_ _09368_ _09447_ VGND VGND VPWR VPWR _09448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26659_ clknet_leaf_77_clk_sys _00276_ net635 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_168_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19200_ top0.matmul0.alpha_pass\[3\] _11141_ VGND VGND VPWR VPWR _11151_ sky130_fd_sc_hd__nand2_1
X_16412_ net1028 net444 VGND VGND VPWR VPWR _08501_ sky130_fd_sc_hd__nand2b_2
X_13624_ _05819_ _05836_ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__xnor2_1
X_17392_ _09378_ VGND VGND VPWR VPWR _09379_ sky130_fd_sc_hd__buf_2
XFILLER_0_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19131_ top0.kid\[0\] _11098_ _11100_ top0.kpd\[0\] VGND VGND VPWR VPWR _11101_ sky130_fd_sc_hd__a22o_1
X_13555_ _05764_ _05767_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__xnor2_2
X_16343_ _08431_ _08432_ VGND VGND VPWR VPWR _08433_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16274_ net467 net500 VGND VGND VPWR VPWR _08365_ sky130_fd_sc_hd__nand2_2
XFILLER_0_125_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19062_ _11033_ _11034_ VGND VGND VPWR VPWR _11035_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13486_ _05697_ _05698_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__xor2_1
XFILLER_0_180_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18013_ _09992_ _09997_ VGND VGND VPWR VPWR _09998_ sky130_fd_sc_hd__nor2_1
X_15225_ _07320_ _07323_ VGND VGND VPWR VPWR _07324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15156_ _07253_ _07254_ VGND VGND VPWR VPWR _07255_ sky130_fd_sc_hd__nand2_2
XFILLER_0_196_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14107_ _06317_ _06318_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19964_ _11612_ _11574_ VGND VGND VPWR VPWR _11833_ sky130_fd_sc_hd__or2_1
X_15087_ _07176_ _07185_ VGND VGND VPWR VPWR _07186_ sky130_fd_sc_hd__nand2_1
X_14038_ _06242_ _06250_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__nor2_1
X_18915_ _10875_ _10889_ VGND VGND VPWR VPWR _10890_ sky130_fd_sc_hd__xnor2_2
X_19895_ _11759_ _11768_ _11769_ VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18846_ _10738_ _10739_ _10733_ VGND VGND VPWR VPWR _10822_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18777_ _10684_ _10753_ VGND VGND VPWR VPWR _10754_ sky130_fd_sc_hd__xor2_2
X_15989_ top0.pid_q.curr_int\[4\] _08078_ _08082_ VGND VGND VPWR VPWR _08083_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17728_ _09702_ _09705_ _09713_ VGND VGND VPWR VPWR _09715_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_171_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17659_ _09644_ _09645_ VGND VGND VPWR VPWR _09646_ sky130_fd_sc_hd__xor2_1
XFILLER_0_175_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20670_ _12517_ _12518_ _12480_ VGND VGND VPWR VPWR _12519_ sky130_fd_sc_hd__a21bo_1
X_19329_ _11266_ _11267_ VGND VGND VPWR VPWR _11268_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_174_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22340_ _01839_ _01856_ _01857_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22271_ _01829_ _01828_ _01830_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24010_ _03366_ _03367_ _03248_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__a21oi_1
Xhold110 top0.svm0.tC\[7\] VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__dlygate4sd3_1
X_21222_ _12620_ VGND VGND VPWR VPWR _13066_ sky130_fd_sc_hd__inv_2
Xhold121 top0.svm0.tB\[5\] VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold132 top0.periodTop\[11\] VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold143 top0.kpq\[0\] VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 top0.matmul0.matmul_stage_inst.c\[10\] VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 top0.pid_q.curr_error\[14\] VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__dlygate4sd3_1
X_21153_ _12967_ _12997_ VGND VGND VPWR VPWR _12998_ sky130_fd_sc_hd__xnor2_2
Xhold176 top0.pid_d.prev_error\[8\] VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold187 top0.matmul0.matmul_stage_inst.b\[1\] VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 net602 VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold198 top0.pid_q.prev_error\[11\] VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 net615 VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__clkbuf_4
X_20104_ _11649_ _11961_ _11954_ VGND VGND VPWR VPWR _11963_ sky130_fd_sc_hd__a21o_1
Xfanout623 net624 VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__clkbuf_4
X_25961_ top0.matmul0.beta_pass\[0\] _05169_ _05170_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__a21o_1
X_21084_ _11727_ net225 _11788_ _12851_ VGND VGND VPWR VPWR _12930_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout634 net635 VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__clkbuf_4
Xfanout645 net654 VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout656 net658 VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__clkbuf_4
X_24912_ _04222_ _04225_ _04258_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__a21o_1
Xfanout667 net669 VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__clkbuf_4
X_20035_ top0.cordic0.slte0.opA\[7\] _11785_ VGND VGND VPWR VPWR _11900_ sky130_fd_sc_hd__nor2_1
X_25892_ _05109_ _12014_ net840 _05029_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__a2bb2o_1
Xfanout678 net679 VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__clkbuf_4
Xfanout689 net693 VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__clkbuf_2
X_24843_ _04185_ _04194_ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24774_ _04028_ _04029_ _03991_ _03992_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__o211a_1
XFILLER_0_197_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21986_ net147 _01311_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__nand2_1
X_23725_ _03042_ _03044_ _03075_ _03082_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__a22o_1
X_26513_ clknet_leaf_65_clk_sys _00136_ net657 VGND VGND VPWR VPWR top0.pid_q.out\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_200_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20937_ _12700_ VGND VGND VPWR VPWR _12785_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23656_ _03008_ _03009_ _03013_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_3_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26444_ clknet_leaf_87_clk_sys _00085_ net644 VGND VGND VPWR VPWR top0.kiq\[1\] sky130_fd_sc_hd__dfrtp_1
X_20868_ _12095_ _12716_ VGND VGND VPWR VPWR _12717_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22607_ _02159_ _02154_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__or2b_1
X_26375_ _05419_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__clkbuf_1
X_23587_ _02960_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20799_ _12546_ _12579_ _12606_ _12647_ VGND VGND VPWR VPWR _12648_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25326_ _03900_ _04182_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__nor2_1
X_13340_ _05549_ _05550_ _05552_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22538_ _02007_ _02084_ _02085_ _02082_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25257_ _04539_ _04603_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__xnor2_1
X_13271_ _05483_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__clkbuf_4
X_22469_ net85 _02025_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15010_ _07130_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__clkbuf_1
X_24208_ _03563_ _03565_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__and2_1
X_25188_ top0.matmul0.matmul_stage_inst.mult2\[10\] _04535_ _03146_ VGND VGND VPWR
+ VPWR _04536_ sky130_fd_sc_hd__mux2_1
X_24139_ _03496_ _03161_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__nor2_2
X_16961_ _09017_ _09005_ top0.pid_q.prev_error\[9\] VGND VGND VPWR VPWR _09018_ sky130_fd_sc_hd__o21ba_1
X_18700_ _10676_ _10677_ VGND VGND VPWR VPWR _10678_ sky130_fd_sc_hd__or2_1
X_15912_ net502 _08005_ _08006_ net499 VGND VGND VPWR VPWR _08007_ sky130_fd_sc_hd__a22o_1
X_19680_ _11565_ _11566_ VGND VGND VPWR VPWR _11567_ sky130_fd_sc_hd__xnor2_2
X_16892_ _08951_ _08952_ VGND VGND VPWR VPWR _08954_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18631_ net382 _09518_ _09689_ _10074_ VGND VGND VPWR VPWR _10609_ sky130_fd_sc_hd__a22o_1
X_15843_ net451 net529 VGND VGND VPWR VPWR _07939_ sky130_fd_sc_hd__nand2_1
X_18562_ _10537_ _10540_ VGND VGND VPWR VPWR _10541_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_188_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15774_ _07732_ _07736_ _07870_ VGND VGND VPWR VPWR _07871_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17513_ _09498_ _09499_ VGND VGND VPWR VPWR _09500_ sky130_fd_sc_hd__nand2_1
X_14725_ _06832_ _06927_ net20 VGND VGND VPWR VPWR _06928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18493_ net331 net373 VGND VGND VPWR VPWR _10473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17444_ net407 net357 VGND VGND VPWR VPWR _09431_ sky130_fd_sc_hd__nand2_2
XFILLER_0_28_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14656_ net848 _06280_ _06860_ _06381_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13607_ _05816_ _05817_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__nand2_1
X_17375_ net354 net358 VGND VGND VPWR VPWR _09362_ sky130_fd_sc_hd__nand2_1
X_14587_ _06742_ _06744_ VGND VGND VPWR VPWR _06793_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19114_ _11083_ _11085_ _11033_ VGND VGND VPWR VPWR _11086_ sky130_fd_sc_hd__mux2_1
X_16326_ _07230_ net444 VGND VGND VPWR VPWR _08416_ sky130_fd_sc_hd__nand2_2
XFILLER_0_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13538_ _05749_ _05750_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19045_ net371 net370 _10495_ VGND VGND VPWR VPWR _11018_ sky130_fd_sc_hd__and3_1
X_13469_ _05483_ _05485_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__and2_1
X_16257_ _08337_ _08347_ VGND VGND VPWR VPWR _08348_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15208_ net542 net470 VGND VGND VPWR VPWR _07307_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16188_ _08277_ _08279_ VGND VGND VPWR VPWR _08280_ sky130_fd_sc_hd__xor2_1
XFILLER_0_50_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15139_ _07220_ _07221_ VGND VGND VPWR VPWR _07238_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19947_ _11431_ _11817_ net177 VGND VGND VPWR VPWR _11818_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19878_ _11742_ _11753_ VGND VGND VPWR VPWR _11754_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18829_ _10801_ _10803_ VGND VGND VPWR VPWR _10805_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21840_ _01398_ _01399_ _01391_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__and3_1
XFILLER_0_179_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21771_ _01331_ _01332_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_188_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23510_ _02920_ VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__clkbuf_1
X_20722_ net268 _12570_ VGND VGND VPWR VPWR _12571_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24490_ _03840_ _03845_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23441_ top0.cordic0.vec\[1\]\[15\] _02868_ _02876_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__a21o_1
X_20653_ _12470_ _12481_ VGND VGND VPWR VPWR _12502_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26160_ spi0.data_packed\[5\] _05300_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23372_ _02791_ _02813_ _02799_ net120 VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_12_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20584_ _12430_ _12431_ _12432_ VGND VGND VPWR VPWR _12433_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25111_ _04457_ _04459_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22323_ _01684_ _01737_ _01804_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__or3_1
X_26091_ _05270_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25042_ _04305_ _04312_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__or2_1
X_22254_ _01803_ _01809_ _01813_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21205_ _13045_ _13048_ VGND VGND VPWR VPWR _13049_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22185_ _01711_ _01718_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__nand2_1
X_21136_ _11739_ net228 VGND VGND VPWR VPWR _12981_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26993_ clknet_leaf_26_clk_sys _00610_ net625 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout420 net421 VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__buf_4
Xfanout431 top0.pid_d.state\[5\] VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__clkbuf_4
Xfanout442 top0.pid_d.state\[1\] VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__buf_2
Xfanout453 net454 VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__clkbuf_2
X_25944_ _05151_ _05156_ _05150_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_21_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21067_ _11787_ _12912_ VGND VGND VPWR VPWR _12913_ sky130_fd_sc_hd__xnor2_1
Xfanout464 net465 VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__buf_4
Xfanout475 net478 VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__clkbuf_4
Xfanout486 net488 VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__buf_2
X_20018_ top0.cordic0.slte0.opA\[5\] _11866_ _11865_ VGND VGND VPWR VPWR _11884_ sky130_fd_sc_hd__o21a_1
XFILLER_0_198_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout497 net498 VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__buf_4
X_25875_ _05083_ _05084_ _05089_ _05093_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__a22o_1
X_24826_ _03161_ _04174_ _03975_ _04177_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__o31a_2
XFILLER_0_198_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24757_ _04108_ _04109_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__xor2_1
X_21969_ _01511_ _01513_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__nand2_1
X_14510_ _05822_ _06716_ _06640_ net28 VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_178_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23708_ net568 top0.matmul0.matmul_stage_inst.b\[2\] top0.matmul0.matmul_stage_inst.a\[2\]
+ net564 VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__a22o_2
XFILLER_0_51_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15490_ _07293_ _07588_ VGND VGND VPWR VPWR _07589_ sky130_fd_sc_hd__nor2_1
X_24688_ _03910_ _03911_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14441_ _06642_ _06647_ VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23639_ net569 top0.matmul0.matmul_stage_inst.b\[6\] top0.matmul0.matmul_stage_inst.a\[6\]
+ net564 VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__a22o_1
X_26427_ clknet_leaf_78_clk_sys _00068_ net632 VGND VGND VPWR VPWR top0.kid\[0\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_30_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout60 top0.periodTop_r\[2\] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_4
Xfanout71 top0.matmul0.op\[1\] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_2
X_14372_ _06574_ _06580_ VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__xnor2_4
Xfanout82 net84 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17160_ _09172_ _09173_ VGND VGND VPWR VPWR _09174_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26358_ spi0.data_packed\[77\] spi0.data_packed\[78\] net690 VGND VGND VPWR VPWR
+ _05411_ sky130_fd_sc_hd__mux2_1
Xfanout93 net94 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_2
X_13323_ net54 VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__inv_2
X_16111_ _08202_ _08203_ VGND VGND VPWR VPWR _08204_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25309_ _04610_ _04654_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17091_ top0.pid_q.curr_error\[4\] _00011_ _09117_ VGND VGND VPWR VPWR _09122_ sky130_fd_sc_hd__and3_1
X_26289_ _05376_ VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13254_ net173 top0.svm0.state\[1\] top0.svm0.state\[0\] VGND VGND VPWR VPWR _05467_
+ sky130_fd_sc_hd__nor3b_4
X_16042_ _08121_ _08135_ VGND VGND VPWR VPWR _08136_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19801_ net259 _11664_ _11667_ VGND VGND VPWR VPWR _11682_ sky130_fd_sc_hd__o21a_1
X_17993_ top0.pid_d.out\[1\] _09978_ net14 VGND VGND VPWR VPWR _09979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19732_ _11612_ _11614_ _11615_ _11448_ _11445_ VGND VGND VPWR VPWR _11616_ sky130_fd_sc_hd__o221a_2
X_16944_ _09000_ _09001_ net547 VGND VGND VPWR VPWR _09002_ sky130_fd_sc_hd__and3b_1
XFILLER_0_193_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19663_ net291 VGND VGND VPWR VPWR _11550_ sky130_fd_sc_hd__inv_2
X_16875_ _08936_ _08922_ _08924_ _08937_ VGND VGND VPWR VPWR _08938_ sky130_fd_sc_hd__a31o_1
X_18614_ _05449_ _10592_ VGND VGND VPWR VPWR _10593_ sky130_fd_sc_hd__and2_1
X_15826_ _07819_ _07824_ _07817_ VGND VGND VPWR VPWR _07922_ sky130_fd_sc_hd__o21a_1
X_19594_ _11468_ _11473_ _11477_ _11482_ VGND VGND VPWR VPWR _11483_ sky130_fd_sc_hd__or4_4
XFILLER_0_56_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18545_ net390 net312 VGND VGND VPWR VPWR _10524_ sky130_fd_sc_hd__nand2_1
X_15757_ _07754_ _07755_ _07756_ VGND VGND VPWR VPWR _07854_ sky130_fd_sc_hd__o21a_1
XFILLER_0_176_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14708_ _06876_ VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__inv_2
X_18476_ net344 net348 VGND VGND VPWR VPWR _10456_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15688_ net481 _07784_ _07785_ VGND VGND VPWR VPWR _07786_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_173_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17427_ net413 net340 VGND VGND VPWR VPWR _09414_ sky130_fd_sc_hd__and2_2
X_14639_ _06840_ _06843_ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_51_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17358_ net417 net343 VGND VGND VPWR VPWR _09345_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16309_ net545 _08328_ _08329_ net548 _08399_ VGND VGND VPWR VPWR _08400_ sky130_fd_sc_hd__a32o_1
X_17289_ _09285_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19028_ net316 _10384_ _10074_ VGND VGND VPWR VPWR _11001_ sky130_fd_sc_hd__nand3_1
XFILLER_0_152_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23990_ _03317_ _03318_ _03347_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__a21o_1
X_22941_ _02306_ _02454_ _02309_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22872_ top0.svm0.tB\[7\] _02390_ net170 VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__o21ba_1
X_25660_ net71 _04933_ _04934_ net74 _04878_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__a221o_1
X_24611_ _03948_ _03952_ _03964_ VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__o21ba_1
X_21823_ net130 net1031 VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__nand2_2
X_25591_ net69 VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_174_Right_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24542_ _03887_ _03896_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__xnor2_2
X_21754_ _01298_ _01315_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_149_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20705_ net301 net296 VGND VGND VPWR VPWR _12554_ sky130_fd_sc_hd__nor2_1
X_24473_ _03828_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27261_ clknet_3_0__leaf_clk_mosi _00875_ VGND VGND VPWR VPWR spi0.data_packed\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_21685_ _01229_ _01246_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_11_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23424_ _02858_ _02861_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__xor2_1
X_26212_ spi0.data_packed\[4\] spi0.data_packed\[5\] net694 VGND VGND VPWR VPWR _05338_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27192_ clknet_leaf_56_clk_sys _00806_ net668 VGND VGND VPWR VPWR top0.currT_r\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_20636_ _12480_ _12482_ VGND VGND VPWR VPWR _12485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26143_ _05287_ top0.cordic0.slte0.opB\[3\] _12006_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23355_ _11513_ _02797_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20567_ _12411_ _12414_ VGND VGND VPWR VPWR _12416_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22306_ _01863_ _01865_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__xnor2_2
X_26074_ top0.a_in_matmul\[10\] _05257_ _05230_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__mux2_1
X_23286_ _02730_ _02733_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__xor2_2
X_20498_ net295 net287 VGND VGND VPWR VPWR _12347_ sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_72_clk_sys clknet_3_5__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_72_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_25025_ _04368_ _04374_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__xnor2_2
X_22237_ _01643_ net95 VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__nor2_1
X_22168_ _01249_ _01247_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__nand2_1
X_21119_ _12897_ _12933_ _12892_ VGND VGND VPWR VPWR _12964_ sky130_fd_sc_hd__o21a_1
X_26976_ clknet_leaf_28_clk_sys _00593_ net622 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_14990_ spi0.data_packed\[1\] top0.periodTop\[1\] _07108_ VGND VGND VPWR VPWR _07120_
+ sky130_fd_sc_hd__mux2_1
Xfanout250 top0.cordic0.vec\[0\]\[10\] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__buf_2
X_22099_ _01653_ _01660_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__nor2_1
Xfanout261 net262 VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout272 net273 VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__buf_2
X_13941_ _06152_ _06153_ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__and2b_1
X_25927_ _05138_ _05141_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__xnor2_1
Xfanout283 net284 VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__buf_2
Xfanout294 net295 VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__buf_2
XFILLER_0_191_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16660_ _08690_ _08735_ _08736_ VGND VGND VPWR VPWR _08745_ sky130_fd_sc_hd__a21bo_1
X_13872_ _05751_ _05785_ _06084_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__o21a_2
X_25858_ _05439_ _05065_ _05078_ _05067_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_201_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15611_ net1019 VGND VGND VPWR VPWR _07710_ sky130_fd_sc_hd__buf_4
XFILLER_0_202_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24809_ _04159_ _04160_ VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__or2b_1
X_16591_ _08676_ _08677_ VGND VGND VPWR VPWR _08678_ sky130_fd_sc_hd__nand2_1
XFILLER_0_198_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25789_ net208 _05009_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18330_ _10311_ _10210_ _10211_ VGND VGND VPWR VPWR _10312_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15542_ _07639_ _07640_ VGND VGND VPWR VPWR _07641_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18261_ net434 _10161_ _10243_ net436 _07138_ VGND VGND VPWR VPWR _10244_ sky130_fd_sc_hd__a221o_1
X_15473_ _07282_ _07570_ _07571_ VGND VGND VPWR VPWR _07572_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_84_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17212_ net548 _09029_ _09219_ net554 VGND VGND VPWR VPWR _09220_ sky130_fd_sc_hd__a22o_1
X_14424_ _06565_ _06630_ _06631_ VGND VGND VPWR VPWR _06632_ sky130_fd_sc_hd__o21a_2
XFILLER_0_182_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18192_ net328 net388 VGND VGND VPWR VPWR _10175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17143_ _09157_ _09158_ VGND VGND VPWR VPWR _09159_ sky130_fd_sc_hd__nand2_1
X_14355_ _06562_ _06563_ VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_181_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13306_ net49 net1015 VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__nand2_2
XFILLER_0_24_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14286_ _05565_ _05608_ _05609_ VGND VGND VPWR VPWR _06496_ sky130_fd_sc_hd__or3_2
X_17074_ _08403_ _09111_ VGND VGND VPWR VPWR _09112_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16025_ _08113_ _08118_ VGND VGND VPWR VPWR _08119_ sky130_fd_sc_hd__xnor2_1
X_13237_ _05454_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__buf_1
XFILLER_0_21_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17976_ _09874_ _09877_ VGND VGND VPWR VPWR _09962_ sky130_fd_sc_hd__nand2_1
X_19715_ _11451_ _11446_ _11594_ net84 _11599_ VGND VGND VPWR VPWR _11600_ sky130_fd_sc_hd__a221o_1
X_16927_ top0.currT_r\[8\] _08985_ VGND VGND VPWR VPWR _08986_ sky130_fd_sc_hd__xnor2_1
X_19646_ _11408_ _11438_ _11424_ _11452_ _11511_ VGND VGND VPWR VPWR _11534_ sky130_fd_sc_hd__o2111ai_4
X_16858_ _08908_ _08909_ _08921_ VGND VGND VPWR VPWR _08922_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15809_ _07810_ _07893_ _07892_ VGND VGND VPWR VPWR _07905_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19577_ top0.cordic0.slte0.opA\[12\] top0.cordic0.slte0.opB\[12\] VGND VGND VPWR
+ VPWR _11466_ sky130_fd_sc_hd__and2b_1
X_16789_ top0.kiq\[4\] _08863_ _08866_ VGND VGND VPWR VPWR _08868_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18528_ _10434_ _10507_ VGND VGND VPWR VPWR _10508_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18459_ _10436_ _10438_ VGND VGND VPWR VPWR _10439_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21470_ _00977_ _01008_ net218 VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20421_ _12267_ _12269_ net269 VGND VGND VPWR VPWR _12270_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23140_ _02598_ _02628_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20352_ net283 net276 VGND VGND VPWR VPWR _12201_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23071_ _02570_ _02571_ net46 VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__a21o_1
X_20283_ _12130_ _12131_ VGND VGND VPWR VPWR _12132_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22022_ net152 net136 VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26830_ clknet_leaf_43_clk_sys _00447_ net680 VGND VGND VPWR VPWR top0.svm0.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold14 top0.matmul0.matmul_stage_inst.c\[13\] VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold25 top0.matmul0.matmul_stage_inst.d\[7\] VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 top0.svm0.tC\[0\] VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 top0.matmul0.matmul_stage_inst.d\[4\] VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 top0.pid_q.prev_error\[15\] VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__dlygate4sd3_1
X_26761_ clknet_leaf_7_clk_sys _00378_ net593 VGND VGND VPWR VPWR top0.cordic0.domain\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_23973_ _03237_ _03246_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__xnor2_1
Xhold69 top0.cordic0.sin\[7\] VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__dlygate4sd3_1
X_25712_ net784 _04964_ _04936_ _04972_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__a22o_1
X_22924_ _02439_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__buf_2
XFILLER_0_39_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26692_ clknet_leaf_83_clk_sys _00309_ net641 VGND VGND VPWR VPWR top0.pid_d.curr_error\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25643_ top0.matmul0.sin\[4\] _04914_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__nor2_1
X_22855_ _02374_ top0.svm0.tA\[12\] _02319_ _02318_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21806_ net147 _01294_ net162 VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__mux2_1
X_22786_ _07115_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_151_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25574_ _04874_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24525_ _03809_ _03869_ _03804_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_148_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21737_ net147 net142 VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__nand2_2
XFILLER_0_66_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27244_ clknet_3_5__leaf_clk_mosi _00858_ VGND VGND VPWR VPWR spi0.data_packed\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24456_ _03804_ _03811_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21668_ net88 VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_164_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20619_ net288 net282 VGND VGND VPWR VPWR _12468_ sky130_fd_sc_hd__nor2_1
X_23407_ _02835_ _02836_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__or2_1
X_24387_ _03161_ _03743_ VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__nor2_1
X_27175_ clknet_leaf_32_clk_sys _00789_ net618 VGND VGND VPWR VPWR top0.periodTop_r\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_62_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21599_ _01141_ _01145_ _01134_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14140_ _06351_ _06193_ _06191_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26126_ spi0.data_packed\[21\] _05281_ _05282_ net905 VGND VGND VPWR VPWR _00802_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23338_ net134 _02780_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14071_ net1025 _05726_ _05727_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23269_ net1016 _02716_ _02708_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__or3_1
X_26057_ top0.matmul0.alpha_pass\[6\] _05237_ _05244_ VGND VGND VPWR VPWR _05245_
+ sky130_fd_sc_hd__a21o_1
X_25008_ _04356_ _04357_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__xnor2_1
X_17830_ _09809_ _09816_ VGND VGND VPWR VPWR _09817_ sky130_fd_sc_hd__xnor2_1
X_17761_ _09406_ _09368_ _09446_ VGND VGND VPWR VPWR _09748_ sky130_fd_sc_hd__a21bo_1
X_26959_ clknet_leaf_15_clk_sys _00576_ net613 VGND VGND VPWR VPWR top0.matmul0.b\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14973_ spi0.data_packed\[28\] top0.kiq\[12\] _07108_ VGND VGND VPWR VPWR _07109_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19500_ top0.pid_d.curr_int\[13\] top0.pid_d.prev_int\[13\] VGND VGND VPWR VPWR _11392_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_57_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16712_ top0.pid_q.out\[14\] _07705_ _08796_ net544 VGND VGND VPWR VPWR _08797_ sky130_fd_sc_hd__a22o_1
X_13924_ _06133_ _06136_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__xnor2_1
X_17692_ net398 net345 net349 net392 VGND VGND VPWR VPWR _09679_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_199_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19431_ top0.pid_d.curr_int\[6\] top0.pid_d.prev_int\[6\] VGND VGND VPWR VPWR _11331_
+ sky130_fd_sc_hd__xor2_1
X_16643_ _08662_ _08666_ _08660_ VGND VGND VPWR VPWR _08729_ sky130_fd_sc_hd__a21o_1
X_13855_ _06020_ _06017_ _06012_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19362_ net433 _07137_ _05441_ VGND VGND VPWR VPWR _11284_ sky130_fd_sc_hd__o21a_2
XFILLER_0_186_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16574_ _08582_ _08585_ _08579_ VGND VGND VPWR VPWR _08661_ sky130_fd_sc_hd__a21o_1
X_13786_ _05996_ _05997_ _05998_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18313_ _10168_ _10170_ _10294_ VGND VGND VPWR VPWR _10295_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15525_ net478 net514 VGND VGND VPWR VPWR _07624_ sky130_fd_sc_hd__nand2_2
X_19293_ top0.pid_d.prev_error\[12\] top0.pid_d.curr_error\[12\] VGND VGND VPWR VPWR
+ _11235_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18244_ net421 net310 _10082_ _10226_ VGND VGND VPWR VPWR _10227_ sky130_fd_sc_hd__a31o_1
X_15456_ _07267_ _07268_ _07269_ VGND VGND VPWR VPWR _07555_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14407_ net45 _06131_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__nand2_2
XFILLER_0_167_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18175_ top0.pid_d.curr_int\[3\] _10069_ top0.pid_d.out\[3\] VGND VGND VPWR VPWR
+ _10158_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15387_ _07438_ _07483_ _07182_ _07484_ _07485_ VGND VGND VPWR VPWR _07486_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_108_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17126_ top0.pid_q.curr_int\[0\] top0.pid_q.prev_int\[0\] _09142_ VGND VGND VPWR
+ VPWR _09144_ sky130_fd_sc_hd__nand3_1
XFILLER_0_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14338_ _06178_ _06384_ _06472_ _06545_ VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__nand4bb_4
XFILLER_0_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17057_ top0.pid_q.curr_error\[3\] _09100_ _09102_ _08920_ VGND VGND VPWR VPWR _00184_
+ sky130_fd_sc_hd__a22o_1
X_14269_ _06419_ _06420_ _06477_ _06478_ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__or4_2
XFILLER_0_0_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16008_ net453 net521 VGND VGND VPWR VPWR _08102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17959_ _09943_ _09944_ VGND VGND VPWR VPWR _09945_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_174_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20970_ net231 _12698_ _12814_ _12816_ VGND VGND VPWR VPWR _12817_ sky130_fd_sc_hd__a211o_1
XFILLER_0_174_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_20_clk_sys clknet_3_2__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_20_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_196_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19629_ net1016 VGND VGND VPWR VPWR _11518_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_178_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22640_ _01924_ _01821_ net107 VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22571_ _02124_ _02125_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__and2_1
XFILLER_0_180_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24310_ _03110_ _03130_ _03135_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__o21a_1
X_21522_ _01073_ _01077_ _01083_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_69_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25290_ _04634_ _04628_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__or2b_1
XFILLER_0_134_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24241_ _03595_ _03598_ _03588_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21453_ _00984_ _00986_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20404_ net265 net254 VGND VGND VPWR VPWR _12253_ sky130_fd_sc_hd__xor2_2
XFILLER_0_32_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24172_ _03411_ _03529_ _03413_ _03414_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__o211ai_1
X_21384_ _11789_ _13129_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__nor2_1
XFILLER_0_189_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23123_ _07117_ _02616_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20335_ _12181_ _12182_ _12183_ VGND VGND VPWR VPWR _12184_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23054_ _05500_ top0.svm0.counter\[12\] _02550_ _02554_ VGND VGND VPWR VPWR _02555_
+ sky130_fd_sc_hd__a31o_1
X_20266_ _12113_ _12114_ VGND VGND VPWR VPWR _12115_ sky130_fd_sc_hd__nor2_2
XFILLER_0_101_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22005_ _01564_ _01566_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__xnor2_1
X_20197_ _12042_ _12045_ net267 VGND VGND VPWR VPWR _12046_ sky130_fd_sc_hd__o21bai_2
X_26813_ clknet_leaf_67_clk_sys _00430_ net660 VGND VGND VPWR VPWR top0.pid_q.prev_int\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_26744_ clknet_leaf_96_clk_sys _00361_ net588 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_23956_ _03045_ _03046_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__or2_1
X_22907_ net169 _02409_ _02424_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_196_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26675_ clknet_leaf_81_clk_sys _00292_ net636 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_23887_ _03011_ _03060_ _03243_ _03244_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13640_ _05809_ _05850_ _05852_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__a21o_1
X_25626_ _04884_ top0.matmul0.sin\[1\] top0.matmul0.sin\[0\] VGND VGND VPWR VPWR _04906_
+ sky130_fd_sc_hd__and3_1
X_22838_ _02338_ _02344_ _02351_ _02357_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13571_ _05772_ _05783_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__xnor2_1
X_25557_ _04865_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_4_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22769_ top0.pid_q.prev_int\[13\] _02291_ _02294_ top0.pid_q.curr_int\[13\] VGND
+ VGND VPWR VPWR _00432_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15310_ net542 net471 _07407_ VGND VGND VPWR VPWR _07409_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24508_ _03859_ _03860_ _03862_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__or3_2
XFILLER_0_54_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16290_ _08348_ _08380_ VGND VGND VPWR VPWR _08381_ sky130_fd_sc_hd__xnor2_2
X_25488_ top0.matmul0.matmul_stage_inst.mult1\[0\] _03641_ _04829_ VGND VGND VPWR
+ VPWR _04830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15241_ net522 _07314_ _07313_ VGND VGND VPWR VPWR _07340_ sky130_fd_sc_hd__or3_1
X_27227_ clknet_3_4__leaf_clk_mosi _00841_ VGND VGND VPWR VPWR spi0.data_packed\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_24439_ _03788_ _03789_ _03794_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15172_ _07267_ _07270_ VGND VGND VPWR VPWR _07271_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_90_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27158_ clknet_leaf_9_clk_sys _00772_ net596 VGND VGND VPWR VPWR top0.a_in_matmul\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14123_ net1030 _06023_ VGND VGND VPWR VPWR _06335_ sky130_fd_sc_hd__nand2_1
X_26109_ top0.periodTop\[8\] _05276_ _05278_ net43 VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19980_ _11484_ _11504_ _11847_ VGND VGND VPWR VPWR _11848_ sky130_fd_sc_hd__a21oi_1
X_27089_ clknet_leaf_1_clk_sys _00706_ net584 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18931_ _10828_ _10829_ VGND VGND VPWR VPWR _10906_ sky130_fd_sc_hd__nand2_1
X_14054_ _06263_ _06133_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18862_ top0.pid_d.out\[11\] _10833_ _10837_ VGND VGND VPWR VPWR _10838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17813_ net393 net345 net349 net388 VGND VGND VPWR VPWR _09800_ sky130_fd_sc_hd__a22oi_1
X_18793_ _10255_ _10768_ _10699_ _10694_ VGND VGND VPWR VPWR _10769_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_118_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17744_ _09424_ _09730_ VGND VGND VPWR VPWR _09731_ sky130_fd_sc_hd__nand2_1
X_14956_ spi0.data_packed\[20\] top0.kiq\[4\] _07097_ VGND VGND VPWR VPWR _07100_
+ sky130_fd_sc_hd__mux2_1
X_13907_ _06118_ _06102_ _06103_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__and3_1
XFILLER_0_199_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17675_ _09652_ _09661_ VGND VGND VPWR VPWR _09662_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14887_ _07063_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__clkbuf_1
X_19414_ top0.pid_d.curr_int\[3\] VGND VGND VPWR VPWR _11316_ sky130_fd_sc_hd__inv_2
X_16626_ _08648_ _08711_ VGND VGND VPWR VPWR _08712_ sky130_fd_sc_hd__xor2_1
X_13838_ _06024_ _06049_ _06050_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__o21a_1
XFILLER_0_187_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19345_ _11121_ _11162_ _11278_ _11273_ top0.pid_d.curr_error\[4\] VGND VGND VPWR
+ VPWR _00298_ sky130_fd_sc_hd__a32o_1
X_16557_ _08560_ _08565_ _08558_ VGND VGND VPWR VPWR _08644_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_31_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13769_ _05931_ _05935_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__xor2_1
XFILLER_0_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15508_ _07298_ _07599_ _07606_ VGND VGND VPWR VPWR _07607_ sky130_fd_sc_hd__a21o_1
X_19276_ net438 _11218_ _11219_ VGND VGND VPWR VPWR _11220_ sky130_fd_sc_hd__and3_1
X_16488_ net459 _08573_ _08575_ VGND VGND VPWR VPWR _08576_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18227_ net405 net315 VGND VGND VPWR VPWR _10210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15439_ _07276_ _07537_ VGND VGND VPWR VPWR _07538_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18158_ _09593_ net307 _10140_ VGND VGND VPWR VPWR _10142_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold303 top0.cordic0.sin\[1\] VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__dlygate4sd3_1
X_17109_ top0.pid_q.curr_error\[13\] _08860_ _09116_ VGND VGND VPWR VPWR _09131_ sky130_fd_sc_hd__and3_1
X_18089_ _10053_ _10056_ _10072_ VGND VGND VPWR VPWR _10073_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20120_ top0.cordic0.slte0.opA\[14\] _11970_ _11966_ _11965_ VGND VGND VPWR VPWR
+ _11977_ sky130_fd_sc_hd__a211o_1
XFILLER_0_68_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20051_ net932 _11913_ _11914_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23810_ _03139_ _03141_ _03167_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__and3_1
XFILLER_0_175_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24790_ _04038_ _04045_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__nor2_1
X_23741_ _03073_ _03074_ _03098_ VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__a21o_1
X_20953_ _12782_ _12800_ VGND VGND VPWR VPWR _12801_ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26460_ clknet_leaf_91_clk_sys net701 net600 VGND VGND VPWR VPWR spi0.cs_sync\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_23672_ net572 top0.matmul0.matmul_stage_inst.d\[11\] top0.matmul0.matmul_stage_inst.c\[11\]
+ net556 VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__a22o_4
X_20884_ _12161_ _12192_ _12187_ VGND VGND VPWR VPWR _12733_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25411_ _04701_ _04707_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__nor2_1
XFILLER_0_192_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22623_ _01877_ _02175_ _02176_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__or3b_1
X_26391_ clknet_leaf_38_clk_sys _00032_ net677 VGND VGND VPWR VPWR top0.svm0.tC\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25342_ _04614_ _04615_ _04686_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__o21ba_1
X_22554_ _01074_ _01980_ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21505_ _01065_ _01066_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25273_ _04548_ _04549_ _04618_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22485_ _02038_ _02040_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27012_ clknet_leaf_23_clk_sys _00629_ net626 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_24224_ _03575_ _03578_ _03581_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21436_ _00964_ _00997_ _01001_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_146_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_86_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24155_ _03470_ _03512_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21367_ net231 _13170_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23106_ top0.svm0.delta\[1\] net555 top0.svm0.delta\[2\] top0.svm0.delta\[3\] VGND
+ VGND VPWR VPWR _02604_ sky130_fd_sc_hd__or4_2
X_20318_ _12164_ _12166_ VGND VGND VPWR VPWR _12167_ sky130_fd_sc_hd__xnor2_1
X_24086_ _03328_ _03329_ _03332_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__a21oi_1
X_21298_ _13136_ _13140_ VGND VGND VPWR VPWR _13141_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_101_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23037_ net65 net63 net61 VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__or3_1
X_20249_ _12092_ _12093_ _12097_ VGND VGND VPWR VPWR _12098_ sky130_fd_sc_hd__a21bo_1
X_14810_ _06974_ _06977_ VGND VGND VPWR VPWR _07010_ sky130_fd_sc_hd__or2_1
X_15790_ net508 net481 _07767_ VGND VGND VPWR VPWR _07887_ sky130_fd_sc_hd__a21o_1
X_24988_ _03355_ _04131_ _04337_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_95_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14741_ _06942_ _06943_ VGND VGND VPWR VPWR _06944_ sky130_fd_sc_hd__or2_1
X_26727_ clknet_leaf_104_clk_sys _00344_ net576 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_23939_ _03293_ _03294_ _03287_ _03290_ _03291_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__a311o_1
XFILLER_0_200_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17460_ _09406_ _09446_ VGND VGND VPWR VPWR _09447_ sky130_fd_sc_hd__xnor2_1
X_14672_ net39 _06824_ _06874_ _06875_ VGND VGND VPWR VPWR _06876_ sky130_fd_sc_hd__a31o_1
X_26658_ clknet_leaf_77_clk_sys _00275_ net635 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16411_ _08496_ _08499_ VGND VGND VPWR VPWR _08500_ sky130_fd_sc_hd__xnor2_2
X_13623_ _05816_ _05817_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__xnor2_1
X_25609_ _05457_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__clkbuf_4
X_17391_ net423 top0.pid_d.mult0.a\[0\] _09377_ VGND VGND VPWR VPWR _09378_ sky130_fd_sc_hd__and3_1
XFILLER_0_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26589_ clknet_leaf_54_clk_sys _00212_ net669 VGND VGND VPWR VPWR top0.pid_q.prev_error\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19130_ _11099_ VGND VGND VPWR VPWR _11100_ sky130_fd_sc_hd__buf_2
X_16342_ net463 net501 VGND VGND VPWR VPWR _08432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13554_ _05765_ _05766_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__xor2_1
XFILLER_0_183_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19061_ top0.pid_d.out\[14\] top0.pid_d.curr_int\[14\] VGND VGND VPWR VPWR _11034_
+ sky130_fd_sc_hd__xor2_1
X_16273_ _08261_ _08266_ _08363_ VGND VGND VPWR VPWR _08364_ sky130_fd_sc_hd__o21a_1
XFILLER_0_180_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13485_ _05530_ _05543_ _05545_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__or3_1
X_18012_ _09993_ _09996_ VGND VGND VPWR VPWR _09997_ sky130_fd_sc_hd__xnor2_1
X_15224_ net487 _07321_ _07322_ VGND VGND VPWR VPWR _07323_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15155_ _07252_ _07210_ VGND VGND VPWR VPWR _07254_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14106_ _06315_ _06316_ _06310_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19963_ net992 _11831_ _11832_ _11830_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__a22o_1
X_15086_ _07177_ _07180_ _07184_ VGND VGND VPWR VPWR _07185_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_201_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14037_ _06246_ _06249_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__xnor2_1
X_18914_ _10887_ _10888_ VGND VGND VPWR VPWR _10889_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19894_ net227 _11435_ _11767_ VGND VGND VPWR VPWR _11769_ sky130_fd_sc_hd__and3_1
X_18845_ _10808_ _10820_ VGND VGND VPWR VPWR _10821_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18776_ _10751_ _10752_ VGND VGND VPWR VPWR _10753_ sky130_fd_sc_hd__or2b_1
X_15988_ top0.pid_q.curr_int\[4\] _08078_ top0.pid_q.out\[4\] VGND VGND VPWR VPWR
+ _08082_ sky130_fd_sc_hd__a21o_1
XFILLER_0_171_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17727_ _09702_ _09705_ _09713_ VGND VGND VPWR VPWR _09714_ sky130_fd_sc_hd__and3_1
X_14939_ spi0.data_packed\[44\] top0.kid\[12\] _07086_ VGND VGND VPWR VPWR _07091_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17658_ net382 _09362_ _09498_ VGND VGND VPWR VPWR _09645_ sky130_fd_sc_hd__or3_2
XFILLER_0_58_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16609_ net449 net500 VGND VGND VPWR VPWR _08695_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17589_ net425 _09522_ _09523_ VGND VGND VPWR VPWR _09576_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19328_ top0.pid_d.prev_error\[15\] top0.pid_d.curr_error\[15\] VGND VGND VPWR VPWR
+ _11267_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19259_ _11203_ _11196_ top0.pid_d.prev_error\[8\] VGND VGND VPWR VPWR _11204_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_169_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22270_ net77 _01822_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold100 top0.svm0.tA\[15\] VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21221_ _13063_ _13064_ _13056_ _13058_ VGND VGND VPWR VPWR _13065_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold111 top0.svm0.tA\[3\] VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 top0.matmul0.matmul_stage_inst.c\[4\] VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 top0.c_out_calc\[0\] VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold144 top0.c_out_calc\[11\] VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__dlygate4sd3_1
X_21152_ _12995_ _12996_ VGND VGND VPWR VPWR _12997_ sky130_fd_sc_hd__or2b_1
Xhold155 top0.svm0.tC\[3\] VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold166 top0.matmul0.matmul_stage_inst.b\[5\] VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 _00318_ VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 top0.c_out_calc\[7\] VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__dlygate4sd3_1
X_20103_ _11857_ _11961_ VGND VGND VPWR VPWR _11962_ sky130_fd_sc_hd__nor2_1
Xhold199 top0.pid_q.prev_error\[3\] VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 net605 VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__buf_2
Xfanout613 net614 VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__clkbuf_4
X_21083_ _11788_ _12851_ _12928_ _11758_ net229 VGND VGND VPWR VPWR _12929_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25960_ top0.pid_q.out\[0\] _12032_ _05014_ spi0.data_packed\[48\] VGND VGND VPWR
+ VPWR _05170_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout624 net629 VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__buf_2
Xfanout635 net654 VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__buf_2
XFILLER_0_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24911_ _04257_ _04261_ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__xnor2_4
X_20034_ _11431_ _11898_ net178 VGND VGND VPWR VPWR _11899_ sky130_fd_sc_hd__o21ai_1
Xfanout646 net649 VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout657 net658 VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__clkbuf_4
X_25891_ _05102_ _05108_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__xnor2_1
Xfanout668 net669 VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout679 net686 VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__clkbuf_4
X_24842_ _04187_ _04193_ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24773_ _03991_ _03992_ _04028_ _04029_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__a211o_1
X_21985_ _01454_ _01480_ _01543_ _01546_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__a211o_1
X_26512_ clknet_leaf_66_clk_sys _00135_ net659 VGND VGND VPWR VPWR top0.pid_q.out\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_23724_ _03078_ _03081_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__xnor2_4
X_20936_ _12783_ _12708_ VGND VGND VPWR VPWR _12784_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26443_ clknet_leaf_87_clk_sys _00084_ net644 VGND VGND VPWR VPWR top0.kiq\[0\] sky130_fd_sc_hd__dfrtp_1
X_23655_ _03010_ _03011_ _03009_ _03012_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__a31o_1
X_20867_ _12714_ _12715_ VGND VGND VPWR VPWR _12716_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22606_ _02154_ _02159_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__or2b_1
XFILLER_0_193_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26374_ spi0.opcode\[5\] spi0.opcode\[6\] net696 VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23586_ top0.matmul0.alpha_pass\[0\] _09251_ net560 VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__mux2_1
X_20798_ _12644_ _12645_ _12646_ VGND VGND VPWR VPWR _12647_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_113_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25325_ _04272_ _04288_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22537_ net726 _12004_ _12740_ _02092_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25256_ _04601_ _04602_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__and2b_1
X_13270_ top0.matmul0.alpha_pass\[0\] _05435_ _05474_ VGND VGND VPWR VPWR _05483_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_17_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22468_ net92 _01769_ _02023_ _02024_ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__a211o_1
X_24207_ _03564_ _03161_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__nor2_1
X_21419_ _00933_ _00985_ _00947_ net218 VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__o2bb2a_1
X_25187_ _04533_ _04534_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__xnor2_1
X_22399_ _01143_ _01259_ _01954_ net119 _01956_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24138_ _02998_ _03000_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__nor2_2
X_16960_ top0.pid_q.curr_error\[9\] VGND VGND VPWR VPWR _09017_ sky130_fd_sc_hd__inv_2
X_24069_ _03335_ _03426_ _03374_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15911_ net483 net502 _07485_ VGND VGND VPWR VPWR _08006_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16891_ _08951_ _08952_ VGND VGND VPWR VPWR _08953_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_188_Right_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18630_ _10573_ _10577_ _10607_ VGND VGND VPWR VPWR _10608_ sky130_fd_sc_hd__a21oi_1
X_15842_ net455 net523 VGND VGND VPWR VPWR _07938_ sky130_fd_sc_hd__nand2_2
X_18561_ _10538_ _10539_ VGND VGND VPWR VPWR _10540_ sky130_fd_sc_hd__xor2_1
X_15773_ _07732_ _07736_ _07734_ VGND VGND VPWR VPWR _07870_ sky130_fd_sc_hd__a21o_1
X_17512_ net390 net386 net358 net401 VGND VGND VPWR VPWR _09499_ sky130_fd_sc_hd__or4bb_1
X_14724_ _06832_ _05731_ VGND VGND VPWR VPWR _06927_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_67_clk_sys clknet_3_5__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_67_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_108_clk_sys clknet_3_0__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_108_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_18492_ net338 net364 VGND VGND VPWR VPWR _10472_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17443_ net395 _09428_ _09429_ net352 VGND VGND VPWR VPWR _09430_ sky130_fd_sc_hd__a2bb2o_1
X_14655_ _06817_ _06859_ VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_86_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13606_ top0.periodTop_r\[4\] _05517_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17374_ net357 _09358_ _09359_ _09360_ VGND VGND VPWR VPWR _09361_ sky130_fd_sc_hd__a22oi_2
X_14586_ _06749_ _06791_ VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__xor2_4
XFILLER_0_172_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19113_ top0.pid_d.out\[14\] top0.pid_d.curr_int\[14\] _11084_ VGND VGND VPWR VPWR
+ _11085_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16325_ _08351_ _08353_ _08414_ VGND VGND VPWR VPWR _08415_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_40_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13537_ _05747_ _05748_ _05742_ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19044_ net377 _10494_ _10964_ VGND VGND VPWR VPWR _11017_ sky130_fd_sc_hd__or3b_2
XFILLER_0_54_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16256_ _08339_ _08346_ VGND VGND VPWR VPWR _08347_ sky130_fd_sc_hd__xnor2_1
X_13468_ _05677_ _05680_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15207_ net539 net471 VGND VGND VPWR VPWR _07306_ sky130_fd_sc_hd__nand2_1
X_16187_ _08202_ _08203_ _08278_ VGND VGND VPWR VPWR _08279_ sky130_fd_sc_hd__a21oi_2
X_13399_ top0.matmul0.beta_pass\[9\] _05435_ _05470_ _05464_ top0.c_out_calc\[9\]
+ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_3_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15138_ _07220_ _07221_ _07236_ VGND VGND VPWR VPWR _07237_ sky130_fd_sc_hd__or3b_1
XFILLER_0_26_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19946_ _11802_ _11816_ VGND VGND VPWR VPWR _11817_ sky130_fd_sc_hd__xor2_1
X_15069_ _07152_ _07167_ VGND VGND VPWR VPWR _07168_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_120_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19877_ _11713_ _11743_ _11744_ _11752_ VGND VGND VPWR VPWR _11753_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18828_ _10801_ _10803_ VGND VGND VPWR VPWR _10804_ sky130_fd_sc_hd__nand2_1
X_18759_ _10616_ _10617_ VGND VGND VPWR VPWR _10736_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21770_ _01175_ _01259_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_72_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20721_ _11593_ _12569_ VGND VGND VPWR VPWR _12570_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20652_ _12497_ _12500_ VGND VGND VPWR VPWR _12501_ sky130_fd_sc_hd__xnor2_2
X_23440_ net94 _02868_ _02869_ _02870_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23371_ _01217_ _02811_ _02812_ _01408_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__a31o_1
X_20583_ net302 _12264_ VGND VGND VPWR VPWR _12432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25110_ _04382_ _04458_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22322_ net749 _12034_ _12037_ _01881_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__a31o_1
X_26090_ top0.a_in_matmul\[14\] _05269_ _05164_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25041_ _04381_ _04390_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__xnor2_2
X_22253_ _01803_ _01809_ _01742_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__o21a_1
XFILLER_0_182_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21204_ _13046_ _13047_ _11789_ VGND VGND VPWR VPWR _13048_ sky130_fd_sc_hd__a21o_1
XFILLER_0_197_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22184_ _01695_ _01743_ _01744_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__o21a_2
XFILLER_0_197_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21135_ net272 _12975_ _12979_ VGND VGND VPWR VPWR _12980_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26992_ clknet_leaf_26_clk_sys _00609_ net627 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout410 net414 VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__clkbuf_4
Xfanout421 top0.pid_d.mult0.a\[2\] VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__clkbuf_2
Xfanout432 net434 VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__clkbuf_4
X_25943_ _05439_ _05155_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__nand2_1
Xfanout443 top0.pid_q.mult0.b\[15\] VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__buf_4
X_21066_ _11757_ _12911_ _12832_ VGND VGND VPWR VPWR _12912_ sky130_fd_sc_hd__o21a_1
Xfanout454 top0.pid_q.mult0.b\[11\] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__clkbuf_4
Xfanout465 top0.pid_q.mult0.b\[7\] VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__clkbuf_4
Xfanout476 net477 VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__clkbuf_4
X_20017_ _11837_ _11838_ _11853_ _11881_ _11882_ VGND VGND VPWR VPWR _11883_ sky130_fd_sc_hd__o32a_1
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout487 net488 VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__clkbuf_4
X_25874_ _05082_ _05083_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__nand2_1
Xfanout498 net499 VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__clkbuf_4
X_24825_ _03549_ _04176_ _03829_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__o21a_2
XFILLER_0_96_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24756_ _03024_ _03025_ _03061_ _03062_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_169_Left_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21968_ _01523_ _01527_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23707_ _03061_ _03062_ _03063_ _03064_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__o22a_2
XFILLER_0_68_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20919_ net236 _12761_ _12762_ VGND VGND VPWR VPWR _12767_ sky130_fd_sc_hd__or3b_1
X_24687_ _03572_ _04040_ _03549_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21899_ _01459_ _01460_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14440_ _06642_ _06647_ VGND VGND VPWR VPWR _06648_ sky130_fd_sc_hd__and2_1
X_26426_ clknet_leaf_88_clk_sys _00067_ net642 VGND VGND VPWR VPWR top0.kpq\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_23638_ _02995_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_193_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout50 top0.periodTop_r\[6\] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_4
Xfanout61 top0.periodTop_r\[2\] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_4
Xfanout72 net73 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_2
XFILLER_0_65_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14371_ _06576_ _06579_ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout83 net84 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
X_26357_ _05410_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23569_ _02951_ VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout94 top0.cordic0.vec\[1\]\[15\] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_4
XFILLER_0_88_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16110_ net463 net510 VGND VGND VPWR VPWR _08203_ sky130_fd_sc_hd__nand2_1
X_25308_ _04650_ _04653_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_181_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13322_ _05530_ _05534_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17090_ net899 _09115_ _09121_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26288_ spi0.data_packed\[42\] net1011 net689 VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16041_ _08130_ _08134_ VGND VGND VPWR VPWR _08135_ sky130_fd_sc_hd__xnor2_1
X_25239_ _04585_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__inv_2
X_13253_ _05433_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_178_Left_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19800_ net259 _11664_ _11665_ _11666_ _11621_ VGND VGND VPWR VPWR _11681_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_202_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17992_ net434 _09900_ _09901_ _09977_ net439 VGND VGND VPWR VPWR _09978_ sky130_fd_sc_hd__a32o_1
XFILLER_0_102_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16943_ _08998_ _08999_ _08997_ VGND VGND VPWR VPWR _09001_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19731_ _11536_ _11537_ _11573_ VGND VGND VPWR VPWR _11615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16874_ top0.pid_q.prev_error\[3\] VGND VGND VPWR VPWR _08937_ sky130_fd_sc_hd__inv_2
X_19662_ net174 _11525_ _11547_ _11549_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__a31o_1
X_18613_ top0.pid_d.out\[8\] _10591_ net14 VGND VGND VPWR VPWR _10592_ sky130_fd_sc_hd__mux2_1
X_15825_ _07855_ _07857_ _07920_ VGND VGND VPWR VPWR _07921_ sky130_fd_sc_hd__o21ai_1
X_19593_ _11478_ _11479_ _11480_ _11481_ VGND VGND VPWR VPWR _11482_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_187_Left_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18544_ net317 _10521_ _10522_ _10208_ VGND VGND VPWR VPWR _10523_ sky130_fd_sc_hd__a22o_1
X_15756_ _07849_ _07852_ VGND VGND VPWR VPWR _07853_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14707_ _06862_ _06905_ _06908_ _06909_ VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__o211a_2
XFILLER_0_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18475_ _10449_ _10454_ VGND VGND VPWR VPWR _10455_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15687_ net511 net480 _07663_ _07779_ VGND VGND VPWR VPWR _07785_ sky130_fd_sc_hd__a211o_1
XFILLER_0_185_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17426_ _09411_ _09412_ VGND VGND VPWR VPWR _09413_ sky130_fd_sc_hd__xor2_4
XFILLER_0_74_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14638_ _06841_ _06842_ VGND VGND VPWR VPWR _06843_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17357_ _09340_ _09341_ _09343_ VGND VGND VPWR VPWR _09344_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14569_ _06706_ _06711_ _06774_ VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16308_ _08397_ _08398_ VGND VGND VPWR VPWR _08399_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17288_ top0.matmul0.beta_pass\[6\] _09284_ net562 VGND VGND VPWR VPWR _09285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19027_ _10944_ _10947_ VGND VGND VPWR VPWR _11000_ sky130_fd_sc_hd__and2b_1
X_16239_ _08231_ _08249_ _08317_ VGND VGND VPWR VPWR _08330_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19929_ top0.cordic0.slte0.opA\[0\] _11785_ VGND VGND VPWR VPWR _11801_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22940_ top0.svm0.delta\[3\] _02453_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_177_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22871_ _02324_ top0.svm0.tB\[6\] _02389_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24610_ _03948_ _03952_ _03950_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_195_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21822_ _01379_ _01383_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25590_ _04883_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__buf_2
XFILLER_0_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24541_ _03894_ _03895_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21753_ _01309_ _01314_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__xnor2_1
X_20704_ net292 net278 VGND VGND VPWR VPWR _12553_ sky130_fd_sc_hd__xnor2_4
X_27260_ clknet_3_3__leaf_clk_mosi _00874_ VGND VGND VPWR VPWR spi0.data_packed\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_24472_ _03741_ _03827_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21684_ _01242_ _01245_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__xor2_2
XFILLER_0_191_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26211_ _05337_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23423_ _02851_ _02859_ _02860_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__a21o_1
X_27191_ clknet_leaf_56_clk_sys _00805_ net668 VGND VGND VPWR VPWR top0.currT_r\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_20635_ _12480_ _12483_ _12477_ VGND VGND VPWR VPWR _12484_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26142_ spi0.data_packed\[1\] _05286_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20566_ _12411_ _12414_ VGND VGND VPWR VPWR _12415_ sky130_fd_sc_hd__xor2_1
X_23354_ _02788_ _02789_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22305_ _01748_ _01794_ _01864_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__o21ai_2
Xclkbuf_leaf_15_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_15_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_26073_ top0.matmul0.alpha_pass\[10\] _05237_ _05256_ VGND VGND VPWR VPWR _05257_
+ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_7_clk_sys clknet_3_2__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_7_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_20497_ net298 _12065_ _12156_ net295 _12345_ VGND VGND VPWR VPWR _12346_ sky130_fd_sc_hd__o221a_1
X_23285_ _11484_ _11504_ _11509_ _02732_ VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__a211o_1
X_25024_ _04370_ _04373_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22236_ _01685_ _01686_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__nor2_1
X_22167_ _01722_ _01728_ VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21118_ net718 _12813_ _12962_ _12963_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__a22o_1
X_26975_ clknet_leaf_28_clk_sys _00592_ net622 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_121_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22098_ _01654_ _01655_ _01632_ _01656_ _01659_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__o32a_2
Xfanout240 top0.cordic0.vec\[0\]\[12\] VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_8
Xfanout251 net252 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__buf_4
Xfanout262 top0.cordic0.vec\[0\]\[8\] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__buf_4
X_13940_ _06146_ _06151_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__nand2_1
X_25926_ _05139_ _05140_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__xnor2_1
Xfanout273 top0.cordic0.vec\[0\]\[6\] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__buf_4
X_21049_ net221 _12827_ _11759_ VGND VGND VPWR VPWR _12895_ sky130_fd_sc_hd__a21o_1
Xfanout284 top0.cordic0.vec\[0\]\[4\] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__buf_2
Xfanout295 net297 VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__buf_2
X_13871_ _05752_ _05753_ _05785_ _05751_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__a22o_1
X_25857_ top0.matmul0.alpha_pass\[5\] top0.matmul0.beta_pass\[5\] _05438_ _05070_
+ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__o31a_1
X_15610_ top0.pid_q.out\[0\] _07705_ _07708_ net544 VGND VGND VPWR VPWR _07709_ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24808_ _04035_ _04032_ _03942_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_202_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16590_ _08674_ _08675_ _08673_ VGND VGND VPWR VPWR _08677_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_9_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25788_ net208 _12017_ top0.cordic0.in_valid net205 VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_69_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15541_ net460 net528 VGND VGND VPWR VPWR _07640_ sky130_fd_sc_hd__nand2_1
X_24739_ _03564_ _03719_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18260_ _10165_ _10242_ VGND VGND VPWR VPWR _10243_ sky130_fd_sc_hd__xnor2_1
X_15472_ net531 net462 net464 net528 VGND VGND VPWR VPWR _07571_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_167_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17211_ _09217_ _09218_ VGND VGND VPWR VPWR _09219_ sky130_fd_sc_hd__xnor2_1
X_14423_ _06567_ _06572_ VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__nand2_1
X_26409_ clknet_leaf_85_clk_sys _00050_ net634 VGND VGND VPWR VPWR top0.kpd\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_18191_ _10106_ _10108_ _10173_ VGND VGND VPWR VPWR _10174_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_126_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17142_ top0.pid_q.curr_int\[3\] top0.pid_q.prev_int\[3\] VGND VGND VPWR VPWR _09158_
+ sky130_fd_sc_hd__xnor2_1
X_14354_ net45 _05726_ _05727_ VGND VGND VPWR VPWR _06563_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13305_ _05517_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__buf_1
XFILLER_0_135_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17073_ _09063_ top0.pid_q.curr_error\[13\] _09096_ VGND VGND VPWR VPWR _09111_ sky130_fd_sc_hd__mux2_1
X_14285_ net41 _05602_ _05603_ VGND VGND VPWR VPWR _06495_ sky130_fd_sc_hd__and3_2
XFILLER_0_165_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16024_ _08115_ _08117_ VGND VGND VPWR VPWR _08118_ sky130_fd_sc_hd__xor2_1
XFILLER_0_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13236_ net437 _05441_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17975_ _09858_ _09881_ _09880_ VGND VGND VPWR VPWR _09961_ sky130_fd_sc_hd__a21o_1
X_19714_ net179 _11598_ VGND VGND VPWR VPWR _11599_ sky130_fd_sc_hd__nor2_1
X_16926_ top0.matmul0.beta_pass\[8\] _05436_ VGND VGND VPWR VPWR _08985_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19645_ _11529_ _11532_ _11511_ VGND VGND VPWR VPWR _11533_ sky130_fd_sc_hd__a21o_1
X_16857_ top0.pid_q.curr_error\[2\] VGND VGND VPWR VPWR _08921_ sky130_fd_sc_hd__inv_2
X_15808_ _07901_ _07902_ VGND VGND VPWR VPWR _07904_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19576_ top0.cordic0.slte0.opB\[12\] top0.cordic0.slte0.opA\[12\] VGND VGND VPWR
+ VPWR _11465_ sky130_fd_sc_hd__nor2b_1
X_16788_ net533 _08856_ _08859_ net789 _08867_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15739_ _07834_ _07835_ VGND VGND VPWR VPWR _07836_ sky130_fd_sc_hd__xnor2_1
X_18527_ _10441_ _10506_ VGND VGND VPWR VPWR _10507_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18458_ _10400_ _10409_ _10437_ VGND VGND VPWR VPWR _10438_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17409_ net410 _09352_ _09351_ net357 VGND VGND VPWR VPWR _09396_ sky130_fd_sc_hd__and4_1
XFILLER_0_29_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18389_ _10278_ _10280_ _10279_ VGND VGND VPWR VPWR _10370_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20420_ net267 net262 VGND VGND VPWR VPWR _12269_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20351_ _12136_ _12199_ _11689_ VGND VGND VPWR VPWR _12200_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23070_ _02540_ _02566_ _02564_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__or3b_1
XFILLER_0_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20282_ net296 net269 VGND VGND VPWR VPWR _12131_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_178_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22021_ net136 _01301_ _01487_ net166 VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold15 top0.cordic0.cos\[1\] VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 top0.cordic0.sin\[6\] VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 top0.periodTop\[15\] VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__dlygate4sd3_1
X_26760_ clknet_3_0__leaf_clk_sys _00377_ net589 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_23972_ _03328_ _03329_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__nand2_1
Xhold48 top0.matmul0.matmul_stage_inst.start VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 top0.matmul0.matmul_stage_inst.d\[0\] VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25711_ top0.matmul0.sin\[4\] _04971_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__xnor2_1
X_22923_ net171 _02306_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__nand2_1
X_26691_ clknet_leaf_83_clk_sys _00308_ net641 VGND VGND VPWR VPWR top0.pid_d.curr_error\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_190_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25642_ net847 _04904_ _04917_ _04919_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__a22o_1
X_22854_ top0.svm0.counter\[12\] VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__inv_2
XFILLER_0_195_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21805_ _01331_ _01332_ _01326_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25573_ top0.matmul0.a\[9\] top0.matmul0.matmul_stage_inst.e\[9\] _04867_ VGND VGND
+ VPWR VPWR _04874_ sky130_fd_sc_hd__mux2_1
X_22785_ top0.svm0.state\[0\] VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__inv_4
XFILLER_0_79_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24524_ _03868_ _03878_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_93_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21736_ _01296_ _01297_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27243_ clknet_3_7__leaf_clk_mosi _00857_ VGND VGND VPWR VPWR spi0.data_packed\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_24455_ _03809_ _03810_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21667_ _01205_ _01228_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_149_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23406_ net107 _02844_ _02845_ _02843_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__a22o_1
X_27174_ clknet_leaf_32_clk_sys _00788_ net618 VGND VGND VPWR VPWR top0.periodTop_r\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_20618_ _12142_ _12465_ VGND VGND VPWR VPWR _12467_ sky130_fd_sc_hd__nand2_1
X_24386_ _03741_ _03742_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__nor2_2
XFILLER_0_163_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21598_ _01146_ _01153_ _01159_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__a21o_2
X_26125_ spi0.data_packed\[20\] _05281_ _05282_ net918 VGND VGND VPWR VPWR _00801_
+ sky130_fd_sc_hd__a22o_1
X_23337_ _02755_ _02780_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20549_ _12279_ _12266_ _12397_ VGND VGND VPWR VPWR _12398_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14070_ net51 _05723_ _05724_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__and3_1
X_26056_ top0.pid_d.out\[6\] _05232_ _05233_ spi0.data_packed\[70\] VGND VGND VPWR
+ VPWR _05244_ sky130_fd_sc_hd__a22o_1
X_23268_ net1016 _02708_ _02716_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__o21ai_1
X_25007_ net1017 _04190_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22219_ _01223_ _01778_ _01779_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__o21ai_1
X_23199_ net260 net254 net251 net245 net204 net196 VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__mux4_1
X_17760_ _09718_ _09726_ _09737_ VGND VGND VPWR VPWR _09747_ sky130_fd_sc_hd__and3_1
X_14972_ _07041_ VGND VGND VPWR VPWR _07108_ sky130_fd_sc_hd__clkbuf_4
X_26958_ clknet_leaf_13_clk_sys _00575_ net616 VGND VGND VPWR VPWR top0.matmul0.b\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13923_ net65 _06135_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__and2_2
X_16711_ top0.pid_q.out\[14\] _08792_ _08795_ VGND VGND VPWR VPWR _08796_ sky130_fd_sc_hd__mux2_1
X_25909_ _05125_ _12014_ net844 _05029_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__a2bb2o_1
X_17691_ net398 net392 net345 net349 VGND VGND VPWR VPWR _09678_ sky130_fd_sc_hd__nand4_1
XFILLER_0_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26889_ clknet_leaf_37_clk_sys _00506_ net679 VGND VGND VPWR VPWR top0.svm0.tB\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16642_ _08692_ _08727_ VGND VGND VPWR VPWR _08728_ sky130_fd_sc_hd__xnor2_2
X_19430_ top0.pid_d.prev_int\[5\] _11325_ _11329_ VGND VGND VPWR VPWR _11330_ sky130_fd_sc_hd__o21ai_2
X_13854_ _06041_ _06038_ _06043_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16573_ _08629_ _08659_ VGND VGND VPWR VPWR _08660_ sky130_fd_sc_hd__xnor2_2
X_19361_ net722 _11273_ _11281_ _11269_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__a22o_1
X_13785_ _05996_ _05997_ net59 _05496_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18312_ _10168_ _10170_ _10169_ VGND VGND VPWR VPWR _10294_ sky130_fd_sc_hd__o21a_1
X_15524_ _07550_ _07551_ _07622_ VGND VGND VPWR VPWR _07623_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_128_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19292_ top0.pid_d.prev_error\[12\] top0.pid_d.curr_error\[12\] VGND VGND VPWR VPWR
+ _11234_ sky130_fd_sc_hd__and2_1
X_18243_ net416 net410 _09967_ top0.pid_d.mult0.b\[15\] _09567_ VGND VGND VPWR VPWR
+ _10226_ sky130_fd_sc_hd__a32o_1
XFILLER_0_72_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15455_ _07550_ _07553_ VGND VGND VPWR VPWR _07554_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_167_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14406_ _06581_ _06592_ _06613_ VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__a21oi_4
X_18174_ top0.pid_d.out\[3\] _09339_ _10157_ _10067_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15386_ net495 net491 VGND VGND VPWR VPWR _07485_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17125_ top0.pid_q.curr_int\[0\] top0.pid_q.prev_int\[0\] _09142_ VGND VGND VPWR
+ VPWR _09143_ sky130_fd_sc_hd__a21o_1
X_14337_ net855 _06280_ _06546_ _06381_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17056_ _09104_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__clkbuf_1
X_14268_ _06444_ _06445_ _06433_ _06434_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_21_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16007_ net449 net523 VGND VGND VPWR VPWR _08101_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13219_ _05443_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__clkbuf_2
X_14199_ _06313_ _06314_ VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17958_ net424 net313 VGND VGND VPWR VPWR _09944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16909_ net468 _08890_ _08969_ _08930_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17889_ _09798_ _09801_ VGND VGND VPWR VPWR _09876_ sky130_fd_sc_hd__nor2_1
X_19628_ _11484_ _11504_ _11509_ VGND VGND VPWR VPWR _11517_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19559_ _11447_ VGND VGND VPWR VPWR _11448_ sky130_fd_sc_hd__buf_2
XFILLER_0_94_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22570_ _02122_ _02123_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21521_ net131 _01078_ _01079_ _01082_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24240_ _03566_ _03596_ _03597_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__and3b_1
XFILLER_0_113_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21452_ net794 _12034_ _12037_ _01017_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__a31o_1
XFILLER_0_145_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20403_ _12249_ _12251_ VGND VGND VPWR VPWR _12252_ sky130_fd_sc_hd__and2b_1
XFILLER_0_181_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24171_ _03410_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__inv_2
X_21383_ _00933_ _00950_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23122_ top0.svm0.delta\[8\] _02615_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20334_ _12125_ _12150_ _12151_ _12166_ VGND VGND VPWR VPWR _12183_ sky130_fd_sc_hd__nand4_2
XFILLER_0_3_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23053_ net32 top0.svm0.counter\[13\] VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__xnor2_1
X_20265_ _12112_ _12105_ _12106_ VGND VGND VPWR VPWR _12114_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22004_ net106 _01565_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20196_ net262 net257 VGND VGND VPWR VPWR _12045_ sky130_fd_sc_hd__and2_1
X_26812_ clknet_leaf_51_clk_sys _00429_ net670 VGND VGND VPWR VPWR top0.pid_q.prev_int\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26743_ clknet_leaf_96_clk_sys _00360_ net588 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_23955_ _02998_ _03000_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__or2_2
X_22906_ top0.svm0.tC\[9\] _02422_ _02423_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__a21oi_1
X_26674_ clknet_leaf_81_clk_sys _00291_ net636 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_23886_ _02984_ _02986_ _03207_ _03208_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__o22a_1
XFILLER_0_169_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25625_ top0.matmul0.sin\[1\] top0.matmul0.sin\[0\] VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__nor2_1
X_22837_ _02354_ _02355_ _02356_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__or3b_1
XFILLER_0_168_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13570_ _05777_ _05782_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__xnor2_2
X_25556_ top0.matmul0.a\[1\] top0.matmul0.matmul_stage_inst.e\[1\] _04856_ VGND VGND
+ VPWR VPWR _04865_ sky130_fd_sc_hd__mux2_1
X_22768_ top0.pid_q.prev_int\[12\] _02291_ _02294_ top0.pid_q.curr_int\[12\] VGND
+ VGND VPWR VPWR _00431_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24507_ _03846_ _03847_ _03861_ _03652_ _03849_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_52_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21719_ net163 _01266_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__nor2_2
XFILLER_0_66_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25487_ _03148_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__buf_4
XFILLER_0_82_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22699_ _01948_ _02242_ _02243_ _02249_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15240_ net525 _07227_ _07338_ _07241_ VGND VGND VPWR VPWR _07339_ sky130_fd_sc_hd__a31o_1
X_27226_ clknet_3_4__leaf_clk_mosi _00840_ VGND VGND VPWR VPWR spi0.data_packed\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_24438_ _03790_ _03793_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15171_ _07268_ _07269_ VGND VGND VPWR VPWR _07270_ sky130_fd_sc_hd__xnor2_2
X_27157_ clknet_leaf_6_clk_sys _00771_ net596 VGND VGND VPWR VPWR top0.a_in_matmul\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_24369_ _03076_ _03077_ _03103_ _03104_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14122_ net27 _06333_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__and2_1
X_26108_ top0.periodTop\[7\] _05276_ _05278_ net47 VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27088_ clknet_leaf_1_clk_sys _00705_ net584 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14053_ _06260_ _06264_ _06265_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__o21ai_4
X_18930_ _10903_ _10904_ VGND VGND VPWR VPWR _10905_ sky130_fd_sc_hd__or2_2
X_26039_ net979 _05229_ _05230_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18861_ top0.pid_d.curr_int\[11\] _10836_ VGND VGND VPWR VPWR _10837_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_105_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17812_ net393 net388 net345 net349 VGND VGND VPWR VPWR _09799_ sky130_fd_sc_hd__nand4_1
XFILLER_0_100_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18792_ net377 _10690_ _10074_ _10767_ VGND VGND VPWR VPWR _10768_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17743_ _09418_ _09421_ VGND VGND VPWR VPWR _09730_ sky130_fd_sc_hd__nor2_1
X_14955_ _07099_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__clkbuf_1
X_13906_ _06102_ _06103_ _06118_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__a21oi_2
X_17674_ _09655_ _09660_ VGND VGND VPWR VPWR _09661_ sky130_fd_sc_hd__xnor2_1
X_14886_ spi0.data_packed\[51\] top0.kpq\[3\] _07053_ VGND VGND VPWR VPWR _07063_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19413_ top0.pid_d.prev_int\[3\] VGND VGND VPWR VPWR _11315_ sky130_fd_sc_hd__inv_2
X_16625_ _08637_ _08639_ _08710_ VGND VGND VPWR VPWR _08711_ sky130_fd_sc_hd__a21oi_2
X_13837_ _06023_ _06033_ _06030_ _06032_ _06039_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__o32a_1
XFILLER_0_98_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16556_ _08634_ _08642_ VGND VGND VPWR VPWR _08643_ sky130_fd_sc_hd__xnor2_2
X_19344_ top0.pid_d.curr_error\[3\] _11275_ _11278_ _11152_ VGND VGND VPWR VPWR _00297_
+ sky130_fd_sc_hd__a22o_1
X_13768_ _05973_ _05977_ _05980_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_114_Left_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15507_ _07253_ _07254_ _07604_ VGND VGND VPWR VPWR _07606_ sky130_fd_sc_hd__a21bo_1
X_16487_ net497 _08574_ VGND VGND VPWR VPWR _08575_ sky130_fd_sc_hd__nand2_1
X_19275_ _11216_ _11217_ VGND VGND VPWR VPWR _11219_ sky130_fd_sc_hd__or2_1
X_13699_ _05910_ _05911_ net59 _05517_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18226_ net319 _10206_ _10207_ _10208_ VGND VGND VPWR VPWR _10209_ sky130_fd_sc_hd__a22o_2
X_15438_ net480 _07274_ _07366_ VGND VGND VPWR VPWR _07537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18157_ _09593_ net307 _10140_ VGND VGND VPWR VPWR _10141_ sky130_fd_sc_hd__and3_1
X_15369_ net534 _07466_ _07467_ VGND VGND VPWR VPWR _07468_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17108_ net909 _09114_ _09130_ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__a21o_1
Xhold304 top0.b_in_matmul\[5\] VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__dlygate4sd3_1
X_18088_ _10053_ _10056_ _10054_ VGND VGND VPWR VPWR _10072_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17039_ _09073_ _09074_ _09075_ VGND VGND VPWR VPWR _09091_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_123_Left_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20050_ top0.cordic0.slte0.opA\[8\] _11784_ _11912_ VGND VGND VPWR VPWR _11914_ sky130_fd_sc_hd__or3_1
XFILLER_0_175_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23740_ _03092_ _03095_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_139_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20952_ _11788_ _12794_ _12798_ _12799_ VGND VGND VPWR VPWR _12800_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_132_Left_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23671_ net568 top0.matmul0.matmul_stage_inst.b\[11\] top0.matmul0.matmul_stage_inst.a\[11\]
+ net564 VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__a22o_4
XFILLER_0_67_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20883_ _12179_ _12242_ _12731_ VGND VGND VPWR VPWR _12732_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_89_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25410_ _04717_ _04753_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_178_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22622_ _02130_ _02127_ _02003_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__nand3b_1
X_26390_ clknet_leaf_39_clk_sys _00031_ net677 VGND VGND VPWR VPWR top0.svm0.tC\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_191_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25341_ _04614_ _04615_ _04613_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22553_ net102 _02103_ _02105_ _02107_ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__a31o_2
XFILLER_0_75_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21504_ net99 VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__clkinv_4
X_25272_ _04548_ _04549_ _04547_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_146_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22484_ _02038_ _02040_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__nor2_1
XFILLER_0_185_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27011_ clknet_leaf_23_clk_sys _00628_ net626 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_24223_ _03549_ _03580_ _03578_ _03575_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_185_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21435_ _01000_ _00995_ _00966_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24154_ _03483_ _03468_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_141_Left_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21366_ _11727_ _13001_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_169_Right_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23105_ _07117_ _02603_ VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__nor2_1
X_20317_ net214 _12165_ VGND VGND VPWR VPWR _12166_ sky130_fd_sc_hd__xnor2_2
X_24085_ _03328_ _03329_ _03332_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__and3_1
X_21297_ _13138_ _13139_ VGND VGND VPWR VPWR _13140_ sky130_fd_sc_hd__xnor2_2
X_23036_ net20 top0.svm0.counter\[15\] VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__or2_1
X_20248_ _12095_ _12096_ VGND VGND VPWR VPWR _12097_ sky130_fd_sc_hd__xnor2_2
X_20179_ _12009_ net208 _12026_ _12029_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__a31o_1
X_24987_ _03234_ _04174_ _03765_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14740_ _06939_ _06941_ VGND VGND VPWR VPWR _06943_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23938_ _03291_ _03270_ _03271_ _03287_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__or4_1
X_26726_ clknet_leaf_104_clk_sys _00343_ net576 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_150_Left_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14671_ _06841_ _06842_ VGND VGND VPWR VPWR _06875_ sky130_fd_sc_hd__nor2_1
X_26657_ clknet_leaf_78_clk_sys _00274_ net631 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_23869_ _03168_ _03169_ _03225_ _03226_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__o211ai_4
X_16410_ _08497_ _08498_ VGND VGND VPWR VPWR _08499_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13622_ _05574_ _05833_ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__or2_1
X_25608_ net725 _00000_ _04895_ VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__o21a_1
XFILLER_0_196_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17390_ net334 net338 VGND VGND VPWR VPWR _09377_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26588_ clknet_leaf_54_clk_sys _00211_ net669 VGND VGND VPWR VPWR top0.pid_q.prev_error\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16341_ net458 net503 VGND VGND VPWR VPWR _08431_ sky130_fd_sc_hd__nand2_1
X_13553_ net39 _05475_ _05476_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__and3_1
X_25539_ _05456_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19060_ top0.pid_d.out\[13\] top0.pid_d.curr_int\[13\] _11032_ VGND VGND VPWR VPWR
+ _11033_ sky130_fd_sc_hd__o21ai_2
X_16272_ _08261_ _08266_ _08259_ VGND VGND VPWR VPWR _08363_ sky130_fd_sc_hd__a21bo_1
X_13484_ _05541_ _05538_ _05539_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__nor3_1
XFILLER_0_192_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18011_ _09994_ _09995_ VGND VGND VPWR VPWR _09996_ sky130_fd_sc_hd__xnor2_1
X_15223_ _07313_ _07315_ VGND VGND VPWR VPWR _07322_ sky130_fd_sc_hd__nand2_1
X_27209_ clknet_leaf_6_clk_sys _00823_ net591 VGND VGND VPWR VPWR top0.cordic0.slte0.opB\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15154_ _07252_ _07210_ _07214_ VGND VGND VPWR VPWR _07253_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_63_clk_sys clknet_3_4__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_63_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_104_clk_sys clknet_3_0__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_104_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_14105_ _06310_ _06315_ _06316_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19962_ top0.cordic0.slte0.opA\[2\] _11785_ VGND VGND VPWR VPWR _11832_ sky130_fd_sc_hd__nor2_1
X_15085_ net540 net465 _07181_ _07177_ _07183_ VGND VGND VPWR VPWR _07184_ sky130_fd_sc_hd__a32o_1
XFILLER_0_200_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14036_ _06155_ _06247_ _06248_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__o21ai_2
X_18913_ _10804_ _10805_ _10722_ VGND VGND VPWR VPWR _10888_ sky130_fd_sc_hd__mux2_1
X_19893_ _11526_ _11767_ net175 VGND VGND VPWR VPWR _11768_ sky130_fd_sc_hd__o21ai_1
X_18844_ _10818_ _10819_ VGND VGND VPWR VPWR _10820_ sky130_fd_sc_hd__nor2_1
X_18775_ _10686_ _10750_ VGND VGND VPWR VPWR _10752_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15987_ top0.pid_q.out\[4\] _07700_ _08081_ _07710_ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17726_ _09698_ _09707_ _09712_ VGND VGND VPWR VPWR _09713_ sky130_fd_sc_hd__a21boi_1
X_14938_ _07090_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17657_ _09642_ _09624_ _09643_ VGND VGND VPWR VPWR _09644_ sky130_fd_sc_hd__a21o_1
XFILLER_0_187_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14869_ _07054_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16608_ _08312_ _08693_ VGND VGND VPWR VPWR _08694_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17588_ net342 net349 net425 _09525_ VGND VGND VPWR VPWR _09575_ sky130_fd_sc_hd__o22ai_1
X_19327_ _11258_ _11254_ _11255_ VGND VGND VPWR VPWR _11266_ sky130_fd_sc_hd__o21ba_1
X_16539_ _08624_ _08614_ _08625_ VGND VGND VPWR VPWR _08626_ sky130_fd_sc_hd__o21a_1
XFILLER_0_174_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19258_ top0.pid_d.curr_error\[8\] VGND VGND VPWR VPWR _11203_ sky130_fd_sc_hd__inv_2
X_18209_ _10115_ _10117_ _10191_ VGND VGND VPWR VPWR _10192_ sky130_fd_sc_hd__a21oi_2
X_19189_ top0.matmul0.alpha_pass\[0\] top0.matmul0.alpha_pass\[1\] top0.matmul0.alpha_pass\[2\]
+ VGND VGND VPWR VPWR _11141_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21220_ _12646_ _13054_ _13055_ _12577_ VGND VGND VPWR VPWR _13064_ sky130_fd_sc_hd__and4b_1
Xhold101 top0.c_out_calc\[8\] VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold112 top0.pid_q.prev_error\[8\] VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 top0.svm0.tB\[4\] VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 top0.svm0.tB\[6\] VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold145 top0.periodTop\[5\] VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__dlygate4sd3_1
X_21151_ _12971_ _12994_ VGND VGND VPWR VPWR _12996_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold156 top0.matmul0.matmul_stage_inst.b\[8\] VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 top0.c_out_calc\[6\] VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold178 top0.pid_d.prev_error\[4\] VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__dlygate4sd3_1
X_20102_ _11957_ _11960_ VGND VGND VPWR VPWR _11961_ sky130_fd_sc_hd__xor2_1
Xfanout603 net605 VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__clkbuf_4
X_21082_ _11788_ _12851_ net221 VGND VGND VPWR VPWR _12928_ sky130_fd_sc_hd__o21ai_1
Xhold189 top0.pid_d.prev_error\[9\] VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout614 net615 VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__buf_2
Xfanout625 net629 VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__clkbuf_4
X_24910_ _04258_ _04260_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__xnor2_2
Xfanout636 net638 VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__clkbuf_4
X_20033_ _11895_ _11897_ VGND VGND VPWR VPWR _11898_ sky130_fd_sc_hd__xor2_1
Xfanout647 net649 VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__clkbuf_4
X_25890_ _05106_ _05107_ _02282_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__a21o_1
Xfanout658 net661 VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__clkbuf_2
Xfanout669 net687 VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__buf_2
X_24841_ _04188_ _04192_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24772_ _04088_ _04124_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__xnor2_2
X_21984_ _01446_ _01428_ _01545_ _01450_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__a22oi_1
X_26511_ clknet_leaf_64_clk_sys _00134_ net656 VGND VGND VPWR VPWR top0.pid_q.out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_23723_ _03079_ _03080_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_179_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20935_ _12704_ _12706_ VGND VGND VPWR VPWR _12783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26442_ clknet_leaf_84_clk_sys _00083_ net640 VGND VGND VPWR VPWR top0.kid\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23654_ _02984_ _02986_ _02997_ _02999_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__o22a_1
X_20866_ net285 net259 VGND VGND VPWR VPWR _12715_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22605_ _02157_ _02158_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26373_ _05418_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23585_ _02959_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20797_ _12583_ _12605_ VGND VGND VPWR VPWR _12646_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25324_ _03280_ _03936_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22536_ _12036_ _02091_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25255_ _04596_ _04600_ _04595_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__a21o_1
X_22467_ _01643_ net92 _01119_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24206_ _03207_ _03208_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__nor2_2
XFILLER_0_122_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21418_ _00947_ _00948_ net219 VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__o21ai_1
X_25186_ _04404_ _04466_ _04468_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__a21o_1
X_22398_ _01918_ _01955_ _01259_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_103_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24137_ _03017_ _03114_ _03493_ _03494_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_32_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21349_ _13141_ _13146_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24068_ _03359_ _03362_ VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23019_ _02516_ _02520_ _02521_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_60_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15910_ net499 _07367_ _08002_ _08004_ net483 VGND VGND VPWR VPWR _08005_ sky130_fd_sc_hd__a32o_1
XFILLER_0_194_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16890_ top0.pid_q.prev_error\[5\] top0.pid_q.curr_error\[5\] VGND VGND VPWR VPWR
+ _08952_ sky130_fd_sc_hd__xor2_1
X_15841_ _07933_ _07936_ VGND VGND VPWR VPWR _07937_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18560_ net323 net376 VGND VGND VPWR VPWR _10539_ sky130_fd_sc_hd__nand2_1
X_15772_ _07738_ _07761_ _07868_ VGND VGND VPWR VPWR _07869_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17511_ net391 net385 VGND VGND VPWR VPWR _09498_ sky130_fd_sc_hd__nand2_1
X_14723_ _06924_ _06925_ VGND VGND VPWR VPWR _06926_ sky130_fd_sc_hd__xor2_2
XFILLER_0_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26709_ clknet_leaf_71_clk_sys _00326_ net657 VGND VGND VPWR VPWR top0.pid_d.curr_int\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_18491_ _10372_ _10374_ _10470_ VGND VGND VPWR VPWR _10471_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_3_7__f_clk_mosi clknet_0_clk_mosi VGND VGND VPWR VPWR clknet_3_7__leaf_clk_mosi
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_200_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14654_ _06819_ _06858_ VGND VGND VPWR VPWR _06859_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_184_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17442_ _09351_ net392 VGND VGND VPWR VPWR _09429_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13605_ _05816_ _05817_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14585_ _06751_ _06790_ VGND VGND VPWR VPWR _06791_ sky130_fd_sc_hd__xnor2_4
X_17373_ net395 net357 VGND VGND VPWR VPWR _09360_ sky130_fd_sc_hd__nand2_2
XFILLER_0_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19112_ _11082_ VGND VGND VPWR VPWR _11084_ sky130_fd_sc_hd__inv_2
X_13536_ _05742_ _05747_ _05748_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__and3_1
X_16324_ _08351_ _08353_ _08352_ VGND VGND VPWR VPWR _08414_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16255_ _08344_ _08345_ net497 VGND VGND VPWR VPWR _08346_ sky130_fd_sc_hd__or3b_2
X_19043_ _10950_ _10952_ _11015_ VGND VGND VPWR VPWR _11016_ sky130_fd_sc_hd__a21o_1
X_13467_ _05678_ _05679_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__xor2_1
XFILLER_0_180_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15206_ top0.pid_q.mult0.a\[2\] net475 VGND VGND VPWR VPWR _07305_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16186_ _08202_ _08203_ _08201_ VGND VGND VPWR VPWR _08278_ sky130_fd_sc_hd__o21ba_1
X_13398_ top0.matmul0.alpha_pass\[9\] _05435_ _05474_ VGND VGND VPWR VPWR _05611_
+ sky130_fd_sc_hd__nand3_4
XFILLER_0_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15137_ _07222_ _07235_ VGND VGND VPWR VPWR _07236_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19945_ _11806_ _11815_ _11426_ VGND VGND VPWR VPWR _11816_ sky130_fd_sc_hd__o21a_1
X_15068_ _07150_ _07151_ VGND VGND VPWR VPWR _07167_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14019_ _06229_ _06231_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__xnor2_1
X_19876_ _11732_ _11746_ _11748_ _11717_ _11751_ VGND VGND VPWR VPWR _11752_ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18827_ _10709_ _10714_ _10802_ VGND VGND VPWR VPWR _10803_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18758_ _10494_ _09771_ _10495_ VGND VGND VPWR VPWR _10735_ sky130_fd_sc_hd__and3_1
XFILLER_0_175_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17709_ _09493_ _09690_ _09694_ net352 _09695_ VGND VGND VPWR VPWR _09696_ sky130_fd_sc_hd__a221o_2
XFILLER_0_76_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18689_ _10666_ VGND VGND VPWR VPWR _10667_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20720_ net298 _12508_ _12567_ _12568_ VGND VGND VPWR VPWR _12569_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20651_ net249 _12499_ VGND VGND VPWR VPWR _12500_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23370_ _11518_ _02796_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20582_ _12201_ _12429_ _11550_ VGND VGND VPWR VPWR _12431_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22321_ _12036_ _01880_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25040_ _04387_ _04389_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22252_ net721 _12034_ _12037_ _01812_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21203_ net222 _12910_ VGND VGND VPWR VPWR _13047_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22183_ _01698_ _01720_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21134_ net251 _12917_ _12976_ _12977_ _12978_ VGND VGND VPWR VPWR _12979_ sky130_fd_sc_hd__a41o_1
X_26991_ clknet_leaf_26_clk_sys _00608_ net625 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout400 net401 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_4
Xfanout411 net414 VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__clkbuf_2
Xfanout422 net423 VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__clkbuf_4
X_25942_ _05145_ _05146_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__nand2_1
X_21065_ net230 _12072_ VGND VGND VPWR VPWR _12911_ sky130_fd_sc_hd__nand2_1
Xfanout433 net434 VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__buf_2
XFILLER_0_100_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout444 top0.pid_q.mult0.b\[15\] VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__buf_4
Xfanout455 net457 VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__buf_4
Xfanout466 net467 VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__clkbuf_4
Xfanout477 net478 VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__buf_2
X_20016_ top0.cordic0.slte0.opA\[5\] _11852_ _11868_ VGND VGND VPWR VPWR _11882_ sky130_fd_sc_hd__and3_1
X_25873_ _05083_ _05088_ _05089_ _05091_ _08900_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__a311o_1
Xfanout488 top0.pid_q.mult0.b\[2\] VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__buf_4
Xfanout499 top0.pid_q.mult0.a\[15\] VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__buf_4
X_24824_ _03017_ _03185_ _04175_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_198_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_11_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_11_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_3_clk_sys clknet_3_2__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_3_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_24755_ _03054_ _03055_ _03029_ _03030_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__o22a_1
XFILLER_0_69_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21967_ _01493_ _01514_ _01519_ _01528_ VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__o211a_1
X_23706_ net572 top0.matmul0.matmul_stage_inst.d\[1\] top0.matmul0.matmul_stage_inst.c\[1\]
+ net556 VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__a22o_4
X_20918_ _12764_ _12765_ net241 VGND VGND VPWR VPWR _12766_ sky130_fd_sc_hd__a21oi_1
X_24686_ _03910_ _03911_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__or2_1
X_21898_ _01081_ _01458_ net167 VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23637_ net565 net557 top0.matmul0.matmul_stage_inst.e\[6\] VGND VGND VPWR VPWR _02995_
+ sky130_fd_sc_hd__o21a_1
X_26425_ clknet_leaf_57_clk_sys _00066_ net644 VGND VGND VPWR VPWR top0.kpq\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_20849_ _12696_ _12697_ VGND VGND VPWR VPWR _12698_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout40 top0.periodTop_r\[10\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_4
Xfanout51 net1027 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_4
XFILLER_0_37_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout62 top0.periodTop_r\[1\] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_4
X_14370_ _06521_ _06577_ _06578_ VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__a21o_1
X_26356_ spi0.data_packed\[76\] spi0.data_packed\[77\] net690 VGND VGND VPWR VPWR
+ _05410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23568_ top0.b_in_matmul\[7\] top0.matmul0.b\[7\] _02948_ VGND VGND VPWR VPWR _02951_
+ sky130_fd_sc_hd__mux2_1
Xfanout73 net74 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_2
Xfanout84 net85 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_2
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout95 net96 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_2
X_25307_ _04651_ _04652_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__xnor2_1
X_13321_ _05533_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__buf_6
XFILLER_0_52_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22519_ _02074_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__inv_2
X_26287_ net957 VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__clkbuf_1
X_23499_ _02914_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16040_ _08132_ _08133_ VGND VGND VPWR VPWR _08134_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25238_ _04576_ _04584_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__xnor2_1
X_13252_ _05464_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__buf_4
XFILLER_0_162_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25169_ _04410_ _04516_ _04417_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_102_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17991_ _09893_ _09976_ VGND VGND VPWR VPWR _09977_ sky130_fd_sc_hd__xor2_2
XFILLER_0_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19730_ _11573_ net82 _11535_ _11613_ VGND VGND VPWR VPWR _11614_ sky130_fd_sc_hd__o22a_1
X_16942_ _08997_ _08998_ _08999_ VGND VGND VPWR VPWR _09000_ sky130_fd_sc_hd__and3_1
X_19661_ net1013 _11546_ _11525_ VGND VGND VPWR VPWR _11549_ sky130_fd_sc_hd__a21oi_1
X_16873_ top0.pid_q.curr_error\[3\] VGND VGND VPWR VPWR _08936_ sky130_fd_sc_hd__inv_2
X_18612_ net432 _10516_ _10517_ _10590_ net436 VGND VGND VPWR VPWR _10591_ sky130_fd_sc_hd__a32o_1
X_15824_ _07855_ _07857_ _07853_ VGND VGND VPWR VPWR _07920_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_126_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19592_ top0.cordic0.slte0.opA\[6\] top0.cordic0.slte0.opB\[6\] VGND VGND VPWR VPWR
+ _11481_ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18543_ net382 net317 VGND VGND VPWR VPWR _10522_ sky130_fd_sc_hd__nand2_1
X_15755_ _07850_ _07851_ VGND VGND VPWR VPWR _07852_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14706_ _06865_ _06903_ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__nand2_1
X_18474_ _10452_ _10453_ VGND VGND VPWR VPWR _10454_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15686_ net511 _07779_ _07780_ _07783_ VGND VGND VPWR VPWR _07784_ sky130_fd_sc_hd__a31o_1
XFILLER_0_184_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17425_ net329 net425 VGND VGND VPWR VPWR _09412_ sky130_fd_sc_hd__nand2_2
XFILLER_0_200_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14637_ net36 _05666_ VGND VGND VPWR VPWR _06842_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14568_ _06706_ _06711_ _06704_ VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_138_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17356_ _09340_ _09341_ _09342_ VGND VGND VPWR VPWR _09343_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16307_ _08316_ _08330_ _08396_ VGND VGND VPWR VPWR _08398_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13519_ _05536_ _05731_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14499_ _06623_ _06625_ _06705_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__o21a_1
X_17287_ _09282_ _09283_ VGND VGND VPWR VPWR _09284_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19026_ _10954_ _10997_ _10998_ _10845_ VGND VGND VPWR VPWR _10999_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_70_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16238_ _08326_ _08327_ VGND VGND VPWR VPWR _08329_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16169_ _08185_ _08187_ _08260_ VGND VGND VPWR VPWR _08261_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_11_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19928_ _11431_ _11799_ net177 VGND VGND VPWR VPWR _11800_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_177_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19859_ _11733_ _11735_ VGND VGND VPWR VPWR _11736_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22870_ _02324_ top0.svm0.tB\[6\] top0.svm0.tB\[5\] _02387_ _02388_ VGND VGND VPWR
+ VPWR _02389_ sky130_fd_sc_hd__a221o_1
XFILLER_0_183_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21821_ _01381_ _01382_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__and2_1
XFILLER_0_195_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24540_ _03892_ _03893_ _03890_ _03891_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__o211a_1
X_21752_ _01311_ _01313_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20703_ _12047_ _12551_ net305 VGND VGND VPWR VPWR _12552_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24471_ net556 top0.matmul0.matmul_stage_inst.c\[15\] top0.matmul0.matmul_stage_inst.b\[15\]
+ net568 VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__a22o_2
X_21683_ _01099_ _01243_ _01244_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__o21ai_2
X_26210_ spi0.data_packed\[3\] spi0.data_packed\[4\] net694 VGND VGND VPWR VPWR _05337_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23422_ net103 _02849_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__nor2_1
X_27190_ clknet_leaf_55_clk_sys _00804_ net668 VGND VGND VPWR VPWR top0.currT_r\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20634_ _12471_ _12482_ VGND VGND VPWR VPWR _12483_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26141_ spi0.data_packed\[0\] spi0.data_packed\[15\] net19 VGND VGND VPWR VPWR _05286_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23353_ net216 _02795_ _11560_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__mux2_2
XFILLER_0_184_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20565_ _12370_ _12412_ _12413_ VGND VGND VPWR VPWR _12414_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_34_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22304_ _01774_ _01792_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26072_ top0.pid_d.out\[10\] _05232_ _05233_ spi0.data_packed\[74\] VGND VGND VPWR
+ VPWR _05256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23284_ _02660_ _02669_ _02731_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__nor3_1
X_20496_ _11437_ _12059_ _12344_ VGND VGND VPWR VPWR _12345_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25023_ _04289_ _04291_ _04372_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22235_ _01748_ _01795_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22166_ _01724_ _01727_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__xnor2_1
X_21117_ _12742_ VGND VGND VPWR VPWR _12963_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26974_ clknet_leaf_28_clk_sys _00591_ net624 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[6\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout230 top0.cordic0.vec\[0\]\[14\] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_4
X_22097_ _01657_ _01658_ _01619_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__mux2_1
Xfanout241 net242 VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout252 top0.cordic0.vec\[0\]\[10\] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_6
X_25925_ top0.matmul0.alpha_pass\[13\] top0.matmul0.beta_pass\[13\] VGND VGND VPWR
+ VPWR _05140_ sky130_fd_sc_hd__xnor2_2
Xfanout263 net264 VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__buf_4
X_21048_ _12180_ _12893_ VGND VGND VPWR VPWR _12894_ sky130_fd_sc_hd__nor2_1
Xfanout274 net275 VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_4
Xfanout285 top0.cordic0.vec\[0\]\[4\] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__buf_4
Xfanout296 net297 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__clkbuf_4
X_13870_ _05801_ _05855_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__nor2_1
X_25856_ top0.matmul0.alpha_pass\[6\] _05074_ _05070_ VGND VGND VPWR VPWR _05077_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24807_ _04035_ _04032_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22999_ top0.svm0.delta\[11\] _02504_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25787_ _05018_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15540_ net462 net526 VGND VGND VPWR VPWR _07639_ sky130_fd_sc_hd__nand2_1
X_24738_ _03006_ _03198_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15471_ net531 net528 net462 net464 VGND VGND VPWR VPWR _07570_ sky130_fd_sc_hd__nand4_1
XFILLER_0_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24669_ _02989_ _02991_ _03093_ _03094_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__o22a_1
XFILLER_0_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14422_ _06567_ _06572_ VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__nor2_1
X_17210_ top0.pid_q.curr_int\[11\] top0.pid_q.prev_int\[11\] VGND VGND VPWR VPWR _09218_
+ sky130_fd_sc_hd__xnor2_1
X_26408_ clknet_leaf_79_clk_sys _00049_ net634 VGND VGND VPWR VPWR top0.kpd\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_18190_ _10106_ _10108_ _10107_ VGND VGND VPWR VPWR _10173_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14353_ net44 _05723_ _05724_ VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__and3_1
XFILLER_0_181_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17141_ _09154_ _09156_ VGND VGND VPWR VPWR _09157_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26339_ _05401_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__clkbuf_1
X_13304_ _05472_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17072_ _09110_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14284_ _06395_ _06396_ _06493_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__o21a_2
XFILLER_0_97_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16023_ _08027_ _08029_ _08116_ VGND VGND VPWR VPWR _08117_ sky130_fd_sc_hd__a21oi_2
X_13235_ _05453_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17974_ _09931_ _09959_ VGND VGND VPWR VPWR _09960_ sky130_fd_sc_hd__xnor2_2
X_19713_ _11596_ _11597_ _11576_ VGND VGND VPWR VPWR _11598_ sky130_fd_sc_hd__mux2_1
X_16925_ top0.currT_r\[7\] _08971_ _08983_ VGND VGND VPWR VPWR _08984_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19644_ net306 _11452_ _11424_ VGND VGND VPWR VPWR _11532_ sky130_fd_sc_hd__or3b_1
X_16856_ _08917_ _08919_ VGND VGND VPWR VPWR _08920_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_189_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15807_ _07901_ _07902_ VGND VGND VPWR VPWR _07903_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19575_ top0.cordic0.slte0.opB\[13\] top0.cordic0.slte0.opA\[13\] VGND VGND VPWR
+ VPWR _11464_ sky130_fd_sc_hd__xor2_1
XFILLER_0_177_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16787_ top0.kiq\[3\] _08863_ _08866_ VGND VGND VPWR VPWR _08867_ sky130_fd_sc_hd__and3_1
X_13999_ net27 net22 VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__nand2_4
XFILLER_0_34_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18526_ _10443_ _10505_ VGND VGND VPWR VPWR _10506_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15738_ net454 net528 VGND VGND VPWR VPWR _07835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18457_ _10400_ _10409_ _10399_ VGND VGND VPWR VPWR _10437_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15669_ _07617_ _07618_ _07766_ VGND VGND VPWR VPWR _07767_ sky130_fd_sc_hd__a21o_1
XFILLER_0_200_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17408_ _09394_ VGND VGND VPWR VPWR _09395_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18388_ _10365_ _10368_ VGND VGND VPWR VPWR _10369_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17339_ top0.matmul0.matmul_stage_inst.mult1\[13\] top0.matmul0.matmul_stage_inst.mult2\[13\]
+ VGND VGND VPWR VPWR _09328_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20350_ net247 net238 VGND VGND VPWR VPWR _12199_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19009_ _10892_ _10898_ _10897_ VGND VGND VPWR VPWR _10983_ sky130_fd_sc_hd__a21o_1
XFILLER_0_183_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20281_ _11437_ _12128_ _12129_ VGND VGND VPWR VPWR _12130_ sky130_fd_sc_hd__o21a_1
XFILLER_0_80_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_7__f_clk_sys clknet_0_clk_sys VGND VGND VPWR VPWR clknet_3_7__leaf_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_105_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22020_ _01310_ _01301_ _01496_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_12_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold16 top0.matmul0.matmul_stage_inst.a\[7\] VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold27 top0.cordic0.sin\[4\] VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__dlygate4sd3_1
X_23971_ _03312_ _03321_ _03327_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__nand3_2
Xhold38 top0.cordic0.cos\[6\] VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold49 top0.cordic0.sin\[2\] VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__dlygate4sd3_1
X_22922_ _02306_ _02437_ _02309_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25710_ net72 _04914_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__nand2_1
X_26690_ clknet_leaf_84_clk_sys _00307_ net641 VGND VGND VPWR VPWR top0.pid_d.curr_error\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_22853_ _02346_ _02372_ _02350_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__o21ba_1
X_25641_ net72 _04918_ _04890_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_196_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21804_ _01318_ _01365_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__nand2_1
X_25572_ _04873_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__clkbuf_1
X_22784_ _02297_ _02305_ _02307_ top0.svm0.out_valid VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24523_ _03872_ _03877_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__xnor2_2
X_21735_ _01290_ _01293_ _01295_ VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24454_ _03195_ _03198_ _03722_ _03324_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__o211a_1
X_27242_ clknet_3_7__leaf_clk_mosi _00856_ VGND VGND VPWR VPWR spi0.data_packed\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21666_ _01210_ _01227_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23405_ net108 _11857_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__nor2_1
XFILLER_0_188_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27173_ clknet_leaf_32_clk_sys _00787_ net618 VGND VGND VPWR VPWR top0.periodTop_r\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20617_ _12465_ VGND VGND VPWR VPWR _12466_ sky130_fd_sc_hd__inv_2
X_24385_ net556 top0.matmul0.matmul_stage_inst.c\[14\] top0.matmul0.matmul_stage_inst.b\[14\]
+ net568 VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__a22o_4
X_21597_ _01146_ _01153_ _01158_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26124_ _05277_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23336_ net128 _02774_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20548_ _12396_ _12363_ _12372_ VGND VGND VPWR VPWR _12397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26055_ _05243_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__clkbuf_1
X_23267_ _11425_ _02714_ _02715_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_18_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20479_ _12264_ _12327_ net280 VGND VGND VPWR VPWR _12328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25006_ _03280_ _03200_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22218_ net104 _01224_ net100 VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__mux2_1
X_23198_ net243 net237 net233 net228 net204 net196 VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__mux4_2
X_22149_ _01709_ _01710_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__xnor2_2
X_26957_ clknet_leaf_13_clk_sys _00574_ net616 VGND VGND VPWR VPWR top0.matmul0.b\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_14971_ _07107_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16710_ top0.pid_q.curr_int\[14\] _08794_ VGND VGND VPWR VPWR _08795_ sky130_fd_sc_hd__xnor2_1
X_13922_ top0.matmul0.alpha_pass\[15\] _05436_ _05717_ _06134_ VGND VGND VPWR VPWR
+ _06135_ sky130_fd_sc_hd__a31o_4
X_25908_ _05102_ _05112_ _05119_ _05120_ _05124_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__o221a_1
XFILLER_0_156_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17690_ net417 net332 _09675_ _09676_ VGND VGND VPWR VPWR _09677_ sky130_fd_sc_hd__a31o_1
XFILLER_0_195_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26888_ clknet_leaf_37_clk_sys _00505_ net679 VGND VGND VPWR VPWR top0.svm0.tB\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16641_ _08725_ _08726_ VGND VGND VPWR VPWR _08727_ sky130_fd_sc_hd__nand2_1
X_25839_ _05058_ _05061_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__xnor2_1
X_13853_ _06038_ _06044_ _06065_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_27_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19360_ _11121_ _11264_ _11278_ _11273_ net765 VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__a32o_1
X_16572_ _08653_ _08658_ VGND VGND VPWR VPWR _08659_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_201_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13784_ net54 _05484_ _05486_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__and3_1
X_18311_ _10186_ _10188_ _10292_ VGND VGND VPWR VPWR _10293_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15523_ _07550_ _07551_ _07552_ VGND VGND VPWR VPWR _07622_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19291_ top0.pid_d.mult0.b\[11\] _11094_ _11231_ _11233_ _08889_ VGND VGND VPWR VPWR
+ _00289_ sky130_fd_sc_hd__o221a_1
XFILLER_0_38_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18242_ _10088_ _10093_ _10092_ VGND VGND VPWR VPWR _10225_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_155_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15454_ _07551_ _07552_ VGND VGND VPWR VPWR _07553_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14405_ _06581_ _06592_ _06582_ VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_5_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18173_ net434 _10071_ _10156_ net439 _07138_ VGND VGND VPWR VPWR _10157_ sky130_fd_sc_hd__a221o_1
X_15385_ net539 VGND VGND VPWR VPWR _07484_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17124_ top0.pid_q.curr_int\[1\] top0.pid_q.prev_int\[1\] VGND VGND VPWR VPWR _09142_
+ sky130_fd_sc_hd__xor2_1
X_14336_ _06474_ _06545_ VGND VGND VPWR VPWR _06546_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_135_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14267_ _06433_ _06434_ _06444_ _06445_ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__o211a_1
X_17055_ net1018 _09103_ VGND VGND VPWR VPWR _09104_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16006_ net456 net1028 VGND VGND VPWR VPWR _08100_ sky130_fd_sc_hd__nand2_2
XFILLER_0_110_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13218_ _05442_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__buf_4
X_14198_ _06311_ _06312_ VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17957_ net420 net315 VGND VGND VPWR VPWR _09943_ sky130_fd_sc_hd__nand2_1
X_16908_ net546 _08962_ _08968_ _08882_ VGND VGND VPWR VPWR _08969_ sky130_fd_sc_hd__a211o_1
XFILLER_0_174_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17888_ _09798_ _09801_ VGND VGND VPWR VPWR _09875_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19627_ _11408_ _11515_ VGND VGND VPWR VPWR _11516_ sky130_fd_sc_hd__nand2_1
X_16839_ top0.matmul0.beta_pass\[2\] _08903_ VGND VGND VPWR VPWR _08904_ sky130_fd_sc_hd__xor2_1
XFILLER_0_189_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_58_clk_sys clknet_3_4__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_58_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_19558_ net182 net180 VGND VGND VPWR VPWR _11447_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18509_ _10487_ _10488_ VGND VGND VPWR VPWR _10489_ sky130_fd_sc_hd__xor2_1
XFILLER_0_158_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19489_ _11341_ _11375_ _11382_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__a21o_1
X_21520_ _01080_ net131 _01081_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__o21a_1
XFILLER_0_180_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21451_ _01015_ _01016_ _12740_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20402_ _12067_ _12250_ VGND VGND VPWR VPWR _12251_ sky130_fd_sc_hd__xnor2_2
X_24170_ _03410_ _03526_ _03527_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__mux2_1
X_21382_ _00947_ _00949_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23121_ top0.svm0.delta\[7\] _02612_ _02595_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__o21a_1
X_20333_ _12150_ _12151_ _12177_ _12125_ VGND VGND VPWR VPWR _12182_ sky130_fd_sc_hd__a211o_1
XFILLER_0_189_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23052_ _05500_ _02551_ _02552_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20264_ _12105_ _12106_ _12112_ VGND VGND VPWR VPWR _12113_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22003_ net124 net109 VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__nand2_1
X_20195_ net253 _12042_ _12043_ VGND VGND VPWR VPWR _12044_ sky130_fd_sc_hd__a21boi_1
X_26811_ clknet_leaf_69_clk_sys _00428_ net663 VGND VGND VPWR VPWR top0.pid_q.prev_int\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26742_ clknet_leaf_96_clk_sys _00359_ net587 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_23954_ _03308_ _03311_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22905_ top0.svm0.tC\[9\] _02422_ _02360_ VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__o21a_1
X_23885_ _03004_ _03005_ _02976_ _02977_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__o22a_1
X_26673_ clknet_leaf_81_clk_sys _00290_ net636 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22836_ _02352_ top0.svm0.tA\[1\] VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25624_ _04890_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_196_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25555_ _04864_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__clkbuf_1
X_22767_ net914 _02291_ _02294_ top0.pid_q.curr_int\[11\] VGND VGND VPWR VPWR _00430_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24506_ _03846_ _03858_ _03654_ _03657_ VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__o211a_1
X_21718_ net147 net142 VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__nor2_1
X_25486_ _04828_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22698_ net104 _02244_ _02245_ _01063_ _02248_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27225_ clknet_3_5__leaf_clk_mosi _00839_ VGND VGND VPWR VPWR spi0.data_packed\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_191_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24437_ _03791_ _03792_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21649_ net105 VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_118_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15170_ net526 net470 VGND VGND VPWR VPWR _07269_ sky130_fd_sc_hd__nand2_1
X_24368_ _03060_ _03123_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27156_ clknet_leaf_10_clk_sys _00770_ net594 VGND VGND VPWR VPWR top0.a_in_matmul\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14121_ _05523_ _05524_ _05489_ _05491_ VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__a22o_1
X_26107_ top0.periodTop\[6\] _05276_ _05278_ net50 VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__a22o_1
X_23319_ _02755_ _02764_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__xnor2_1
X_27087_ clknet_leaf_2_clk_sys _00704_ net610 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_24299_ _03624_ _03625_ _03622_ _03620_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14052_ _06263_ _06133_ _06136_ _06130_ _06085_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__o2111ai_4
X_26038_ _05164_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18860_ _10834_ _10758_ _10835_ VGND VGND VPWR VPWR _10836_ sky130_fd_sc_hd__a21o_1
XFILLER_0_197_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17811_ _09658_ _09796_ _09797_ VGND VGND VPWR VPWR _09798_ sky130_fd_sc_hd__a21oi_2
X_18791_ _09356_ _09758_ VGND VGND VPWR VPWR _10767_ sky130_fd_sc_hd__nor2_1
X_17742_ _09505_ _09728_ _09506_ VGND VGND VPWR VPWR _09729_ sky130_fd_sc_hd__mux2_1
X_14954_ spi0.data_packed\[19\] top0.kiq\[3\] _07097_ VGND VGND VPWR VPWR _07099_
+ sky130_fd_sc_hd__mux2_1
X_13905_ _06109_ _06117_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__xnor2_4
X_17673_ _09656_ _09659_ VGND VGND VPWR VPWR _09660_ sky130_fd_sc_hd__xnor2_2
X_14885_ _07062_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19412_ top0.pid_d.curr_int\[3\] _11290_ _11293_ _11314_ VGND VGND VPWR VPWR _00329_
+ sky130_fd_sc_hd__a22o_1
X_16624_ _08637_ _08639_ _08638_ VGND VGND VPWR VPWR _08710_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_100_clk_sys clknet_3_0__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_100_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_13836_ _05567_ _06032_ _06033_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19343_ net986 _11275_ _11278_ _11142_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16555_ _08636_ _08641_ VGND VGND VPWR VPWR _08642_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13767_ _05973_ _05977_ _05979_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_168_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15506_ _07255_ _07600_ _07602_ _07604_ VGND VGND VPWR VPWR _07605_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_31_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19274_ _11216_ _11217_ VGND VGND VPWR VPWR _11218_ sky130_fd_sc_hd__nand2_1
X_16486_ net458 net461 net466 VGND VGND VPWR VPWR _08574_ sky130_fd_sc_hd__or3_1
X_13698_ net54 _05478_ _05479_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18225_ net356 net360 net365 VGND VGND VPWR VPWR _10208_ sky130_fd_sc_hd__o21ai_4
X_15437_ net514 net480 VGND VGND VPWR VPWR _07536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18156_ net416 net315 _10138_ _10139_ VGND VGND VPWR VPWR _10140_ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15368_ net534 net484 _07456_ net537 VGND VGND VPWR VPWR _07467_ sky130_fd_sc_hd__and4b_1
XFILLER_0_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17107_ top0.pid_q.curr_error\[12\] _08860_ _09116_ VGND VGND VPWR VPWR _09130_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14319_ _06513_ _06528_ VGND VGND VPWR VPWR _06529_ sky130_fd_sc_hd__xor2_2
XFILLER_0_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold305 top0.cordic0.sin\[6\] VGND VGND VPWR VPWR net1005 sky130_fd_sc_hd__dlygate4sd3_1
X_18087_ _10069_ _10070_ VGND VGND VPWR VPWR _10071_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15299_ _07380_ _07381_ _07392_ _07396_ VGND VGND VPWR VPWR _07398_ sky130_fd_sc_hd__and4_1
XFILLER_0_111_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17038_ _09087_ _09089_ VGND VGND VPWR VPWR _09090_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18989_ _10861_ _10873_ _10962_ VGND VGND VPWR VPWR _10963_ sky130_fd_sc_hd__o21a_1
XFILLER_0_197_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20951_ _12795_ _12792_ VGND VGND VPWR VPWR _12799_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23670_ net565 net557 top0.matmul0.matmul_stage_inst.e\[1\] VGND VGND VPWR VPWR _03028_
+ sky130_fd_sc_hd__o21a_4
XFILLER_0_49_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20882_ _12161_ _12192_ _12194_ VGND VGND VPWR VPWR _12731_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_191_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22621_ _02138_ _02174_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__xor2_2
XFILLER_0_88_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25340_ _04619_ _04624_ _04684_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22552_ _01069_ _01616_ _02106_ _01643_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21503_ net116 VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__inv_2
X_25271_ _04613_ _04616_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_5_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22483_ _01925_ _02039_ net80 VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27010_ clknet_leaf_23_clk_sys _00627_ net625 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_24222_ _03572_ _03324_ _03579_ _03542_ _03323_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__a32o_1
XFILLER_0_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21434_ _00998_ _00999_ _00987_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24153_ _03490_ _03498_ _03510_ VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21365_ _13169_ _13179_ _13180_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23104_ top0.svm0.delta\[3\] _02602_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20316_ net239 net230 VGND VGND VPWR VPWR _12165_ sky130_fd_sc_hd__nand2_2
X_24084_ _03438_ _03441_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21296_ _13001_ _12990_ VGND VGND VPWR VPWR _13139_ sky130_fd_sc_hd__or2_1
X_23035_ net21 top0.svm0.counter\[15\] VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__nand2_1
X_20247_ net240 net230 VGND VGND VPWR VPWR _12096_ sky130_fd_sc_hd__xnor2_4
X_20178_ _12026_ _12028_ _12009_ VGND VGND VPWR VPWR _12029_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24986_ _04257_ _04260_ _04335_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__o21ai_4
X_26725_ clknet_leaf_103_clk_sys _00342_ net576 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_23937_ _03291_ _03293_ _03294_ _03287_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__and4_1
XFILLER_0_99_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_6__f_clk_mosi clknet_0_clk_mosi VGND VGND VPWR VPWR clknet_3_6__leaf_clk_mosi
+ sky130_fd_sc_hd__clkbuf_16
X_14670_ _06841_ _06842_ VGND VGND VPWR VPWR _06874_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26656_ clknet_leaf_79_clk_sys _00273_ net632 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_23868_ _03193_ _03194_ _03224_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__nand3_4
XFILLER_0_196_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13621_ _05574_ _05833_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__nand2_1
X_25607_ _04886_ top0.matmul0.cos\[7\] _04878_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__or3_1
X_22819_ top0.svm0.counter\[3\] VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__inv_2
X_26587_ clknet_leaf_54_clk_sys _00210_ net667 VGND VGND VPWR VPWR top0.pid_q.prev_error\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_23799_ _03155_ _03156_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__nand2_2
XFILLER_0_95_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16340_ net466 net497 VGND VGND VPWR VPWR _08430_ sky130_fd_sc_hd__nand2_2
X_13552_ net37 _05478_ _05479_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__and3_1
X_25538_ _04855_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13483_ net45 _05585_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__nand2_1
X_16271_ _08350_ _08361_ VGND VGND VPWR VPWR _08362_ sky130_fd_sc_hd__xnor2_2
X_25469_ _04809_ _04811_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__nor2_1
X_18010_ net416 net315 VGND VGND VPWR VPWR _09995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15222_ _07313_ _07315_ VGND VGND VPWR VPWR _07321_ sky130_fd_sc_hd__nor2_2
X_27208_ clknet_leaf_93_clk_sys _00822_ net600 VGND VGND VPWR VPWR top0.cordic0.slte0.opB\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27139_ clknet_leaf_13_clk_sys _00753_ net616 VGND VGND VPWR VPWR top0.b_in_matmul\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15153_ _07211_ _07212_ VGND VGND VPWR VPWR _07252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14104_ _06313_ _06314_ _06311_ _06312_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__o211ai_1
X_19961_ _11431_ _11830_ net177 VGND VGND VPWR VPWR _11831_ sky130_fd_sc_hd__o21ai_1
X_15084_ net460 net464 _07178_ _07182_ VGND VGND VPWR VPWR _07183_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_10_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14035_ _06157_ _06159_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__or2b_1
X_18912_ _10880_ _10886_ VGND VGND VPWR VPWR _10887_ sky130_fd_sc_hd__xnor2_1
X_19892_ _11764_ _11766_ VGND VGND VPWR VPWR _11767_ sky130_fd_sc_hd__xnor2_1
X_18843_ _10816_ _10817_ VGND VGND VPWR VPWR _10819_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18774_ _10686_ _10750_ VGND VGND VPWR VPWR _10751_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15986_ net548 _08075_ _08080_ net545 _07705_ VGND VGND VPWR VPWR _08081_ sky130_fd_sc_hd__a221o_1
X_17725_ net382 net357 _09708_ _09711_ net352 VGND VGND VPWR VPWR _09712_ sky130_fd_sc_hd__a32o_1
XFILLER_0_145_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14937_ spi0.data_packed\[43\] top0.kid\[11\] _07086_ VGND VGND VPWR VPWR _07090_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17656_ _09627_ _09630_ VGND VGND VPWR VPWR _09643_ sky130_fd_sc_hd__nor2_1
X_14868_ spi0.data_packed\[74\] top0.kpd\[10\] _07053_ VGND VGND VPWR VPWR _07054_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16607_ _08534_ _08657_ _08526_ VGND VGND VPWR VPWR _08693_ sky130_fd_sc_hd__a21oi_1
X_13819_ _05735_ _05501_ _06031_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__or3b_1
X_17587_ net354 _09571_ _09573_ VGND VGND VPWR VPWR _09574_ sky130_fd_sc_hd__a21oi_1
X_14799_ _06989_ _06999_ VGND VGND VPWR VPWR _07000_ sky130_fd_sc_hd__xor2_2
XFILLER_0_86_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19326_ _10311_ _11125_ _11261_ _11265_ _05430_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__a221oi_2
X_16538_ _08624_ _08614_ top0.pid_q.out\[11\] VGND VGND VPWR VPWR _08625_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_85_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19257_ net329 _11117_ _11200_ _11202_ _08889_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__o221a_1
X_16469_ _08555_ _08556_ VGND VGND VPWR VPWR _08557_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18208_ _10115_ _10117_ _10116_ VGND VGND VPWR VPWR _10191_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19188_ top0.matmul0.alpha_pass\[0\] top0.matmul0.alpha_pass\[1\] top0.matmul0.alpha_pass\[2\]
+ VGND VGND VPWR VPWR _11140_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18139_ _10016_ _10018_ _10122_ VGND VGND VPWR VPWR _10123_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_5_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold102 top0.currT_r\[15\] VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 top0.matmul0.matmul_stage_inst.b\[12\] VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 top0.svm0.tC\[14\] VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold135 top0.svm0.tB\[2\] VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__dlygate4sd3_1
X_21150_ _12971_ _12994_ VGND VGND VPWR VPWR _12995_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold146 top0.matmul0.matmul_stage_inst.d\[1\] VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 top0.svm0.tC\[11\] VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 top0.svm0.tC\[12\] VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__dlygate4sd3_1
X_20101_ _11942_ _11950_ _11958_ _11959_ VGND VGND VPWR VPWR _11960_ sky130_fd_sc_hd__o31a_1
XFILLER_0_106_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold179 top0.pid_d.prev_error\[6\] VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__dlygate4sd3_1
X_21081_ _12180_ _12923_ _12925_ _12926_ _11739_ VGND VGND VPWR VPWR _12927_ sky130_fd_sc_hd__a221o_1
Xfanout604 net605 VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__buf_2
XFILLER_0_81_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout615 net629 VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__buf_2
Xfanout626 net629 VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__buf_2
XFILLER_0_0_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20032_ _11880_ _11886_ _11896_ VGND VGND VPWR VPWR _11897_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_176_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout637 net638 VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__clkbuf_4
Xfanout648 net649 VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout659 net660 VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__clkbuf_4
X_24840_ _04189_ _04191_ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24771_ _04089_ _04123_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__xnor2_1
X_21983_ _01544_ _01429_ _01446_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26510_ clknet_leaf_66_clk_sys _00133_ net660 VGND VGND VPWR VPWR top0.pid_q.out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_23722_ _03069_ _03071_ _03057_ _03058_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__o22a_1
X_20934_ _12760_ _12781_ VGND VGND VPWR VPWR _12782_ sky130_fd_sc_hd__xnor2_2
X_26441_ clknet_leaf_80_clk_sys _00082_ net640 VGND VGND VPWR VPWR top0.kid\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_23653_ _02993_ _02995_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__or2_1
X_20865_ _12101_ _12713_ net291 VGND VGND VPWR VPWR _12714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22604_ net79 _01115_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__xnor2_1
X_23584_ top0.b_in_matmul\[15\] net943 _05460_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__mux2_1
X_26372_ spi0.opcode\[4\] spi0.opcode\[5\] net691 VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__mux2_1
X_20796_ _12620_ _12638_ _12618_ VGND VGND VPWR VPWR _12645_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25323_ _04639_ _04638_ _04667_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22535_ _02083_ _02090_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_187_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25254_ _04595_ _04596_ _04600_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22466_ _01852_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24205_ _03560_ _03561_ _03562_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__a21o_1
X_21417_ _00968_ _00983_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__xnor2_1
X_25185_ _04474_ _04532_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__xor2_1
X_22397_ net119 _01917_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24136_ _03491_ _03492_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21348_ _13188_ _00916_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__or2b_1
X_24067_ _03424_ _03371_ _03335_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21279_ net242 _11727_ VGND VGND VPWR VPWR _13122_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23018_ top0.svm0.counter\[13\] top0.svm0.delta\[13\] VGND VGND VPWR VPWR _02521_
+ sky130_fd_sc_hd__nand2_1
X_15840_ _07934_ _07935_ VGND VGND VPWR VPWR _07936_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_200_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15771_ _07738_ _07761_ _07656_ VGND VGND VPWR VPWR _07868_ sky130_fd_sc_hd__o21ba_1
X_24969_ _04316_ _04319_ _04170_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17510_ _09352_ net395 _09355_ VGND VGND VPWR VPWR _09497_ sky130_fd_sc_hd__a21oi_1
X_14722_ net20 _05626_ _06833_ VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__and3_1
X_26708_ clknet_leaf_84_clk_sys net723 net645 VGND VGND VPWR VPWR top0.pid_d.prev_error\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_18490_ _10372_ _10374_ _10373_ VGND VGND VPWR VPWR _10470_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17441_ net392 net357 VGND VGND VPWR VPWR _09428_ sky130_fd_sc_hd__nand2_1
X_14653_ _06852_ _06857_ VGND VGND VPWR VPWR _06858_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_196_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26639_ clknet_leaf_81_clk_sys _00256_ net638 VGND VGND VPWR VPWR top0.pid_d.out\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_200_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13604_ net50 _05523_ _05524_ VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__and3_1
X_17372_ net400 net353 VGND VGND VPWR VPWR _09359_ sky130_fd_sc_hd__nand2_1
X_14584_ _06758_ _06789_ VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_82_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19111_ top0.pid_d.out\[14\] top0.pid_d.curr_int\[14\] _11082_ VGND VGND VPWR VPWR
+ _11083_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16323_ _08377_ _08379_ _08412_ VGND VGND VPWR VPWR _08413_ sky130_fd_sc_hd__a21o_1
X_13535_ _05743_ _05744_ _05745_ _05746_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__nand4bb_2
XFILLER_0_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19042_ _10950_ _10952_ _10848_ VGND VGND VPWR VPWR _11015_ sky130_fd_sc_hd__o21a_1
X_16254_ _08340_ _08343_ _08048_ VGND VGND VPWR VPWR _08345_ sky130_fd_sc_hd__a21oi_1
X_13466_ net39 _05523_ _05524_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15205_ _07166_ _07303_ VGND VGND VPWR VPWR _07304_ sky130_fd_sc_hd__xnor2_4
X_16185_ _08192_ _08194_ _08276_ VGND VGND VPWR VPWR _08277_ sky130_fd_sc_hd__a21oi_2
X_13397_ _05607_ _05608_ _05609_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__or3_2
XFILLER_0_2_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15136_ _07226_ _07234_ VGND VGND VPWR VPWR _07235_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19944_ _11809_ _11814_ net189 VGND VGND VPWR VPWR _11815_ sky130_fd_sc_hd__o21a_1
X_15067_ _07162_ _07165_ VGND VGND VPWR VPWR _07166_ sky130_fd_sc_hd__xnor2_4
X_14018_ _06113_ _06114_ _06230_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__o21a_1
X_19875_ net243 _11749_ _11750_ _11720_ VGND VGND VPWR VPWR _11751_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_65_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18826_ _10709_ _10714_ _10633_ VGND VGND VPWR VPWR _10802_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18757_ _09771_ _10495_ _10494_ VGND VGND VPWR VPWR _10734_ sky130_fd_sc_hd__a21oi_1
X_15969_ _07964_ _07976_ _07977_ VGND VGND VPWR VPWR _08064_ sky130_fd_sc_hd__o21a_1
X_17708_ net352 _09459_ _09687_ VGND VGND VPWR VPWR _09695_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18688_ _10657_ _10665_ VGND VGND VPWR VPWR _10666_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17639_ net403 net344 net348 net398 VGND VGND VPWR VPWR _09626_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20650_ _12498_ VGND VGND VPWR VPWR _12499_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19309_ top0.pid_d.prev_error\[13\] top0.pid_d.curr_error\[13\] VGND VGND VPWR VPWR
+ _11250_ sky130_fd_sc_hd__xor2_1
XFILLER_0_74_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20581_ net275 _12429_ _12274_ VGND VGND VPWR VPWR _12430_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22320_ _01814_ _01879_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22251_ _12036_ _01811_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21202_ _12911_ _12910_ _11759_ VGND VGND VPWR VPWR _13046_ sky130_fd_sc_hd__a21o_1
XFILLER_0_182_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22182_ _01698_ _01720_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__nor2_1
X_21133_ _12917_ _12972_ VGND VGND VPWR VPWR _12978_ sky130_fd_sc_hd__and2b_1
XFILLER_0_197_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26990_ clknet_leaf_25_clk_sys _00607_ net627 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout401 net402 VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout412 net413 VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__clkbuf_4
X_25941_ _05439_ _05150_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__nand2_1
X_21064_ net235 _12207_ _12703_ _12909_ VGND VGND VPWR VPWR _12910_ sky130_fd_sc_hd__a211o_2
Xfanout423 net424 VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__clkbuf_4
Xfanout434 top0.pid_d.state\[4\] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__clkbuf_4
Xfanout445 net446 VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__clkbuf_4
Xfanout456 net457 VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__clkbuf_4
X_20015_ _11852_ _11865_ _11868_ VGND VGND VPWR VPWR _11881_ sky130_fd_sc_hd__and3_1
Xfanout467 top0.pid_q.mult0.b\[7\] VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__buf_2
X_25872_ _05088_ _05090_ _05089_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__nor3_1
Xfanout478 top0.pid_q.mult0.b\[4\] VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__buf_2
Xfanout489 net492 VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__buf_2
X_24823_ _03157_ _03572_ _03315_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__a21oi_1
X_24754_ _03018_ _03019_ _03069_ _03071_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__o22a_1
XFILLER_0_96_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21966_ _01523_ _01527_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23705_ net568 top0.matmul0.matmul_stage_inst.b\[1\] top0.matmul0.matmul_stage_inst.a\[1\]
+ net564 VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__a22o_4
XFILLER_0_139_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20917_ net232 net228 VGND VGND VPWR VPWR _12765_ sky130_fd_sc_hd__nand2_1
X_24685_ _03908_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21897_ net160 _01458_ net155 VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26424_ clknet_leaf_56_clk_sys _00065_ net664 VGND VGND VPWR VPWR top0.kpq\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_23636_ _02993_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__buf_2
X_20848_ net213 net225 VGND VGND VPWR VPWR _12697_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_83_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout30 net31 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_4
Xfanout41 top0.periodTop_r\[9\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_194_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout52 net1027 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_153_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout63 net64 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_4
X_26355_ _05409_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__clkbuf_1
X_23567_ _02950_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__clkbuf_1
Xfanout74 top0.matmul0.op\[0\] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_2
X_20779_ _12622_ _12627_ _12626_ VGND VGND VPWR VPWR _12628_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout85 top0.cordic0.vec\[1\]\[17\] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
X_25306_ _04382_ _04580_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__nand2_1
X_13320_ _05531_ _05532_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__or2_1
Xfanout96 net97 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_2
X_22518_ _02071_ _02072_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__nor2_1
X_26286_ spi0.data_packed\[41\] net956 net688 VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__mux2_1
X_23498_ net1002 top0.matmul0.cos\[4\] _02904_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25237_ _04582_ _04583_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__and2b_1
X_13251_ _05463_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22449_ _01895_ _01943_ _01988_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25168_ _03007_ _04039_ _04067_ _03305_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__or4b_4
X_24119_ _03456_ _03471_ _03476_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25099_ _04436_ _04447_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__xnor2_1
X_17990_ _09902_ _09975_ VGND VGND VPWR VPWR _09976_ sky130_fd_sc_hd__xnor2_2
X_16941_ top0.currT_r\[9\] _08899_ top0.matmul0.beta_pass\[9\] VGND VGND VPWR VPWR
+ _08999_ sky130_fd_sc_hd__or3b_1
XFILLER_0_198_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19660_ _11434_ VGND VGND VPWR VPWR _11548_ sky130_fd_sc_hd__clkbuf_2
X_16872_ top0.currT_r\[4\] _08934_ VGND VGND VPWR VPWR _08935_ sky130_fd_sc_hd__xnor2_2
X_18611_ _10579_ _10589_ VGND VGND VPWR VPWR _10590_ sky130_fd_sc_hd__xnor2_1
X_15823_ _07910_ _07918_ VGND VGND VPWR VPWR _07919_ sky130_fd_sc_hd__xnor2_4
X_19591_ top0.cordic0.slte0.opB\[9\] top0.cordic0.slte0.opA\[9\] VGND VGND VPWR VPWR
+ _11480_ sky130_fd_sc_hd__xor2_1
X_18542_ net382 net367 _10520_ _09689_ _09364_ VGND VGND VPWR VPWR _10521_ sky130_fd_sc_hd__a32o_1
X_15754_ net461 net521 VGND VGND VPWR VPWR _07851_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14705_ _06861_ _06905_ VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18473_ net401 net309 VGND VGND VPWR VPWR _10453_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15685_ _07663_ _07782_ _07667_ VGND VGND VPWR VPWR _07783_ sky130_fd_sc_hd__a21oi_1
X_17424_ _09407_ _09410_ VGND VGND VPWR VPWR _09411_ sky130_fd_sc_hd__xnor2_4
X_14636_ net34 _05619_ VGND VGND VPWR VPWR _06841_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17355_ net415 net348 VGND VGND VPWR VPWR _09342_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14567_ _06764_ _06772_ VGND VGND VPWR VPWR _06773_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_144_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16306_ _08316_ _08330_ _08396_ VGND VGND VPWR VPWR _08397_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13518_ _05611_ _05612_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__nand2_4
X_17286_ top0.matmul0.matmul_stage_inst.mult1\[6\] top0.matmul0.matmul_stage_inst.mult2\[6\]
+ VGND VGND VPWR VPWR _09283_ sky130_fd_sc_hd__xor2_1
X_14498_ _06623_ _06625_ _06624_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__a21bo_1
X_19025_ _10954_ _10955_ _10957_ VGND VGND VPWR VPWR _10998_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16237_ _08326_ _08327_ VGND VGND VPWR VPWR _08328_ sky130_fd_sc_hd__nand2_1
X_13449_ top0.matmul0.beta_pass\[13\] VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16168_ _08185_ _08187_ _08186_ VGND VGND VPWR VPWR _08260_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15119_ _07215_ _07216_ _07210_ VGND VGND VPWR VPWR _07218_ sky130_fd_sc_hd__a21o_1
X_16099_ net456 net516 VGND VGND VPWR VPWR _08192_ sky130_fd_sc_hd__nand2_2
X_19927_ _11796_ _11798_ net181 VGND VGND VPWR VPWR _11799_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_167_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19858_ _11713_ _11721_ _11734_ VGND VGND VPWR VPWR _11735_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_183_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18809_ _10772_ _10784_ VGND VGND VPWR VPWR _10785_ sky130_fd_sc_hd__xnor2_2
X_19789_ net260 _11435_ _11669_ VGND VGND VPWR VPWR _11671_ sky130_fd_sc_hd__and3_1
X_21820_ _01123_ _01380_ net152 VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__o21bai_1
X_21751_ _01090_ _01312_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20702_ net289 net278 VGND VGND VPWR VPWR _12551_ sky130_fd_sc_hd__xor2_2
XFILLER_0_149_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24470_ _03825_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__clkbuf_4
X_21682_ _01110_ _01128_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20633_ _12469_ _12470_ _12481_ VGND VGND VPWR VPWR _12482_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_58_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23421_ net103 _02849_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23352_ _02663_ _02664_ _11654_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26140_ _05285_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__clkbuf_1
X_20564_ _12370_ _12412_ _12387_ VGND VGND VPWR VPWR _12413_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22303_ _01776_ _01862_ net77 VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23283_ _11425_ _02714_ _02715_ _02692_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__a211o_1
X_26071_ _05255_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__clkbuf_1
X_20495_ net282 net288 VGND VGND VPWR VPWR _12344_ sky130_fd_sc_hd__and2b_1
XFILLER_0_132_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25022_ _04289_ _04291_ _04371_ _03758_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__o211a_1
X_22234_ _01793_ _01794_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22165_ net86 _01232_ _01725_ _01726_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__o211a_1
X_21116_ _12952_ _12961_ VGND VGND VPWR VPWR _12962_ sky130_fd_sc_hd__xnor2_2
X_26973_ clknet_leaf_28_clk_sys _00590_ net622 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_22096_ _01628_ _01632_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout220 top0.cordic0.vec\[0\]\[17\] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_2
Xfanout231 net232 VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__buf_2
Xfanout242 net243 VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__buf_2
X_25924_ top0.matmul0.alpha_pass\[12\] top0.matmul0.beta_pass\[12\] VGND VGND VPWR
+ VPWR _05139_ sky130_fd_sc_hd__or2_1
Xfanout253 net256 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_4
X_21047_ _11758_ _12820_ VGND VGND VPWR VPWR _12893_ sky130_fd_sc_hd__nor2_1
Xfanout264 net268 VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__buf_4
Xfanout275 net279 VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__buf_4
Xfanout286 top0.cordic0.vec\[0\]\[4\] VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__buf_2
XFILLER_0_198_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout297 top0.cordic0.vec\[0\]\[2\] VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkbuf_4
X_25855_ _05070_ _05073_ _05075_ _02282_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__a211o_1
XFILLER_0_119_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24806_ _04064_ _04156_ _04157_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25786_ _05012_ top0.matmul0.start _05017_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__mux2_1
X_22998_ top0.svm0.delta\[10\] _02499_ _02503_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_55_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24737_ _03114_ _03826_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21949_ net156 _01441_ _01494_ _01500_ _01510_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__o311a_1
XFILLER_0_55_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15470_ _07565_ _07568_ VGND VGND VPWR VPWR _07569_ sky130_fd_sc_hd__xnor2_1
X_24668_ _02998_ _03000_ _03090_ _03091_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__o22a_2
XFILLER_0_37_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14421_ _06619_ _06628_ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__xnor2_4
X_26407_ clknet_leaf_79_clk_sys _00048_ net632 VGND VGND VPWR VPWR top0.kpd\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_23619_ net564 net557 top0.matmul0.matmul_stage_inst.e\[4\] VGND VGND VPWR VPWR _02977_
+ sky130_fd_sc_hd__o21a_4
XFILLER_0_182_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24599_ _03948_ _03953_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17140_ _09153_ _09147_ _09148_ _09155_ VGND VGND VPWR VPWR _09156_ sky130_fd_sc_hd__a31o_1
X_14352_ net48 _06131_ VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__nand2_2
X_26338_ spi0.data_packed\[67\] spi0.data_packed\[68\] net692 VGND VGND VPWR VPWR
+ _05401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13303_ _05513_ _05514_ _05515_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__o21a_1
X_17071_ net1018 _09109_ VGND VGND VPWR VPWR _09110_ sky130_fd_sc_hd__and2_1
X_14283_ net45 _05625_ _06395_ _06396_ VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26269_ _05366_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16022_ _08027_ _08029_ _08028_ VGND VGND VPWR VPWR _08116_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13234_ net543 _05442_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17973_ _09957_ _09958_ VGND VGND VPWR VPWR _09959_ sky130_fd_sc_hd__or2b_1
X_16924_ top0.currT_r\[7\] _08971_ _08972_ VGND VGND VPWR VPWR _08983_ sky130_fd_sc_hd__o21a_1
X_19712_ net188 _11441_ VGND VGND VPWR VPWR _11597_ sky130_fd_sc_hd__nand2_1
X_16855_ top0.currT_r\[3\] _08918_ VGND VGND VPWR VPWR _08919_ sky130_fd_sc_hd__xnor2_1
X_19643_ _11424_ _11527_ _11530_ VGND VGND VPWR VPWR _11531_ sky130_fd_sc_hd__a21oi_1
X_15806_ top0.pid_q.out\[3\] top0.pid_q.curr_int\[3\] VGND VGND VPWR VPWR _07902_
+ sky130_fd_sc_hd__xor2_1
X_19574_ top0.cordic0.slte0.opB\[3\] _11457_ _11458_ _11462_ VGND VGND VPWR VPWR _11463_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_172_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16786_ _08854_ VGND VGND VPWR VPWR _08866_ sky130_fd_sc_hd__clkbuf_2
X_13998_ _06210_ _05493_ _05494_ _05490_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__or4b_1
XFILLER_0_149_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18525_ _10504_ VGND VGND VPWR VPWR _10505_ sky130_fd_sc_hd__inv_2
X_15737_ net451 net532 VGND VGND VPWR VPWR _07834_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18456_ _10406_ _10407_ _10435_ VGND VGND VPWR VPWR _10436_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_34_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15668_ _07617_ _07618_ _07619_ VGND VGND VPWR VPWR _07766_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17407_ net357 VGND VGND VPWR VPWR _09394_ sky130_fd_sc_hd__inv_2
X_14619_ _06351_ VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__buf_6
XFILLER_0_157_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18387_ _10366_ _10367_ VGND VGND VPWR VPWR _10368_ sky130_fd_sc_hd__xor2_1
XFILLER_0_157_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15599_ net553 net543 VGND VGND VPWR VPWR _07698_ sky130_fd_sc_hd__or2_2
XFILLER_0_16_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17338_ top0.matmul0.matmul_stage_inst.mult1\[13\] top0.matmul0.matmul_stage_inst.mult2\[13\]
+ VGND VGND VPWR VPWR _09327_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17269_ _09268_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19008_ _10930_ _10981_ VGND VGND VPWR VPWR _10982_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20280_ net299 net283 net276 VGND VGND VPWR VPWR _12129_ sky130_fd_sc_hd__or3b_1
XFILLER_0_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_54_clk_sys clknet_3_6__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_54_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_51_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold17 top0.matmul0.matmul_stage_inst.a\[4\] VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold28 top0.pid_q.prev_error\[14\] VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__dlygate4sd3_1
X_23970_ _03312_ _03321_ _03327_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__a21o_1
Xhold39 top0.matmul0.matmul_stage_inst.d\[8\] VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__dlygate4sd3_1
X_22921_ top0.svm0.delta\[1\] _02436_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__xor2_1
X_25640_ net69 top0.matmul0.sin\[3\] VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22852_ _02371_ _02343_ _02342_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21803_ _01335_ _01348_ _01353_ _01363_ _01364_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__a311o_1
X_25571_ top0.matmul0.a\[8\] top0.matmul0.matmul_stage_inst.e\[8\] _04867_ VGND VGND
+ VPWR VPWR _04873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22783_ net171 _02306_ _02305_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24522_ _03873_ _03876_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_137_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21734_ _01290_ _01293_ _01295_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27241_ clknet_3_7__leaf_clk_mosi _00855_ VGND VGND VPWR VPWR spi0.data_packed\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_24453_ _03807_ _03808_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__xnor2_2
X_21665_ _01220_ _01226_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23404_ net1014 _02843_ net178 VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__o21ai_1
X_27172_ clknet_leaf_12_clk_sys _00786_ net618 VGND VGND VPWR VPWR top0.periodTop_r\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_20616_ net275 net263 VGND VGND VPWR VPWR _12465_ sky130_fd_sc_hd__xor2_2
X_24384_ net573 net564 top0.matmul0.matmul_stage_inst.a\[14\] VGND VGND VPWR VPWR
+ _03741_ sky130_fd_sc_hd__o21a_4
X_21596_ _01154_ _01157_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26123_ _05275_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20547_ _12390_ _12276_ _12280_ VGND VGND VPWR VPWR _12396_ sky130_fd_sc_hd__mux2_1
X_23335_ _01135_ net1013 _02777_ _02779_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26054_ top0.a_in_matmul\[5\] _05242_ _05230_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20478_ net300 net297 VGND VGND VPWR VPWR _12327_ sky130_fd_sc_hd__xnor2_1
X_23266_ net180 _02289_ net215 VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25005_ _03343_ _04097_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__nor2_2
X_22217_ _01213_ net100 VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__nor2_1
X_23197_ _05719_ _07038_ _02648_ net839 VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22148_ _01144_ _01456_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__xnor2_1
X_26956_ clknet_leaf_13_clk_sys _00573_ net616 VGND VGND VPWR VPWR top0.matmul0.b\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14970_ spi0.data_packed\[27\] top0.kiq\[11\] _07097_ VGND VGND VPWR VPWR _07107_
+ sky130_fd_sc_hd__mux2_1
X_22079_ _01621_ _01622_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13921_ top0.matmul0.beta_pass\[15\] _05436_ _05719_ _05465_ top0.c_out_calc\[15\]
+ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__a32o_1
X_25907_ _05122_ _05123_ top0.matmul0.alpha_pass\[10\] _02282_ VGND VGND VPWR VPWR
+ _05124_ sky130_fd_sc_hd__a211o_1
XFILLER_0_96_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26887_ clknet_leaf_38_clk_sys _00504_ net677 VGND VGND VPWR VPWR top0.svm0.tB\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16640_ _08694_ _08724_ VGND VGND VPWR VPWR _08726_ sky130_fd_sc_hd__or2_1
X_25838_ _05059_ _05060_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__xnor2_1
X_13852_ _06045_ _06048_ _06061_ _06064_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16571_ _08527_ _08657_ VGND VGND VPWR VPWR _08658_ sky130_fd_sc_hd__xor2_2
XFILLER_0_198_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13783_ net58 _05489_ _05491_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__and3_1
X_25769_ _05005_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18310_ _10186_ _10188_ _10187_ VGND VGND VPWR VPWR _10292_ sky130_fd_sc_hd__o21a_1
X_15522_ _07617_ _07620_ VGND VGND VPWR VPWR _07621_ sky130_fd_sc_hd__xnor2_2
X_19290_ _11121_ _11232_ _11123_ VGND VGND VPWR VPWR _11233_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18241_ _10095_ _10223_ _10129_ VGND VGND VPWR VPWR _10224_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15453_ net522 net470 VGND VGND VPWR VPWR _07552_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14404_ net869 _06280_ _06612_ _06381_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18172_ _10064_ _10155_ VGND VGND VPWR VPWR _10156_ sky130_fd_sc_hd__xnor2_1
X_15384_ net534 net487 VGND VGND VPWR VPWR _07483_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17123_ _09136_ _09139_ _09141_ top0.pid_q.curr_int\[0\] VGND VGND VPWR VPWR _00213_
+ sky130_fd_sc_hd__a22o_1
X_14335_ _06543_ _06544_ VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__nor2_4
XFILLER_0_52_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17054_ _08907_ top0.pid_q.curr_error\[2\] _09096_ VGND VGND VPWR VPWR _09103_ sky130_fd_sc_hd__mux2_1
X_14266_ _06464_ _06467_ _06475_ VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__o21a_1
X_16005_ _08020_ _08022_ _08098_ VGND VGND VPWR VPWR _08099_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13217_ _05441_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14197_ _06398_ _06407_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_148_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17956_ net426 net310 VGND VGND VPWR VPWR _09942_ sky130_fd_sc_hd__nand2_2
XFILLER_0_100_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16907_ _08967_ net550 VGND VGND VPWR VPWR _08968_ sky130_fd_sc_hd__and2b_1
X_17887_ _09866_ _09873_ VGND VGND VPWR VPWR _09874_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_174_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19626_ _11514_ VGND VGND VPWR VPWR _11515_ sky130_fd_sc_hd__clkbuf_4
X_16838_ _08891_ _08901_ _08902_ VGND VGND VPWR VPWR _08903_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_189_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16769_ _00011_ _07700_ _08842_ _08852_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__a31o_1
X_19557_ net138 net133 net129 net125 net197 net191 VGND VGND VPWR VPWR _11446_ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18508_ _10380_ _10392_ _10391_ VGND VGND VPWR VPWR _10488_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19488_ top0.pid_d.curr_int\[12\] _11289_ _11292_ _11381_ VGND VGND VPWR VPWR _11382_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_180_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18439_ _10323_ _10418_ _10419_ VGND VGND VPWR VPWR _10420_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21450_ net1021 _00994_ _01014_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_111_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20401_ net261 net249 VGND VGND VPWR VPWR _12250_ sky130_fd_sc_hd__xnor2_2
X_21381_ _11789_ _00948_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23120_ net933 _02613_ _02614_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__a21o_1
X_20332_ _12180_ _12073_ VGND VGND VPWR VPWR _12181_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23051_ net34 top0.svm0.counter\[12\] _02550_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__or3_1
X_20263_ _12068_ _12107_ _12110_ _12111_ VGND VGND VPWR VPWR _12112_ sky130_fd_sc_hd__o211a_1
X_22002_ net118 net102 VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__nand2_1
X_20194_ net258 net253 VGND VGND VPWR VPWR _12043_ sky130_fd_sc_hd__or2_1
X_26810_ clknet_leaf_68_clk_sys _00427_ net663 VGND VGND VPWR VPWR top0.pid_q.prev_int\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_26741_ clknet_leaf_96_clk_sys _00358_ net587 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_23953_ _03309_ _03310_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__xnor2_4
X_22904_ _02367_ top0.svm0.tC\[8\] _02421_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__a21o_1
X_26672_ clknet_leaf_82_clk_sys _00289_ net646 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_3_5__f_clk_mosi clknet_0_clk_mosi VGND VGND VPWR VPWR clknet_3_5__leaf_clk_mosi
+ sky130_fd_sc_hd__clkbuf_16
X_23884_ _03238_ _03241_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__xnor2_4
X_25623_ _04903_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__clkbuf_1
X_22835_ _02298_ top0.svm0.tA\[0\] VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25554_ top0.matmul0.a\[0\] top0.matmul0.matmul_stage_inst.e\[0\] _04856_ VGND VGND
+ VPWR VPWR _04864_ sky130_fd_sc_hd__mux2_1
X_22766_ net988 _02291_ _02294_ top0.pid_q.curr_int\[10\] VGND VGND VPWR VPWR _00429_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24505_ _03751_ _03846_ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21717_ _01262_ _01264_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__nor2_1
X_25485_ top0.matmul0.matmul_stage_inst.mult2\[15\] _04827_ _03146_ VGND VGND VPWR
+ VPWR _04828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22697_ net104 _02247_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27224_ clknet_3_4__leaf_clk_mosi _00838_ VGND VGND VPWR VPWR spi0.data_packed\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_24436_ _02979_ _02980_ _03054_ _03055_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__o22a_1
XFILLER_0_191_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21648_ _01207_ _01209_ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_136_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27155_ clknet_leaf_6_clk_sys _00769_ net594 VGND VGND VPWR VPWR top0.a_in_matmul\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_24367_ _03721_ _03723_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__nor2_1
X_21579_ _01137_ _01138_ _01140_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__or3_2
X_14120_ net22 _05497_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__nand2_1
X_26106_ net845 _05276_ _05278_ net1027 VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23318_ _02756_ _02762_ _02763_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__or3_2
XFILLER_0_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27086_ clknet_leaf_8_clk_sys _00703_ net584 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_24298_ _03624_ _03625_ _03622_ _03630_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14051_ _06263_ _06133_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__nand2_1
X_26037_ top0.matmul0.alpha_pass\[2\] _05203_ _05228_ VGND VGND VPWR VPWR _05229_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_162_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23249_ _02697_ _02698_ net156 VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17810_ net409 net335 net337 net404 VGND VGND VPWR VPWR _09797_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_24_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18790_ _10731_ _10741_ _10765_ VGND VGND VPWR VPWR _10766_ sky130_fd_sc_hd__o21ai_4
X_17741_ _09418_ _09421_ VGND VGND VPWR VPWR _09728_ sky130_fd_sc_hd__xnor2_1
X_26939_ clknet_leaf_8_clk_sys _00556_ net595 VGND VGND VPWR VPWR top0.matmul0.a\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14953_ _07098_ VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__clkbuf_1
X_13904_ _06111_ _06116_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__xor2_2
X_17672_ _09657_ _09658_ VGND VGND VPWR VPWR _09659_ sky130_fd_sc_hd__xnor2_1
X_14884_ spi0.data_packed\[50\] top0.kpq\[2\] _07053_ VGND VGND VPWR VPWR _07062_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16623_ _08636_ _08641_ _08708_ VGND VGND VPWR VPWR _08709_ sky130_fd_sc_hd__o21a_1
X_19411_ net431 _10156_ _11313_ net442 _11149_ VGND VGND VPWR VPWR _11314_ sky130_fd_sc_hd__a221o_1
X_13835_ net68 net62 _06023_ _06047_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__and4_1
XFILLER_0_187_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16554_ _08637_ _08640_ VGND VGND VPWR VPWR _08641_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19342_ top0.pid_d.curr_error\[1\] _11275_ _11278_ _11131_ VGND VGND VPWR VPWR _00295_
+ sky130_fd_sc_hd__a22o_1
X_13766_ _05960_ _05978_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15505_ _07226_ _07249_ _07597_ _07603_ VGND VGND VPWR VPWR _07604_ sky130_fd_sc_hd__or4_2
X_19273_ top0.pid_d.prev_error\[10\] top0.pid_d.curr_error\[10\] VGND VGND VPWR VPWR
+ _11217_ sky130_fd_sc_hd__xnor2_1
X_16485_ net466 _08141_ _08572_ VGND VGND VPWR VPWR _08573_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13697_ net57 _05475_ _05476_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18224_ net401 net319 VGND VGND VPWR VPWR _10207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15436_ net494 net489 net508 VGND VGND VPWR VPWR _07535_ sky130_fd_sc_hd__and3_1
XFILLER_0_183_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18155_ _09993_ _09994_ VGND VGND VPWR VPWR _10139_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15367_ _07228_ _07456_ net537 _07227_ VGND VGND VPWR VPWR _07466_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_142_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17106_ net898 _09114_ _09129_ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14318_ _06516_ _06527_ VGND VGND VPWR VPWR _06528_ sky130_fd_sc_hd__xor2_2
X_18086_ top0.pid_d.out\[3\] top0.pid_d.curr_int\[3\] VGND VGND VPWR VPWR _10070_
+ sky130_fd_sc_hd__xnor2_1
X_15298_ _07380_ _07381_ _07392_ _07396_ VGND VGND VPWR VPWR _07397_ sky130_fd_sc_hd__a22o_1
Xhold306 top0.periodTop\[15\] VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17037_ top0.currT_r\[15\] _09088_ VGND VGND VPWR VPWR _09089_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14249_ _06450_ _06451_ _06458_ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__nand3_1
XFILLER_0_123_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18988_ _10861_ _10873_ _10848_ VGND VGND VPWR VPWR _10962_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_183_Right_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17939_ _09844_ _09845_ _09924_ VGND VGND VPWR VPWR _09925_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_178_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20950_ _12795_ _12796_ _12797_ _12791_ net213 VGND VGND VPWR VPWR _12798_ sky130_fd_sc_hd__a311o_1
XFILLER_0_108_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19609_ top0.cordic0.slte0.opA\[13\] _11465_ VGND VGND VPWR VPWR _11498_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20881_ _12677_ _12729_ VGND VGND VPWR VPWR _12730_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22620_ _02172_ _02173_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22551_ _01069_ _01616_ _02102_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__a21o_1
XFILLER_0_192_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_46_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21502_ net110 net93 VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__nand2_2
X_25270_ _04614_ _04615_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22482_ _01924_ _01923_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__nor2_1
X_24221_ _03017_ _03323_ _03217_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21433_ _00916_ _00927_ _00956_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24152_ _03490_ _03498_ _03509_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21364_ _13130_ _00930_ _00931_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_47_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23103_ top0.svm0.delta\[1\] net555 top0.svm0.delta\[2\] _02595_ VGND VGND VPWR VPWR
+ _02602_ sky130_fd_sc_hd__o31a_1
X_20315_ _12072_ _12073_ VGND VGND VPWR VPWR _12164_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24083_ _03439_ _03440_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21295_ _13040_ _13042_ _13137_ VGND VGND VPWR VPWR _13138_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23034_ _02522_ _02528_ _02529_ _02535_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__o211ai_1
X_20246_ net244 _12094_ VGND VGND VPWR VPWR _12095_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_12_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_55_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20177_ net209 net206 VGND VGND VPWR VPWR _12028_ sky130_fd_sc_hd__or2_1
X_24985_ _04257_ _04260_ _04258_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26724_ clknet_leaf_78_clk_sys _00341_ net633 VGND VGND VPWR VPWR top0.pid_d.curr_int\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23936_ _03269_ _03266_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26655_ clknet_leaf_81_clk_sys _00272_ net633 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_23867_ _03193_ _03194_ _03224_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__a21o_2
XFILLER_0_54_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13620_ _05571_ _05572_ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__xnor2_1
X_25606_ net755 _00000_ _04887_ _04894_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__o22a_1
X_22818_ _02334_ _02335_ _02336_ _02337_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__a22o_1
X_26586_ clknet_leaf_54_clk_sys _00209_ net667 VGND VGND VPWR VPWR top0.pid_q.prev_error\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_23798_ net565 net557 top0.matmul0.matmul_stage_inst.e\[2\] VGND VGND VPWR VPWR _03156_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_94_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_64_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13551_ net42 _05472_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__nand2_1
X_25537_ top0.matmul0.b\[8\] top0.matmul0.matmul_stage_inst.f\[8\] _04846_ VGND VGND
+ VPWR VPWR _04855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22749_ _11997_ _02289_ _02290_ net180 VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16270_ _08355_ _08360_ VGND VGND VPWR VPWR _08361_ sky130_fd_sc_hd__xnor2_1
X_25468_ _04808_ _04750_ _04721_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__o21a_1
XFILLER_0_165_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13482_ _05499_ _05507_ _05694_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15221_ net527 VGND VGND VPWR VPWR _07320_ sky130_fd_sc_hd__inv_2
X_27207_ clknet_leaf_93_clk_sys _00821_ net600 VGND VGND VPWR VPWR top0.cordic0.slte0.opB\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_24419_ _03686_ _03692_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25399_ _03326_ _04687_ _04371_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27138_ clknet_leaf_12_clk_sys _00752_ net616 VGND VGND VPWR VPWR top0.b_in_matmul\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_15152_ net480 _07248_ _07250_ VGND VGND VPWR VPWR _07251_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_133_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14103_ _06311_ _06312_ _06313_ _06314_ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27069_ clknet_leaf_2_clk_sys _00686_ net584 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.c\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_19960_ _11822_ _11829_ VGND VGND VPWR VPWR _11830_ sky130_fd_sc_hd__xor2_1
X_15083_ net541 VGND VGND VPWR VPWR _07182_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_73_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14034_ _06159_ _06157_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__and2b_1
X_18911_ _10885_ _10884_ _10633_ VGND VGND VPWR VPWR _10886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19891_ _11742_ _11753_ _11765_ VGND VGND VPWR VPWR _11766_ sky130_fd_sc_hd__a21o_1
X_18842_ _10816_ _10817_ VGND VGND VPWR VPWR _10818_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18773_ _10743_ _10749_ VGND VGND VPWR VPWR _10750_ sky130_fd_sc_hd__xnor2_1
X_15985_ _08078_ _08079_ VGND VGND VPWR VPWR _08080_ sky130_fd_sc_hd__xnor2_1
X_17724_ net385 _09709_ _09710_ net391 VGND VGND VPWR VPWR _09711_ sky130_fd_sc_hd__a22o_1
X_14936_ _07089_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17655_ _09627_ _09630_ VGND VGND VPWR VPWR _09642_ sky130_fd_sc_hd__nand2_1
X_14867_ _07041_ VGND VGND VPWR VPWR _07053_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_82_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16606_ _08653_ _08658_ _08691_ VGND VGND VPWR VPWR _08692_ sky130_fd_sc_hd__a21oi_2
X_13818_ net59 _05488_ _05490_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17586_ _09356_ _09572_ net360 net410 VGND VGND VPWR VPWR _09573_ sky130_fd_sc_hd__o211a_1
X_14798_ _06947_ _06991_ _06996_ _06935_ _06998_ VGND VGND VPWR VPWR _06999_ sky130_fd_sc_hd__o221a_1
XFILLER_0_175_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19325_ _11121_ _11264_ _11123_ VGND VGND VPWR VPWR _11265_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16537_ top0.pid_q.curr_int\[11\] VGND VGND VPWR VPWR _08624_ sky130_fd_sc_hd__inv_2
X_13749_ net58 _05478_ _05479_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16468_ net450 net506 VGND VGND VPWR VPWR _08556_ sky130_fd_sc_hd__nand2_1
X_19256_ _11121_ _11201_ _11125_ VGND VGND VPWR VPWR _11202_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18207_ _10186_ _10189_ VGND VGND VPWR VPWR _10190_ sky130_fd_sc_hd__xnor2_1
X_15419_ _07430_ _07454_ _07516_ _07517_ VGND VGND VPWR VPWR _07518_ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19187_ net439 _11137_ _11138_ VGND VGND VPWR VPWR _11139_ sky130_fd_sc_hd__and3_1
X_16399_ _08483_ _08486_ VGND VGND VPWR VPWR _08488_ sky130_fd_sc_hd__or2_1
XFILLER_0_170_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18138_ _10016_ _10018_ _10017_ VGND VGND VPWR VPWR _10122_ sky130_fd_sc_hd__o21a_1
XFILLER_0_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold103 top0.kpq\[14\] VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_91_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold114 top0.svm0.tB\[8\] VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold125 top0.matmul0.matmul_stage_inst.c\[11\] VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__dlygate4sd3_1
X_18069_ _09964_ _09968_ VGND VGND VPWR VPWR _10054_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold136 top0.matmul0.matmul_stage_inst.d\[5\] VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 top0.matmul0.matmul_stage_inst.c\[3\] VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold158 top0.svm0.tC\[15\] VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__dlygate4sd3_1
X_20100_ top0.cordic0.slte0.opA\[12\] _11949_ VGND VGND VPWR VPWR _11959_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold169 top0.svm0.tC\[4\] VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__dlygate4sd3_1
X_21080_ _12072_ _11788_ VGND VGND VPWR VPWR _12926_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout605 net606 VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout616 net620 VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__clkbuf_4
X_20031_ _11879_ _11883_ _11885_ top0.cordic0.slte0.opA\[6\] VGND VGND VPWR VPWR _11896_
+ sky130_fd_sc_hd__o31ai_1
Xfanout627 net628 VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout638 net639 VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__clkbuf_4
Xfanout649 net654 VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24770_ _04104_ _04122_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__xnor2_2
X_21982_ _01428_ _01429_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__nor2_1
X_23721_ _03036_ _03037_ _03054_ _03055_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__o22a_1
X_20933_ _12775_ _12780_ VGND VGND VPWR VPWR _12781_ sky130_fd_sc_hd__xor2_1
XFILLER_0_152_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26440_ clknet_leaf_80_clk_sys _00081_ net633 VGND VGND VPWR VPWR top0.kid\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_23652_ _03004_ _03005_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__or2_2
XFILLER_0_117_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20864_ net265 net271 VGND VGND VPWR VPWR _12713_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22603_ _02155_ _02156_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__nand2_1
X_26371_ _05417_ VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__clkbuf_1
X_23583_ _02958_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20795_ _12618_ _12620_ _12638_ _12643_ VGND VGND VPWR VPWR _12644_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25322_ _04639_ _04638_ _04665_ _04666_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__o22a_1
XFILLER_0_187_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22534_ _02003_ _02007_ _02084_ _02089_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25253_ _04406_ _04599_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22465_ _02019_ _02021_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24204_ _03315_ _03337_ _03323_ _03217_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__and4_1
X_21416_ _00945_ _00982_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__xor2_1
X_25184_ _04525_ _04531_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_162_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22396_ top0.cordic0.vec\[1\]\[10\] _01917_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__nor2_1
X_24135_ _03491_ _03492_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21347_ _13157_ _13187_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__nand2_2
XFILLER_0_60_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24066_ _03350_ VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__inv_2
X_21278_ net262 _13116_ _13120_ VGND VGND VPWR VPWR _13121_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_60_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23017_ top0.svm0.counter\[13\] top0.svm0.delta\[13\] VGND VGND VPWR VPWR _02520_
+ sky130_fd_sc_hd__nor2_1
X_20229_ _12076_ _12077_ VGND VGND VPWR VPWR _12078_ sky130_fd_sc_hd__or2b_1
XFILLER_0_21_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15770_ _07832_ _07866_ VGND VGND VPWR VPWR _07867_ sky130_fd_sc_hd__xor2_2
X_24968_ _04235_ _04317_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__nand2_1
X_14721_ _06920_ _06923_ VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_169_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23919_ _03239_ _03240_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__and2_1
X_26707_ clknet_leaf_85_clk_sys net766 net641 VGND VGND VPWR VPWR top0.pid_d.prev_error\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24899_ _04157_ _04247_ _04248_ _04249_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_58_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17440_ _09413_ _09426_ VGND VGND VPWR VPWR _09427_ sky130_fd_sc_hd__xnor2_4
X_14652_ _06854_ _06856_ VGND VGND VPWR VPWR _06857_ sky130_fd_sc_hd__xor2_1
XFILLER_0_170_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26638_ clknet_leaf_80_clk_sys _00255_ net633 VGND VGND VPWR VPWR top0.pid_d.out\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13603_ net1027 _05520_ _05521_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__and3_1
X_17371_ net405 _09351_ _09354_ _09357_ VGND VGND VPWR VPWR _09358_ sky130_fd_sc_hd__a22o_1
X_14583_ _06785_ _06788_ VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_156_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26569_ clknet_leaf_54_clk_sys _00192_ net667 VGND VGND VPWR VPWR top0.pid_q.curr_error\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_131_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16322_ _08377_ _08379_ _08348_ VGND VGND VPWR VPWR _08412_ sky130_fd_sc_hd__o21ba_1
X_19110_ top0.pid_d.out\[15\] top0.pid_d.curr_int\[15\] VGND VGND VPWR VPWR _11082_
+ sky130_fd_sc_hd__xor2_2
X_13534_ _05743_ _05744_ _05745_ _05746_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_67_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19041_ _11012_ _11013_ VGND VGND VPWR VPWR _11014_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16253_ _08048_ _08340_ _08343_ VGND VGND VPWR VPWR _08344_ sky130_fd_sc_hd__and3_1
X_13465_ net42 _05520_ _05521_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15204_ _07168_ _07173_ VGND VGND VPWR VPWR _07303_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16184_ _08192_ _08194_ _08193_ VGND VGND VPWR VPWR _08276_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13396_ top0.matmul0.beta_pass\[11\] _05434_ _05469_ _05463_ top0.c_out_calc\[11\]
+ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__a32o_2
XFILLER_0_50_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15135_ _07231_ _07232_ _07233_ VGND VGND VPWR VPWR _07234_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19943_ net183 _11810_ _11811_ _11812_ _11813_ VGND VGND VPWR VPWR _11814_ sky130_fd_sc_hd__o221a_1
X_15066_ _07163_ _07164_ VGND VGND VPWR VPWR _07165_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14017_ net39 _05517_ _06113_ _06114_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__a22o_1
X_19874_ _11717_ _11732_ VGND VGND VPWR VPWR _11750_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18825_ _10633_ _10800_ VGND VGND VPWR VPWR _10801_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18756_ _10610_ _10625_ _10627_ VGND VGND VPWR VPWR _10733_ sky130_fd_sc_hd__a21oi_2
X_15968_ _08000_ _08062_ VGND VGND VPWR VPWR _08063_ sky130_fd_sc_hd__xnor2_2
X_17707_ net386 _09394_ _09693_ net391 VGND VGND VPWR VPWR _09694_ sky130_fd_sc_hd__a22o_1
X_14919_ _07080_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__clkbuf_1
X_18687_ _10658_ _10664_ VGND VGND VPWR VPWR _10665_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15899_ _07705_ _07992_ _07994_ _07710_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__o211a_1
X_17638_ net403 net398 net344 net348 VGND VGND VPWR VPWR _09625_ sky130_fd_sc_hd__and4_1
XFILLER_0_37_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17569_ _09551_ _09553_ VGND VGND VPWR VPWR _09556_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19308_ _11248_ _11239_ _11235_ VGND VGND VPWR VPWR _11249_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20580_ net270 net258 VGND VGND VPWR VPWR _12429_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19239_ top0.pid_d.prev_error\[7\] top0.pid_d.curr_error\[7\] VGND VGND VPWR VPWR
+ _11186_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22250_ _01806_ _01810_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21201_ _12967_ _12996_ _12995_ VGND VGND VPWR VPWR _13045_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22181_ _01724_ _01722_ _01741_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__a21o_2
XFILLER_0_197_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21132_ _11673_ _12785_ VGND VGND VPWR VPWR _12977_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout402 top0.pid_d.mult0.a\[6\] VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__clkbuf_2
X_25940_ _05145_ _05152_ _12014_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__a21oi_1
X_21063_ net247 _11726_ _12045_ VGND VGND VPWR VPWR _12909_ sky130_fd_sc_hd__a21oi_1
Xfanout413 net414 VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__clkbuf_4
Xfanout424 top0.pid_d.mult0.a\[1\] VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__buf_4
Xfanout435 net436 VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__clkbuf_4
Xfanout446 top0.pid_q.mult0.b\[14\] VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__buf_4
X_20014_ _11879_ VGND VGND VPWR VPWR _11880_ sky130_fd_sc_hd__inv_2
Xfanout457 top0.pid_q.mult0.b\[10\] VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__buf_4
X_25871_ top0.matmul0.alpha_pass\[7\] top0.matmul0.beta_pass\[7\] top0.matmul0.beta_pass\[8\]
+ net1024 VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__o211a_1
Xfanout468 net469 VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_129_Left_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout479 net482 VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__clkbuf_4
X_24822_ _04173_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24753_ _04020_ _04025_ _04017_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__a21o_1
X_21965_ _01208_ _01526_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23704_ net567 net560 top0.matmul0.matmul_stage_inst.e\[9\] VGND VGND VPWR VPWR _03062_
+ sky130_fd_sc_hd__o21a_4
Xclkbuf_leaf_49_clk_sys clknet_3_6__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_49_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_20916_ net232 net218 VGND VGND VPWR VPWR _12764_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_96_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24684_ _04036_ _03918_ _04037_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_90_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21896_ net150 net128 VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__xor2_2
XFILLER_0_84_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26423_ clknet_leaf_58_clk_sys _00064_ net644 VGND VGND VPWR VPWR top0.kpq\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23635_ net568 net573 top0.matmul0.matmul_stage_inst.f\[6\] VGND VGND VPWR VPWR _02993_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_193_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20847_ net227 net218 VGND VGND VPWR VPWR _12696_ sky130_fd_sc_hd__nor2b_2
Xfanout20 net22 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
XFILLER_0_65_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout31 net32 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_4
XFILLER_0_49_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout42 top0.periodTop_r\[9\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_4
XFILLER_0_7_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout53 top0.periodTop_r\[5\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
X_26354_ spi0.data_packed\[75\] spi0.data_packed\[76\] net690 VGND VGND VPWR VPWR
+ _05409_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_138_Left_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23566_ net966 top0.matmul0.b\[6\] _02948_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__mux2_1
Xfanout64 top0.periodTop_r\[1\] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_4
X_20778_ _12624_ _12625_ VGND VGND VPWR VPWR _12627_ sky130_fd_sc_hd__nor2_1
Xfanout75 top0.matmul0.alpha_pass\[8\] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_2
X_25305_ _04576_ _04582_ _04583_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout86 net89 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_4
XFILLER_0_174_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22517_ _02071_ _02072_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__nand2_1
Xfanout97 top0.cordic0.vec\[1\]\[14\] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_4
XFILLER_0_107_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26285_ net947 VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23497_ _02913_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25236_ _04579_ _04581_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__or2_1
X_13250_ _05462_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__buf_6
XFILLER_0_150_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22448_ _01258_ _01683_ _01738_ _02004_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25167_ _04506_ _04514_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_161_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22379_ _01924_ _01829_ _01937_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24118_ _03473_ _03475_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__nand2_1
X_25098_ _04441_ _04446_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_202_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24049_ _03393_ _03397_ _03406_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__a21o_1
X_16940_ top0.matmul0.beta_pass\[9\] _05437_ top0.currT_r\[9\] VGND VGND VPWR VPWR
+ _08998_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_198_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_147_Left_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16871_ _05438_ _08933_ VGND VGND VPWR VPWR _08934_ sky130_fd_sc_hd__nand2_1
X_18610_ _10505_ _10581_ _10584_ _10585_ _10588_ VGND VGND VPWR VPWR _10589_ sky130_fd_sc_hd__a221o_1
X_15822_ _07913_ _07917_ VGND VGND VPWR VPWR _07918_ sky130_fd_sc_hd__xor2_2
X_19590_ top0.cordic0.slte0.opB\[8\] top0.cordic0.slte0.opA\[8\] VGND VGND VPWR VPWR
+ _11479_ sky130_fd_sc_hd__xor2_1
X_18541_ net387 _10203_ _09364_ VGND VGND VPWR VPWR _10520_ sky130_fd_sc_hd__o21ai_1
X_15753_ net460 net523 VGND VGND VPWR VPWR _07850_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14704_ net817 _06280_ _06907_ _05465_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__a22o_1
X_18472_ _10450_ _10451_ VGND VGND VPWR VPWR _10452_ sky130_fd_sc_hd__xor2_2
X_15684_ _07781_ net511 _07535_ VGND VGND VPWR VPWR _07782_ sky130_fd_sc_hd__or3b_1
X_14635_ net40 _06351_ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__nand2_1
X_17423_ _09408_ _09409_ VGND VGND VPWR VPWR _09410_ sky130_fd_sc_hd__xor2_2
XFILLER_0_158_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14566_ _06766_ _06771_ VGND VGND VPWR VPWR _06772_ sky130_fd_sc_hd__xor2_1
X_17354_ net423 net340 VGND VGND VPWR VPWR _09341_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13517_ _05722_ _05729_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__xnor2_2
X_16305_ _08393_ _08395_ VGND VGND VPWR VPWR _08396_ sky130_fd_sc_hd__nand2_1
X_17285_ _09280_ _09276_ _09281_ VGND VGND VPWR VPWR _09282_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14497_ _06700_ _06703_ VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19024_ _10845_ _10958_ _10939_ VGND VGND VPWR VPWR _10997_ sky130_fd_sc_hd__a21o_1
X_16236_ top0.pid_q.out\[8\] top0.pid_q.curr_int\[8\] VGND VGND VPWR VPWR _08327_
+ sky130_fd_sc_hd__xnor2_1
X_13448_ _05656_ _05660_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16167_ _08255_ _08258_ VGND VGND VPWR VPWR _08259_ sky130_fd_sc_hd__xnor2_4
X_13379_ _05589_ _05591_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15118_ _07210_ _07215_ _07216_ VGND VGND VPWR VPWR _07217_ sky130_fd_sc_hd__nand3_1
X_16098_ _08093_ _08095_ _08190_ VGND VGND VPWR VPWR _08191_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_121_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19926_ net190 _11797_ net201 VGND VGND VPWR VPWR _11798_ sky130_fd_sc_hd__o21ai_1
X_15049_ _07146_ _07147_ VGND VGND VPWR VPWR _07148_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19857_ _11713_ _11721_ net241 VGND VGND VPWR VPWR _11734_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_177_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18808_ _10777_ _10783_ VGND VGND VPWR VPWR _10784_ sky130_fd_sc_hd__xor2_2
X_19788_ net1014 _11669_ net174 VGND VGND VPWR VPWR _11670_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18739_ _10633_ _10715_ VGND VGND VPWR VPWR _10716_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_50_clk_sys clknet_3_6__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_50_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21750_ net119 net102 VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_176_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20701_ net285 net273 _12278_ VGND VGND VPWR VPWR _12550_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21681_ _01128_ _01110_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23420_ _02855_ _02857_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_176_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20632_ net294 _12284_ VGND VGND VPWR VPWR _12481_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_202_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23351_ _01408_ _11548_ _02792_ _02794_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20563_ _12371_ VGND VGND VPWR VPWR _12412_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22302_ _01775_ _01783_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__nor2_1
X_26070_ top0.a_in_matmul\[9\] _05254_ _05230_ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__mux2_1
X_23282_ _11425_ _02728_ _02729_ net215 _11580_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__a32o_1
X_20494_ _12259_ _12342_ VGND VGND VPWR VPWR _12343_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25021_ _03248_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__clkbuf_4
X_22233_ _01774_ _01792_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22164_ _01231_ _01235_ _01232_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_160_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21115_ net1021 _12960_ VGND VGND VPWR VPWR _12961_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26972_ clknet_leaf_29_clk_sys _00589_ net624 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_22095_ _01628_ _01632_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__and2b_1
Xfanout210 net211 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_4
Xfanout221 net224 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_8
Xfanout232 net233 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_2
X_25923_ _05128_ _05134_ _05137_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__o21a_1
X_21046_ _12861_ _12890_ _12891_ VGND VGND VPWR VPWR _12892_ sky130_fd_sc_hd__a21o_1
Xfanout243 top0.cordic0.vec\[0\]\[12\] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_2
Xfanout254 net256 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_4
Xfanout265 net268 VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__buf_4
Xfanout276 net279 VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__buf_4
XFILLER_0_199_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout287 net293 VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__buf_2
X_25854_ _05071_ _05074_ _05070_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__a21oi_1
Xfanout298 net299 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__buf_2
X_24805_ _04066_ _04152_ VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__nand2_1
X_25785_ _05425_ _05014_ _05016_ net207 VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22997_ top0.svm0.delta\[10\] _02499_ net169 VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24736_ _04027_ _04012_ _04011_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_69_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21948_ net160 net137 _01502_ _01507_ _01509_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__a311o_1
X_24667_ _03004_ _03005_ _03103_ _03104_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__o22a_2
X_21879_ net161 net166 VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__or2b_1
XFILLER_0_194_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14420_ _06622_ _06627_ VGND VGND VPWR VPWR _06628_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_37_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26406_ clknet_leaf_98_clk_sys _00047_ net632 VGND VGND VPWR VPWR top0.kpd\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_23618_ net569 net572 top0.matmul0.matmul_stage_inst.f\[4\] VGND VGND VPWR VPWR _02976_
+ sky130_fd_sc_hd__o21a_4
XFILLER_0_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24598_ _03950_ _03952_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__xor2_1
XFILLER_0_181_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14351_ _06510_ _06558_ _06559_ VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26337_ _05400_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__clkbuf_1
X_23549_ top0.a_in_matmul\[14\] top0.matmul0.a\[14\] _02937_ VGND VGND VPWR VPWR _02941_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13302_ net43 _05497_ _05513_ _05514_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__a22o_1
X_17070_ _09045_ top0.pid_q.curr_error\[12\] _09096_ VGND VGND VPWR VPWR _09109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14282_ _06488_ _06491_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_135_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26268_ spi0.data_packed\[32\] spi0.data_packed\[33\] net688 VGND VGND VPWR VPWR
+ _05366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16021_ _08013_ _08015_ _08114_ VGND VGND VPWR VPWR _08115_ sky130_fd_sc_hd__a21oi_2
X_25219_ _04555_ _04564_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13233_ _05452_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__buf_1
XFILLER_0_21_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26199_ net209 top0.svm0.out_valid net206 VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17972_ _09934_ _09956_ VGND VGND VPWR VPWR _09958_ sky130_fd_sc_hd__nand2_1
X_19711_ _11572_ _11440_ _11595_ _11427_ VGND VGND VPWR VPWR _11596_ sky130_fd_sc_hd__o2bb2a_1
X_16923_ net466 _08890_ _08982_ _08930_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19642_ _11424_ _11529_ VGND VGND VPWR VPWR _11530_ sky130_fd_sc_hd__nor2_1
X_16854_ top0.matmul0.beta_pass\[3\] _05438_ VGND VGND VPWR VPWR _08918_ sky130_fd_sc_hd__nand2_1
X_15805_ _07899_ _07900_ VGND VGND VPWR VPWR _07901_ sky130_fd_sc_hd__nor2_1
X_19573_ _11459_ _11460_ _11453_ _11461_ VGND VGND VPWR VPWR _11462_ sky130_fd_sc_hd__a211o_1
X_13997_ top0.matmul0.alpha_pass\[1\] _05435_ _05474_ VGND VGND VPWR VPWR _06210_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_99_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16785_ top0.pid_q.mult0.a\[2\] _08856_ _08859_ net787 _08865_ VGND VGND VPWR VPWR
+ _00151_ sky130_fd_sc_hd__a221o_1
XFILLER_0_189_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18524_ _10490_ _10503_ VGND VGND VPWR VPWR _10504_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15736_ net457 net526 VGND VGND VPWR VPWR _07833_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18455_ _10406_ _10407_ _10402_ VGND VGND VPWR VPWR _10435_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15667_ _07630_ _07634_ _07764_ VGND VGND VPWR VPWR _07765_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17406_ _09392_ _09386_ VGND VGND VPWR VPWR _09393_ sky130_fd_sc_hd__or2b_1
X_14618_ _06773_ _06821_ _06822_ VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__o21ai_2
X_18386_ net334 net373 VGND VGND VPWR VPWR _10367_ sky130_fd_sc_hd__nand2_1
X_15598_ _07616_ _07696_ VGND VGND VPWR VPWR _07697_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14549_ _06701_ _06702_ _06754_ VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__o21a_1
X_17337_ _09326_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17268_ top0.matmul0.beta_pass\[3\] _09267_ net563 VGND VGND VPWR VPWR _09268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19007_ _10979_ _10980_ VGND VGND VPWR VPWR _10981_ sky130_fd_sc_hd__or2b_1
XFILLER_0_180_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16219_ _08304_ _08310_ VGND VGND VPWR VPWR _08311_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17199_ _09207_ _09203_ top0.pid_q.curr_int\[9\] VGND VGND VPWR VPWR _09208_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_11_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19909_ net176 _11648_ VGND VGND VPWR VPWR _11783_ sky130_fd_sc_hd__nand2_1
Xhold18 top0.cordic0.cos\[3\] VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 top0.svm0.tB\[0\] VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__dlygate4sd3_1
X_22920_ top0.svm0.counter\[0\] net555 VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_4__f_clk_mosi clknet_0_clk_mosi VGND VGND VPWR VPWR clknet_3_4__leaf_clk_mosi
+ sky130_fd_sc_hd__clkbuf_16
X_22851_ _02360_ top0.svm0.tA\[9\] _02370_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21802_ _01335_ _01353_ _01348_ _01362_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__o211a_1
X_25570_ _04872_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__clkbuf_1
X_22782_ _07113_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24521_ _03874_ _03875_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__xnor2_1
X_21733_ net141 _01294_ VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27240_ clknet_3_7__leaf_clk_mosi _00854_ VGND VGND VPWR VPWR spi0.data_packed\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_24452_ _03076_ _03077_ _03196_ _03197_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21664_ _01223_ _01225_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__xor2_1
XFILLER_0_176_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23403_ _02838_ _02842_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__xor2_1
X_27171_ clknet_leaf_12_clk_sys _00785_ net618 VGND VGND VPWR VPWR top0.periodTop_r\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_20615_ net274 net263 net249 VGND VGND VPWR VPWR _12464_ sky130_fd_sc_hd__and3_1
XFILLER_0_188_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24383_ _03186_ _03187_ _03739_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_145_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21595_ net164 _01155_ _01156_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26122_ spi0.data_packed\[19\] _05279_ _05280_ net934 VGND VGND VPWR VPWR _00800_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23334_ _01135_ _02778_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__nor2_1
X_20546_ _12386_ _12392_ _12393_ _12394_ _12375_ VGND VGND VPWR VPWR _12395_ sky130_fd_sc_hd__o221a_1
XFILLER_0_104_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26053_ net76 _05237_ _05241_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23265_ _02709_ _02710_ _02712_ _02713_ _11572_ net182 VGND VGND VPWR VPWR _02714_
+ sky130_fd_sc_hd__mux4_1
X_20477_ net298 net282 VGND VGND VPWR VPWR _12326_ sky130_fd_sc_hd__nor2_1
X_25004_ _04273_ _04274_ _04353_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_197_Right_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22216_ _01211_ net102 VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__nand2_4
X_23196_ _05719_ _07034_ _02648_ net838 VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__a22o_1
X_22147_ _01707_ _01708_ net149 VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__mux2_1
X_26955_ clknet_leaf_13_clk_sys _00572_ net613 VGND VGND VPWR VPWR top0.matmul0.b\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_22078_ _01190_ _01639_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__xnor2_2
X_13920_ _05725_ _05728_ _06132_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__a21o_2
X_25906_ net429 _05114_ _05121_ _05110_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__a211o_1
X_21029_ _12749_ _12746_ _12802_ VGND VGND VPWR VPWR _12876_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_199_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26886_ clknet_leaf_38_clk_sys _00503_ net677 VGND VGND VPWR VPWR top0.svm0.tB\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13851_ _06060_ _06063_ _06053_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25837_ net76 top0.matmul0.beta_pass\[5\] VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16570_ net497 _08656_ VGND VGND VPWR VPWR _08657_ sky130_fd_sc_hd__nand2_1
X_13782_ _05979_ _05994_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__xnor2_2
X_25768_ top0.matmul0.matmul_stage_inst.a\[12\] _04901_ _05457_ VGND VGND VPWR VPWR
+ _05005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15521_ _07618_ _07619_ VGND VGND VPWR VPWR _07620_ sky130_fd_sc_hd__xnor2_1
X_24719_ _03765_ _03743_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25699_ net862 _04925_ _04963_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18240_ _10097_ _10127_ VGND VGND VPWR VPWR _10223_ sky130_fd_sc_hd__or2_1
X_15452_ net520 net471 VGND VGND VPWR VPWR _07551_ sky130_fd_sc_hd__nand2_1
X_14403_ _06551_ _06611_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_182_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18171_ _10073_ _10154_ VGND VGND VPWR VPWR _10155_ sky130_fd_sc_hd__xnor2_1
X_15383_ _07456_ _07481_ VGND VGND VPWR VPWR _07482_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14334_ _06476_ _06542_ VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17122_ _09140_ VGND VGND VPWR VPWR _09141_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17053_ net983 _09100_ _09102_ _08894_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__a22o_1
X_14265_ _06464_ _06467_ _06393_ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16004_ _08020_ _08022_ _08021_ VGND VGND VPWR VPWR _08098_ sky130_fd_sc_hd__o21a_1
X_13216_ _05440_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__clkbuf_4
X_14196_ _06401_ _06406_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_164_Right_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17955_ _09863_ _09864_ _09940_ VGND VGND VPWR VPWR _09941_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16906_ _08965_ _08966_ VGND VGND VPWR VPWR _08967_ sky130_fd_sc_hd__xnor2_1
X_17886_ _09869_ _09872_ VGND VGND VPWR VPWR _09873_ sky130_fd_sc_hd__xor2_1
X_19625_ _11513_ VGND VGND VPWR VPWR _11514_ sky130_fd_sc_hd__buf_2
X_16837_ top0.currT_r\[1\] top0.matmul0.beta_pass\[1\] VGND VGND VPWR VPWR _08902_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19556_ net179 _11444_ VGND VGND VPWR VPWR _11445_ sky130_fd_sc_hd__nand2_2
X_16768_ net544 net1019 _08848_ _08851_ VGND VGND VPWR VPWR _08852_ sky130_fd_sc_hd__a31o_1
X_18507_ _10480_ _10486_ VGND VGND VPWR VPWR _10487_ sky130_fd_sc_hd__xnor2_1
X_15719_ _07814_ _07815_ VGND VGND VPWR VPWR _07816_ sky130_fd_sc_hd__xnor2_1
X_19487_ net435 _11240_ _11380_ net441 VGND VGND VPWR VPWR _11381_ sky130_fd_sc_hd__a22o_1
X_16699_ _08746_ _08783_ VGND VGND VPWR VPWR _08784_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18438_ _10318_ _10322_ VGND VGND VPWR VPWR _10419_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18369_ net390 net364 _10349_ _09429_ _09363_ VGND VGND VPWR VPWR _10350_ sky130_fd_sc_hd__a32o_1
XFILLER_0_84_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20400_ net289 _12047_ VGND VGND VPWR VPWR _12249_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21380_ _12705_ _12853_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20331_ _12072_ VGND VGND VPWR VPWR _12180_ sky130_fd_sc_hd__buf_6
XFILLER_0_4_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23050_ top0.svm0.counter\[12\] _02550_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__xnor2_1
X_20262_ _11408_ _11550_ net282 _12068_ VGND VGND VPWR VPWR _12111_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22001_ _01313_ _01561_ _01562_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20193_ net252 net240 VGND VGND VPWR VPWR _12042_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_179_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23952_ _03243_ _03244_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__xnor2_2
X_26740_ clknet_leaf_101_clk_sys _00357_ net587 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[15\]
+ sky130_fd_sc_hd__dfstp_1
X_22903_ _02367_ top0.svm0.tC\[8\] _02419_ _02420_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__o22a_1
X_26671_ clknet_leaf_82_clk_sys _00288_ net646 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_23883_ _03239_ _03240_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__xnor2_2
X_22834_ _02298_ top0.svm0.tA\[0\] _02353_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__a21o_1
X_25622_ top0.matmul0.matmul_stage_inst.a\[14\] _04902_ _05458_ VGND VGND VPWR VPWR
+ _04903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25553_ _04863_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__clkbuf_1
X_22765_ net970 _02292_ _02295_ top0.pid_q.curr_int\[9\] VGND VGND VPWR VPWR _00428_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24504_ _03751_ _03846_ _03857_ _03652_ _03858_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_137_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21716_ _01262_ _01264_ VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__and2_1
X_25484_ _04820_ _04826_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22696_ _01924_ _02246_ _01948_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24435_ _02998_ _03000_ _03061_ _03062_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27223_ clknet_3_5__leaf_clk_mosi _00837_ VGND VGND VPWR VPWR spi0.data_packed\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21647_ _01076_ _01208_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_151_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27154_ clknet_leaf_10_clk_sys _00768_ net602 VGND VGND VPWR VPWR top0.a_in_matmul\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_191_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24366_ _03252_ _03198_ _03722_ _03120_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21578_ _01135_ _01139_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__nor2_1
X_26105_ net741 _05276_ _05278_ net1025 VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23317_ _02707_ _02719_ _02744_ net140 _01123_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__o221a_1
XFILLER_0_160_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27085_ clknet_leaf_8_clk_sys _00702_ net592 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20529_ _12283_ _12314_ _12322_ VGND VGND VPWR VPWR _12378_ sky130_fd_sc_hd__a21o_1
X_24297_ _03301_ _03653_ _03630_ _03620_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__a211o_2
XFILLER_0_34_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14050_ _06261_ _06262_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__nor2_2
XFILLER_0_120_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26036_ top0.pid_d.out\[2\] _05198_ _05199_ spi0.data_packed\[66\] VGND VGND VPWR
+ VPWR _05228_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23248_ _11649_ _02696_ _11954_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23179_ _07115_ _02642_ _02308_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17740_ _09413_ VGND VGND VPWR VPWR _09727_ sky130_fd_sc_hd__inv_2
X_14952_ spi0.data_packed\[18\] top0.kiq\[2\] _07097_ VGND VGND VPWR VPWR _07098_
+ sky130_fd_sc_hd__mux2_1
X_26938_ clknet_leaf_9_clk_sys _00555_ net595 VGND VGND VPWR VPWR top0.matmul0.a\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13903_ _06112_ _06115_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_199_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17671_ net414 net330 VGND VGND VPWR VPWR _09658_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26869_ clknet_leaf_40_clk_sys _00486_ net678 VGND VGND VPWR VPWR top0.svm0.tA\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14883_ _07061_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19410_ _11311_ _11312_ VGND VGND VPWR VPWR _11313_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16622_ _08636_ _08641_ _08634_ VGND VGND VPWR VPWR _08708_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_134_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13834_ _05501_ _06046_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__nor2_1
XFILLER_0_202_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19341_ _11277_ VGND VGND VPWR VPWR _11278_ sky130_fd_sc_hd__buf_2
XFILLER_0_187_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16553_ _08638_ _08639_ VGND VGND VPWR VPWR _08640_ sky130_fd_sc_hd__xor2_1
X_13765_ _05962_ _05961_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_97_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_97_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15504_ net517 _07258_ VGND VGND VPWR VPWR _07603_ sky130_fd_sc_hd__and2_1
X_19272_ _11214_ _11205_ _11215_ VGND VGND VPWR VPWR _11216_ sky130_fd_sc_hd__a21o_1
X_13696_ _05805_ _05731_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__nor2_1
X_16484_ net466 _08141_ net461 VGND VGND VPWR VPWR _08572_ sky130_fd_sc_hd__o21a_1
XFILLER_0_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18223_ net400 net366 _10204_ _10205_ VGND VGND VPWR VPWR _10206_ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15435_ _07266_ _07280_ _07294_ VGND VGND VPWR VPWR _07534_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_72_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18154_ _09993_ _09994_ VGND VGND VPWR VPWR _10138_ sky130_fd_sc_hd__nand2_1
X_15366_ _07450_ _07464_ VGND VGND VPWR VPWR _07465_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17105_ top0.pid_q.curr_error\[11\] _08860_ _09116_ VGND VGND VPWR VPWR _09129_ sky130_fd_sc_hd__and3_1
X_14317_ _06521_ _06526_ VGND VGND VPWR VPWR _06527_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15297_ _07390_ _07391_ _07395_ VGND VGND VPWR VPWR _07396_ sky130_fd_sc_hd__o21bai_1
X_18085_ top0.pid_d.curr_int\[2\] _09983_ _10068_ VGND VGND VPWR VPWR _10069_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold307 top0.cordic0.sin\[13\] VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14248_ _06450_ _06451_ _06458_ VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__a21o_1
X_17036_ top0.matmul0.beta_pass\[15\] _05438_ VGND VGND VPWR VPWR _09088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14179_ _06358_ _06366_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18987_ _10939_ _10960_ VGND VGND VPWR VPWR _10961_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17938_ _09844_ _09845_ _09846_ VGND VGND VPWR VPWR _09924_ sky130_fd_sc_hd__o21a_1
XFILLER_0_178_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17869_ _09848_ _09855_ VGND VGND VPWR VPWR _09856_ sky130_fd_sc_hd__xnor2_2
X_19608_ top0.cordic0.slte0.opA\[13\] _11465_ top0.cordic0.slte0.opB\[13\] VGND VGND
+ VPWR VPWR _11497_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_36_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20880_ _12727_ _12728_ VGND VGND VPWR VPWR _12729_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19539_ _11426_ _11428_ VGND VGND VPWR VPWR _11429_ sky130_fd_sc_hd__nor2_1
XFILLER_0_191_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22550_ net104 _02102_ _02104_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_200_Right_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21501_ _01062_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_101_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22481_ _01953_ _01976_ _02037_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__o21a_1
X_24220_ _03576_ _03577_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__xor2_1
XFILLER_0_134_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21432_ _00916_ _00927_ _00956_ _00954_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__a31o_1
XFILLER_0_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24151_ _03500_ _03505_ _03508_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__or3_2
XFILLER_0_115_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21363_ _00929_ _13182_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23102_ net896 _02600_ _02601_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__a21o_1
X_20314_ _12097_ _12091_ _12162_ VGND VGND VPWR VPWR _12163_ sky130_fd_sc_hd__a21oi_4
X_24082_ _03279_ _03281_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21294_ _13040_ _13042_ _13018_ VGND VGND VPWR VPWR _13137_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23033_ _02309_ top0.svm0.counter\[15\] _02306_ _02534_ VGND VGND VPWR VPWR _02535_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_13_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20245_ net255 net250 VGND VGND VPWR VPWR _12094_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_122_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_110_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20176_ _12027_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24984_ _04315_ _04318_ _04333_ _04235_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26723_ clknet_leaf_78_clk_sys _00340_ net633 VGND VGND VPWR VPWR top0.pid_d.curr_int\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_23935_ _03269_ _03266_ _03231_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__o21ai_2
X_23866_ _03206_ _03223_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__xnor2_2
X_26654_ clknet_leaf_76_clk_sys _00271_ net639 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22817_ top0.svm0.counter\[9\] top0.svm0.tA\[9\] VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25605_ net70 top0.matmul0.cos\[6\] VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23797_ net569 net573 top0.matmul0.matmul_stage_inst.f\[2\] VGND VGND VPWR VPWR _03155_
+ sky130_fd_sc_hd__o21ai_2
X_26585_ clknet_leaf_54_clk_sys _00208_ net673 VGND VGND VPWR VPWR top0.pid_q.prev_error\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13550_ _05689_ _05761_ _05762_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25536_ _04854_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__clkbuf_1
X_22748_ _11413_ _02289_ net176 VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25467_ _04721_ _04809_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__nand2_1
X_13481_ _05499_ _05507_ _05482_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__a21o_1
X_22679_ _02209_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15220_ _07309_ _07312_ _07318_ VGND VGND VPWR VPWR _07319_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_192_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24418_ _03763_ _03773_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__xnor2_2
X_27206_ clknet_leaf_92_clk_sys _00820_ net600 VGND VGND VPWR VPWR top0.cordic0.slte0.opB\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_25398_ _04683_ _04740_ _04741_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15151_ _07222_ _07225_ _07249_ VGND VGND VPWR VPWR _07250_ sky130_fd_sc_hd__and3_1
X_24349_ _03210_ _03211_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__nor2_1
X_27137_ clknet_leaf_12_clk_sys _00751_ net616 VGND VGND VPWR VPWR top0.b_in_matmul\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14102_ _06206_ _06207_ net37 _05472_ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27068_ clknet_leaf_2_clk_sys _00685_ net583 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.c\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15082_ net535 net460 VGND VGND VPWR VPWR _07181_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14033_ _06244_ _06245_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__xor2_1
X_26019_ _05215_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__clkbuf_1
X_18910_ _10800_ _10884_ VGND VGND VPWR VPWR _10885_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19890_ _11742_ _11753_ _11739_ VGND VGND VPWR VPWR _11765_ sky130_fd_sc_hd__o21a_1
X_18841_ _10707_ _10729_ _10727_ VGND VGND VPWR VPWR _10817_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18772_ _10747_ _10748_ VGND VGND VPWR VPWR _10749_ sky130_fd_sc_hd__and2b_1
X_15984_ top0.pid_q.out\[4\] top0.pid_q.curr_int\[4\] VGND VGND VPWR VPWR _08079_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17723_ net386 _09360_ _09692_ VGND VGND VPWR VPWR _09710_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_145_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14935_ spi0.data_packed\[42\] top0.kid\[10\] _07086_ VGND VGND VPWR VPWR _07089_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17654_ _09636_ _09640_ VGND VGND VPWR VPWR _09641_ sky130_fd_sc_hd__xnor2_1
X_14866_ _07052_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__clkbuf_1
X_16605_ _08653_ _08658_ _08629_ VGND VGND VPWR VPWR _08691_ sky130_fd_sc_hd__o21a_1
XFILLER_0_202_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13817_ net62 _05496_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__nand2_1
X_17585_ net418 net423 net415 VGND VGND VPWR VPWR _09572_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14797_ _06942_ _06946_ _06997_ VGND VGND VPWR VPWR _06998_ sky130_fd_sc_hd__or3b_1
XFILLER_0_86_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19324_ _11262_ _11263_ VGND VGND VPWR VPWR _11264_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16536_ _08622_ _08621_ top0.pid_q.out\[12\] VGND VGND VPWR VPWR _08623_ sky130_fd_sc_hd__mux2_1
X_13748_ net59 _05520_ _05521_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__and3_1
XFILLER_0_174_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19255_ net1024 _11190_ VGND VGND VPWR VPWR _11201_ sky130_fd_sc_hd__xor2_1
X_16467_ net452 net503 VGND VGND VPWR VPWR _08555_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13679_ _05890_ _05891_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18206_ _10187_ _10188_ VGND VGND VPWR VPWR _10189_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15418_ _07427_ _07429_ VGND VGND VPWR VPWR _07517_ sky130_fd_sc_hd__nor2_1
X_19186_ _11135_ _11136_ VGND VGND VPWR VPWR _11138_ sky130_fd_sc_hd__nand2_1
X_16398_ _08483_ _08486_ VGND VGND VPWR VPWR _08487_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18137_ _10025_ _10027_ _10120_ VGND VGND VPWR VPWR _10121_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_26_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15349_ net533 net482 _07403_ _07447_ VGND VGND VPWR VPWR _07448_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold104 top0.svm0.tB\[13\] VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold115 top0.pid_d.prev_int\[15\] VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 top0.pid_q.prev_error\[10\] VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__dlygate4sd3_1
X_18068_ _10039_ _10052_ VGND VGND VPWR VPWR _10053_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_106_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold137 top0.svm0.tB\[3\] VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 top0.svm0.tC\[8\] VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__dlygate4sd3_1
X_17019_ top0.pid_q.prev_error\[13\] top0.pid_q.curr_error\[13\] VGND VGND VPWR VPWR
+ _09072_ sky130_fd_sc_hd__and2_1
Xhold159 top0.matmul0.matmul_stage_inst.c\[2\] VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout606 net630 VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout617 net620 VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20030_ _11518_ _11891_ _11894_ _11426_ VGND VGND VPWR VPWR _11895_ sky130_fd_sc_hd__o211a_1
Xfanout628 net629 VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__clkbuf_2
Xfanout639 net654 VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__clkbuf_4
X_21981_ _01454_ _01480_ _01529_ _01541_ _01542_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__o221a_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23720_ _03061_ _03062_ _03076_ _03077_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__o22a_4
X_20932_ _12135_ _12779_ VGND VGND VPWR VPWR _12780_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_179_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23651_ _02976_ _02977_ _02988_ _02990_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__o22a_2
XFILLER_0_89_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20863_ _12709_ _12710_ _12701_ VGND VGND VPWR VPWR _12712_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22602_ net112 net95 _01166_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__or3_1
XFILLER_0_193_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26370_ spi0.opcode\[3\] spi0.opcode\[4\] net691 VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23582_ net1009 top0.matmul0.b\[14\] _02948_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20794_ _12642_ VGND VGND VPWR VPWR _12643_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25321_ _04521_ _04643_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22533_ net210 _02086_ _02088_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_107_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25252_ _04597_ _04526_ _04598_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__o21a_1
XFILLER_0_173_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22464_ _01312_ _02020_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24203_ _03017_ _03252_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__nor2_1
X_21415_ _00975_ _00981_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25183_ _04382_ _04528_ _04529_ _04530_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22395_ _01921_ _01928_ _01952_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24134_ _03045_ _03046_ _03076_ _03077_ VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__o22a_1
X_21346_ _13157_ _13187_ VGND VGND VPWR VPWR _13188_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_45_clk_sys clknet_3_7__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_45_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24065_ _03378_ _03418_ _03422_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__a21boi_1
X_21277_ net239 _13031_ _13118_ _13119_ VGND VGND VPWR VPWR _13120_ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23016_ top0.svm0.counter\[13\] _02306_ _02517_ _02519_ VGND VGND VPWR VPWR _00455_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20228_ _11758_ _12075_ _12074_ VGND VGND VPWR VPWR _12077_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_60_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20159_ _05437_ top0.svm0.out_valid net206 VGND VGND VPWR VPWR _12011_ sky130_fd_sc_hd__mux2_1
X_24967_ _04170_ _04316_ _04317_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14720_ _06921_ _06922_ VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__xor2_1
X_26706_ clknet_leaf_84_clk_sys _00323_ net641 VGND VGND VPWR VPWR top0.pid_d.prev_error\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_23918_ _03272_ _03273_ _03274_ _03275_ _03233_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__a32o_2
X_24898_ _04156_ _04247_ _04245_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14651_ _06755_ _06756_ _06855_ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__o21a_1
XFILLER_0_157_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26637_ clknet_leaf_82_clk_sys _00254_ net638 VGND VGND VPWR VPWR top0.pid_d.out\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_23849_ _03036_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13602_ _05810_ _05813_ _05814_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_68_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17370_ _09351_ _09356_ VGND VGND VPWR VPWR _09357_ sky130_fd_sc_hd__nor2_1
X_14582_ _06723_ _06786_ _06787_ VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__and3_1
X_26568_ clknet_leaf_52_clk_sys _00191_ net673 VGND VGND VPWR VPWR top0.pid_q.curr_error\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16321_ _08393_ _08410_ VGND VGND VPWR VPWR _08411_ sky130_fd_sc_hd__nand2_1
X_25519_ _04845_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__clkbuf_1
X_13533_ _05672_ _05661_ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__nand2_1
X_26499_ clknet_leaf_74_clk_sys _00122_ net655 VGND VGND VPWR VPWR top0.pid_d.prev_int\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19040_ _10957_ _10955_ _10845_ VGND VGND VPWR VPWR _11013_ sky130_fd_sc_hd__mux2_2
XFILLER_0_165_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13464_ net43 _05517_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__nand2_1
X_16252_ net469 _08342_ VGND VGND VPWR VPWR _08343_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15203_ _07240_ _07301_ VGND VGND VPWR VPWR _07302_ sky130_fd_sc_hd__xor2_1
XFILLER_0_63_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13395_ top0.matmul0.alpha_pass\[11\] _05434_ _05467_ VGND VGND VPWR VPWR _05608_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16183_ _08271_ _08274_ VGND VGND VPWR VPWR _08275_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15134_ net479 VGND VGND VPWR VPWR _07233_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19942_ net202 net183 VGND VGND VPWR VPWR _11813_ sky130_fd_sc_hd__nand2_1
X_15065_ net520 net489 VGND VGND VPWR VPWR _07164_ sky130_fd_sc_hd__nand2_2
XFILLER_0_50_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14016_ _06096_ _06227_ _06228_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__o21a_1
X_19873_ _11519_ _11718_ _11732_ net237 VGND VGND VPWR VPWR _11749_ sky130_fd_sc_hd__o31a_1
X_18824_ net362 _10797_ _10798_ _10799_ VGND VGND VPWR VPWR _10800_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_156_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18755_ _10629_ _10653_ _10652_ VGND VGND VPWR VPWR _10732_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15967_ _08010_ _08061_ VGND VGND VPWR VPWR _08062_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17706_ _09360_ _09691_ _09692_ VGND VGND VPWR VPWR _09693_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_175_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14918_ spi0.data_packed\[34\] top0.kid\[2\] _07075_ VGND VGND VPWR VPWR _07080_
+ sky130_fd_sc_hd__mux2_1
X_18686_ _10662_ _10663_ VGND VGND VPWR VPWR _10664_ sky130_fd_sc_hd__xor2_1
X_15898_ _07993_ _07705_ VGND VGND VPWR VPWR _07994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17637_ _09620_ _09623_ VGND VGND VPWR VPWR _09624_ sky130_fd_sc_hd__xnor2_2
X_14849_ spi0.data_packed\[65\] top0.kpd\[1\] _07042_ VGND VGND VPWR VPWR _07044_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17568_ _09540_ _09541_ VGND VGND VPWR VPWR _09555_ sky130_fd_sc_hd__xor2_2
XFILLER_0_86_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19307_ top0.pid_d.prev_error\[12\] top0.pid_d.curr_error\[12\] VGND VGND VPWR VPWR
+ _11248_ sky130_fd_sc_hd__nand2_1
X_16519_ _08489_ _08606_ _08546_ VGND VGND VPWR VPWR _08607_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_46_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17499_ _09482_ _09485_ VGND VGND VPWR VPWR _09486_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19238_ _11183_ _11175_ _11184_ VGND VGND VPWR VPWR _11185_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19169_ _11122_ VGND VGND VPWR VPWR _11123_ sky130_fd_sc_hd__buf_2
XFILLER_0_121_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21200_ _13018_ _13043_ VGND VGND VPWR VPWR _13044_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22180_ _01724_ _01722_ _01727_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21131_ _11673_ _12785_ VGND VGND VPWR VPWR _12976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout403 top0.pid_d.mult0.a\[6\] VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkbuf_4
X_21062_ _11593_ _12904_ _12906_ _12847_ _12907_ VGND VGND VPWR VPWR _12908_ sky130_fd_sc_hd__o221a_1
Xfanout414 top0.pid_d.mult0.a\[4\] VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__buf_2
Xfanout425 net427 VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__clkbuf_4
Xfanout436 top0.pid_d.state\[2\] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__buf_2
X_20013_ _11426_ _11875_ _11878_ VGND VGND VPWR VPWR _11879_ sky130_fd_sc_hd__and3_1
Xfanout447 net448 VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__clkbuf_4
X_25870_ net1024 top0.matmul0.beta_pass\[8\] VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__nor2_1
Xfanout458 net459 VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__clkbuf_4
Xfanout469 net470 VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__buf_2
X_24821_ _03741_ _03742_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24752_ _04020_ _04025_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__or2_1
X_21964_ _01320_ _01524_ _01525_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23703_ net570 net575 top0.matmul0.matmul_stage_inst.f\[9\] VGND VGND VPWR VPWR _03061_
+ sky130_fd_sc_hd__o21a_4
X_20915_ _12761_ _12762_ net241 VGND VGND VPWR VPWR _12763_ sky130_fd_sc_hd__and3b_1
X_24683_ _04036_ _03918_ _03915_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__o21a_1
XFILLER_0_194_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21895_ _01455_ _01456_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__xnor2_2
X_23634_ _02985_ _02987_ _02989_ _02991_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__o22a_1
X_26422_ clknet_leaf_58_clk_sys _00063_ net653 VGND VGND VPWR VPWR top0.kpq\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_194_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20846_ net296 _12690_ _12694_ VGND VGND VPWR VPWR _12695_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout10 _12744_ VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__clkbuf_4
Xfanout21 net22 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_154_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout32 top0.periodTop_r\[13\] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_4
XFILLER_0_92_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout43 top0.periodTop_r\[8\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_4
X_23565_ _02949_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26353_ _05408_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__clkbuf_1
Xfanout54 top0.periodTop_r\[4\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_4
X_20777_ _12624_ _12625_ VGND VGND VPWR VPWR _12626_ sky130_fd_sc_hd__nand2_1
Xfanout65 net67 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout76 top0.matmul0.alpha_pass\[5\] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_4
X_25304_ _04612_ _04649_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22516_ _01980_ _01967_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26284_ net946 spi0.data_packed\[41\] net688 VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__mux2_1
Xfanout87 net89 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_2
Xfanout98 top0.cordic0.vec\[1\]\[14\] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23496_ net718 top0.matmul0.cos\[3\] _02904_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25235_ _04579_ _04581_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22447_ _01944_ _01891_ _01737_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_51_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25166_ _04508_ _04513_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__xnor2_1
X_22378_ net91 _01230_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__nand2_1
X_24117_ _03474_ _03161_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21329_ _13001_ _13170_ VGND VGND VPWR VPWR _13171_ sky130_fd_sc_hd__or2_1
X_25097_ _04443_ _04445_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24048_ _03404_ _03405_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__nor2_1
XFILLER_0_202_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16870_ top0.matmul0.beta_pass\[4\] _08932_ VGND VGND VPWR VPWR _08933_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15821_ _07915_ _07916_ VGND VGND VPWR VPWR _07917_ sky130_fd_sc_hd__xor2_2
XFILLER_0_99_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25999_ top0.pid_q.out\[9\] _05198_ _05199_ spi0.data_packed\[57\] VGND VGND VPWR
+ VPWR _05200_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18540_ _10255_ _10518_ _10454_ _10449_ VGND VGND VPWR VPWR _10519_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15752_ net465 net518 VGND VGND VPWR VPWR _07849_ sky130_fd_sc_hd__nand2_1
X_14703_ _06863_ _06906_ VGND VGND VPWR VPWR _06907_ sky130_fd_sc_hd__xnor2_4
X_18471_ net393 net315 VGND VGND VPWR VPWR _10451_ sky130_fd_sc_hd__nand2_1
X_15683_ net506 VGND VGND VPWR VPWR _07781_ sky130_fd_sc_hd__inv_2
X_17422_ net330 net422 VGND VGND VPWR VPWR _09409_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14634_ _06760_ _06762_ _06838_ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17353_ net418 net344 VGND VGND VPWR VPWR _09340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14565_ _06767_ _06770_ VGND VGND VPWR VPWR _06771_ sky130_fd_sc_hd__xnor2_2
X_16304_ _08394_ VGND VGND VPWR VPWR _08395_ sky130_fd_sc_hd__inv_2
X_13516_ _05725_ _05728_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__xnor2_1
X_17284_ _09280_ _09276_ top0.matmul0.matmul_stage_inst.mult1\[5\] VGND VGND VPWR
+ VPWR _09281_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14496_ _06701_ _06702_ VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19023_ _10968_ _10969_ _10995_ VGND VGND VPWR VPWR _10996_ sky130_fd_sc_hd__o21ai_2
X_16235_ _08324_ _08245_ _08325_ VGND VGND VPWR VPWR _08326_ sky130_fd_sc_hd__a21o_1
X_13447_ _05658_ _05659_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13378_ net57 net54 _05586_ _05588_ _05590_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__a41o_1
X_16166_ _08256_ _08257_ VGND VGND VPWR VPWR _08258_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15117_ _07211_ _07212_ _07214_ VGND VGND VPWR VPWR _07216_ sky130_fd_sc_hd__a21o_1
XFILLER_0_142_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16097_ _08093_ _08095_ _08094_ VGND VGND VPWR VPWR _08190_ sky130_fd_sc_hd__o21a_1
XFILLER_0_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19925_ net194 _11576_ VGND VGND VPWR VPWR _11797_ sky130_fd_sc_hd__nor2_1
X_15048_ net514 net494 VGND VGND VPWR VPWR _07147_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19856_ _11729_ _11732_ VGND VGND VPWR VPWR _11733_ sky130_fd_sc_hd__xor2_2
XFILLER_0_177_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_3__f_clk_mosi clknet_0_clk_mosi VGND VGND VPWR VPWR clknet_3_3__leaf_clk_mosi
+ sky130_fd_sc_hd__clkbuf_16
X_18807_ _10208_ _10778_ _10782_ net316 VGND VGND VPWR VPWR _10783_ sky130_fd_sc_hd__a22o_1
X_19787_ _11664_ _11668_ VGND VGND VPWR VPWR _11669_ sky130_fd_sc_hd__xor2_1
X_16999_ top0.pid_q.prev_error\[12\] top0.pid_q.curr_error\[12\] _09052_ VGND VGND
+ VPWR VPWR _09053_ sky130_fd_sc_hd__a21o_1
XFILLER_0_183_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18738_ _10709_ _10714_ VGND VGND VPWR VPWR _10715_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18669_ _10642_ _10645_ VGND VGND VPWR VPWR _10647_ sky130_fd_sc_hd__nand2_1
X_20700_ _12547_ _12548_ VGND VGND VPWR VPWR _12549_ sky130_fd_sc_hd__xnor2_1
X_21680_ _01231_ _01241_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__xor2_2
XFILLER_0_47_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20631_ _12453_ _12479_ VGND VGND VPWR VPWR _12480_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_178_Right_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23350_ _01408_ _02793_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20562_ _12115_ _12410_ VGND VGND VPWR VPWR _12411_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22301_ _01818_ _01860_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_172_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23281_ _11572_ _02650_ _02657_ _11574_ _11576_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__a221o_1
XFILLER_0_171_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20493_ _12245_ _12247_ VGND VGND VPWR VPWR _12342_ sky130_fd_sc_hd__xor2_2
XFILLER_0_144_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25020_ _04279_ _04281_ _04369_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22232_ _01774_ _01792_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22163_ net105 net90 _01235_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21114_ _12957_ _12959_ _12804_ VGND VGND VPWR VPWR _12960_ sky130_fd_sc_hd__mux2_1
X_26971_ clknet_leaf_27_clk_sys _00588_ net621 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[3\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout200 top0.cordic0.gm0.iter\[0\] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_2
X_22094_ _01635_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout211 top0.cordic0.domain\[1\] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__buf_2
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout222 net224 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25922_ _05110_ _05127_ _05135_ _05136_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__a31o_1
X_21045_ _12835_ _12863_ VGND VGND VPWR VPWR _12891_ sky130_fd_sc_hd__and2b_1
Xfanout233 top0.cordic0.vec\[0\]\[14\] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_2
Xfanout244 net245 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__buf_4
Xfanout255 net256 VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout266 net268 VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_201_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout277 net278 VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__buf_2
X_25853_ top0.matmul0.alpha_pass\[6\] top0.matmul0.beta_pass\[6\] VGND VGND VPWR VPWR
+ _05074_ sky130_fd_sc_hd__nor2_1
Xfanout288 net293 VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkbuf_2
Xfanout299 net301 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24804_ _04066_ _04152_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25784_ top0.pid_d.out_valid _12030_ _05015_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__o21ai_1
X_22996_ net169 _02501_ _02502_ _02500_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24735_ _04078_ _04087_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__xor2_4
XFILLER_0_119_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21947_ _01199_ _01508_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24666_ _03874_ _04018_ _04019_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__a21oi_2
X_21878_ _01437_ _01439_ net166 VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26405_ clknet_leaf_79_clk_sys _00046_ net632 VGND VGND VPWR VPWR top0.kpd\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_23617_ _02975_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__clkbuf_1
X_20829_ _12223_ _12226_ _12217_ VGND VGND VPWR VPWR _12678_ sky130_fd_sc_hd__a21o_1
XFILLER_0_166_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24597_ _03834_ _03951_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14350_ _06513_ _06528_ VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26336_ spi0.data_packed\[66\] spi0.data_packed\[67\] net690 VGND VGND VPWR VPWR
+ _05400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23548_ _02940_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__clkbuf_1
X_13301_ net40 _05484_ _05486_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__and3_1
X_14281_ _06489_ _06490_ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26267_ _05365_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23479_ _05460_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__buf_4
XFILLER_0_150_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16020_ _08013_ _08015_ _08014_ VGND VGND VPWR VPWR _08114_ sky130_fd_sc_hd__o21a_1
X_13232_ net547 _05441_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__and2_1
X_25218_ _04555_ _04564_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26198_ _05330_ VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25149_ _04428_ _04430_ _04429_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17971_ _09934_ _09956_ VGND VGND VPWR VPWR _09957_ sky130_fd_sc_hd__nor2_1
X_19710_ net188 net82 VGND VGND VPWR VPWR _11595_ sky130_fd_sc_hd__nand2_1
X_16922_ net546 _08974_ _08981_ _08882_ VGND VGND VPWR VPWR _08982_ sky130_fd_sc_hd__a211o_1
X_19641_ _11438_ _11528_ VGND VGND VPWR VPWR _11529_ sky130_fd_sc_hd__nand2_1
X_16853_ _08915_ _08916_ _05601_ VGND VGND VPWR VPWR _08917_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15804_ top0.pid_q.out\[2\] top0.pid_q.curr_int\[2\] VGND VGND VPWR VPWR _07900_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19572_ top0.cordic0.slte0.opA\[4\] top0.cordic0.slte0.opB\[4\] VGND VGND VPWR VPWR
+ _11461_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16784_ top0.kiq\[2\] _08863_ _08861_ VGND VGND VPWR VPWR _08865_ sky130_fd_sc_hd__and3_1
X_13996_ _06205_ _06208_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_137_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18523_ _10492_ _10502_ VGND VGND VPWR VPWR _10503_ sky130_fd_sc_hd__xor2_1
X_15735_ _07826_ _07831_ VGND VGND VPWR VPWR _07832_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_87_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18454_ _10421_ _10433_ VGND VGND VPWR VPWR _10434_ sky130_fd_sc_hd__nand2_1
X_15666_ _07630_ _07634_ _07632_ VGND VGND VPWR VPWR _07764_ sky130_fd_sc_hd__a21o_1
X_17405_ _09350_ _09390_ VGND VGND VPWR VPWR _09392_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14617_ _06782_ _06775_ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__or2b_1
XFILLER_0_200_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18385_ net331 net376 VGND VGND VPWR VPWR _10366_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15597_ _07694_ _07695_ VGND VGND VPWR VPWR _07696_ sky130_fd_sc_hd__or2_1
XFILLER_0_173_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17336_ top0.matmul0.beta_pass\[13\] _09325_ net563 VGND VGND VPWR VPWR _09326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14548_ net44 _06351_ _06701_ _06702_ VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17267_ _09265_ _09266_ VGND VGND VPWR VPWR _09267_ sky130_fd_sc_hd__xnor2_1
X_14479_ _06608_ _06609_ _06672_ VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19006_ _10976_ _10978_ VGND VGND VPWR VPWR _10980_ sky130_fd_sc_hd__nand2_1
X_16218_ _08305_ _08309_ VGND VGND VPWR VPWR _08310_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17198_ top0.pid_q.prev_int\[9\] VGND VGND VPWR VPWR _09207_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16149_ top0.pid_q.out\[6\] _07705_ _08241_ net545 VGND VGND VPWR VPWR _08242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19908_ _11431_ _11781_ net175 VGND VGND VPWR VPWR _11782_ sky130_fd_sc_hd__o21ai_1
Xhold19 top0.kpq\[6\] VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19839_ _11415_ _11714_ _11716_ _11654_ _11675_ VGND VGND VPWR VPWR _11717_ sky130_fd_sc_hd__o221a_2
XFILLER_0_190_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22850_ _02360_ top0.svm0.tA\[9\] _02368_ _02369_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_166_Left_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21801_ _01335_ _01353_ _01348_ _01362_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__a211oi_2
X_22781_ _02296_ _02304_ VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24520_ _03076_ _03077_ _03717_ _03718_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__o22a_1
X_21732_ net152 net147 VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24451_ _03805_ _03806_ _03088_ _03089_ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__a211o_2
X_21663_ _01066_ _01224_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_136_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20614_ _12445_ _12462_ VGND VGND VPWR VPWR _12463_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23402_ _01065_ _02810_ _02839_ _02840_ _02841_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__a311o_1
X_24382_ _03186_ _03187_ _03188_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__a21oi_1
X_27170_ clknet_leaf_12_clk_sys _00784_ net618 VGND VGND VPWR VPWR top0.periodTop_r\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_21594_ net164 _01093_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23333_ _11526_ _02777_ net176 VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__o21a_1
X_26121_ spi0.data_packed\[18\] _05279_ _05280_ top0.currT_r\[2\] VGND VGND VPWR VPWR
+ _00799_ sky130_fd_sc_hd__a22o_1
X_20545_ _12279_ _12266_ VGND VGND VPWR VPWR _12394_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_175_Left_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23264_ net244 net243 net237 net233 net204 net196 VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__mux4_2
X_26052_ top0.pid_d.out\[5\] _05232_ _05233_ spi0.data_packed\[69\] VGND VGND VPWR
+ VPWR _05241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20476_ _12261_ _12324_ VGND VGND VPWR VPWR _12325_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25003_ _04273_ _04274_ _04271_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__a21bo_1
X_22215_ net90 net96 VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__nor2b_1
X_23195_ _05719_ _07028_ _02648_ net804 VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__a22o_1
X_22146_ net132 _01135_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__nand2_1
X_26954_ clknet_leaf_16_clk_sys _00571_ net613 VGND VGND VPWR VPWR top0.matmul0.b\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_22077_ _01193_ _01184_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__xnor2_1
X_25905_ _05102_ _05110_ _05121_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__nand3_1
X_21028_ _12865_ _12874_ VGND VGND VPWR VPWR _12875_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_22_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26885_ clknet_leaf_38_clk_sys _00502_ net678 VGND VGND VPWR VPWR top0.svm0.tB\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_184_Left_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25836_ top0.matmul0.alpha_pass\[4\] top0.matmul0.beta_pass\[4\] VGND VGND VPWR VPWR
+ _05059_ sky130_fd_sc_hd__or2_2
X_13850_ _06056_ _06059_ _06062_ net68 VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_199_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_202_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13781_ _05973_ _05977_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__xor2_1
X_25767_ _05004_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__clkbuf_1
X_22979_ top0.svm0.delta\[8\] _02487_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_201_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15520_ net495 net505 VGND VGND VPWR VPWR _07619_ sky130_fd_sc_hd__nand2_1
X_24718_ _03985_ _03986_ _04070_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__o21a_2
XFILLER_0_84_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25698_ net69 top0.matmul0.sin\[0\] _04896_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15451_ net518 net475 VGND VGND VPWR VPWR _07550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24649_ _03864_ _03865_ _03866_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__a21oi_2
X_14402_ _06557_ _06610_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__xor2_2
XFILLER_0_139_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18170_ _10149_ _10153_ VGND VGND VPWR VPWR _10154_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15382_ _07457_ _07480_ VGND VGND VPWR VPWR _07481_ sky130_fd_sc_hd__xor2_1
XFILLER_0_182_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_193_Left_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17121_ net15 _09134_ VGND VGND VPWR VPWR _09140_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14333_ _06476_ _06542_ VGND VGND VPWR VPWR _06543_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26319_ _05391_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27299_ clknet_3_1__leaf_clk_mosi _00913_ VGND VGND VPWR VPWR spi0.opcode\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17052_ _09101_ VGND VGND VPWR VPWR _09102_ sky130_fd_sc_hd__clkbuf_4
X_14264_ _06387_ _06471_ _06470_ VGND VGND VPWR VPWR _06474_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16003_ _08093_ _08096_ VGND VGND VPWR VPWR _08097_ sky130_fd_sc_hd__xnor2_2
X_13215_ spi0.cs_sync\[2\] _05428_ _05429_ spi0.cs_sync\[1\] VGND VGND VPWR VPWR _05440_
+ sky130_fd_sc_hd__or4b_1
X_14195_ _06402_ _06405_ VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_93_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_93_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_104_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17954_ _09863_ _09864_ _09862_ VGND VGND VPWR VPWR _09940_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16905_ top0.pid_q.prev_error\[6\] top0.pid_q.curr_error\[6\] VGND VGND VPWR VPWR
+ _08966_ sky130_fd_sc_hd__xor2_1
X_17885_ _09870_ _09871_ VGND VGND VPWR VPWR _09872_ sky130_fd_sc_hd__xor2_2
XFILLER_0_174_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16836_ top0.matmul0.beta_pass\[1\] top0.currT_r\[1\] VGND VGND VPWR VPWR _08901_
+ sky130_fd_sc_hd__or2b_1
X_19624_ _11512_ VGND VGND VPWR VPWR _11513_ sky130_fd_sc_hd__clkbuf_4
X_19555_ net81 VGND VGND VPWR VPWR _11444_ sky130_fd_sc_hd__inv_2
X_16767_ _05448_ _07700_ _08849_ _08850_ VGND VGND VPWR VPWR _08851_ sky130_fd_sc_hd__a31o_1
XFILLER_0_189_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13979_ net56 _05663_ _05664_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__and3_1
X_18506_ _10481_ _10485_ VGND VGND VPWR VPWR _10486_ sky130_fd_sc_hd__xor2_1
X_15718_ net477 net509 VGND VGND VPWR VPWR _07815_ sky130_fd_sc_hd__nand2_1
X_19486_ _11376_ _11379_ VGND VGND VPWR VPWR _11380_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16698_ _08747_ _08782_ VGND VGND VPWR VPWR _08783_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18437_ _10346_ _10417_ VGND VGND VPWR VPWR _10418_ sky130_fd_sc_hd__xnor2_1
X_15649_ _07638_ _07639_ _07746_ VGND VGND VPWR VPWR _07747_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_186_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18368_ net397 _10203_ _09363_ VGND VGND VPWR VPWR _10349_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17319_ _09310_ _09306_ top0.matmul0.matmul_stage_inst.mult1\[10\] VGND VGND VPWR
+ VPWR _09311_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_71_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18299_ _10279_ _10280_ VGND VGND VPWR VPWR _10281_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20330_ _12176_ _12178_ VGND VGND VPWR VPWR _12179_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20261_ _11408_ _12067_ _12108_ _12109_ _11571_ VGND VGND VPWR VPWR _12110_ sky130_fd_sc_hd__a32oi_1
XFILLER_0_3_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22000_ _01290_ _01293_ _01295_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_109_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20192_ _12038_ _12040_ VGND VGND VPWR VPWR _12041_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23951_ _03007_ _03114_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__nor2_2
X_22902_ top0.svm0.tC\[7\] _02418_ VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__and2_1
X_26670_ clknet_leaf_82_clk_sys _00287_ net647 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_23882_ _03022_ _03023_ _02988_ _02990_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__o22a_1
X_25621_ net742 _04896_ _04887_ _04902_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__o22a_1
X_22833_ _02352_ top0.svm0.tA\[1\] VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25552_ net943 top0.matmul0.matmul_stage_inst.f\[15\] _04856_ VGND VGND VPWR VPWR
+ _04863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22764_ top0.pid_q.prev_int\[8\] _02292_ _02295_ net924 VGND VGND VPWR VPWR _00427_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24503_ _03663_ _03676_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__and2_1
X_21715_ _01262_ _01264_ _01276_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__o21a_1
X_25483_ _04661_ _04756_ _04822_ _04823_ _04825_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__a311o_1
X_22695_ _01643_ _01248_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27222_ clknet_3_4__leaf_clk_mosi _00836_ VGND VGND VPWR VPWR spi0.data_packed\[8\]
+ sky130_fd_sc_hd__dfxtp_2
X_24434_ _02989_ _02991_ _03069_ _03071_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__o22a_1
X_21646_ net150 net128 VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_118_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27153_ clknet_leaf_9_clk_sys _00767_ net594 VGND VGND VPWR VPWR top0.a_in_matmul\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_24365_ _03717_ _03718_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__or2_2
XFILLER_0_145_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21577_ net139 net131 VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_23_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26104_ net782 _05276_ _05278_ net58 VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__a22o_1
X_20528_ _12369_ _12376_ VGND VGND VPWR VPWR _12377_ sky130_fd_sc_hd__xnor2_2
X_23316_ _02707_ _02759_ _02761_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__a21o_1
X_24296_ _03624_ _03625_ _03622_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__a21o_1
X_27084_ clknet_leaf_8_clk_sys _00701_ net592 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26035_ _05227_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__clkbuf_1
X_20459_ net295 net275 VGND VGND VPWR VPWR _12308_ sky130_fd_sc_hd__or2_1
X_23247_ _11857_ _02696_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23178_ _05719_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22129_ _01215_ _01219_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26937_ clknet_leaf_9_clk_sys _00554_ net595 VGND VGND VPWR VPWR top0.matmul0.a\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14951_ _07041_ VGND VGND VPWR VPWR _07097_ sky130_fd_sc_hd__buf_4
X_13902_ _06113_ _06114_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__xor2_1
X_17670_ net409 net333 VGND VGND VPWR VPWR _09657_ sky130_fd_sc_hd__nand2_1
X_26868_ clknet_leaf_40_clk_sys _00485_ net677 VGND VGND VPWR VPWR top0.svm0.tA\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14882_ spi0.data_packed\[49\] top0.kpq\[1\] _07053_ VGND VGND VPWR VPWR _07061_
+ sky130_fd_sc_hd__mux2_1
X_16621_ _08698_ _08706_ VGND VGND VPWR VPWR _08707_ sky130_fd_sc_hd__xnor2_1
X_13833_ _05489_ _05491_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__nand2_2
X_25819_ _05033_ _05039_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__nand2_1
X_26799_ clknet_leaf_102_clk_sys _00416_ net589 VGND VGND VPWR VPWR top0.cordic0.gm0.iter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_6__f_clk_sys clknet_0_clk_sys VGND VGND VPWR VPWR clknet_3_6__leaf_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19340_ _05442_ _11276_ VGND VGND VPWR VPWR _11277_ sky130_fd_sc_hd__and2_1
XFILLER_0_202_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16552_ net452 net501 VGND VGND VPWR VPWR _08639_ sky130_fd_sc_hd__nand2_1
X_13764_ _05974_ _05975_ _05976_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15503_ _07255_ _07601_ _07298_ VGND VGND VPWR VPWR _07602_ sky130_fd_sc_hd__o21ba_1
X_19271_ _11214_ _11205_ top0.pid_d.prev_error\[9\] VGND VGND VPWR VPWR _11215_ sky130_fd_sc_hd__o21ba_1
X_16483_ _08497_ _08498_ _08570_ VGND VGND VPWR VPWR _08571_ sky130_fd_sc_hd__a21boi_2
X_13695_ _05875_ _05878_ _05907_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_183_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18222_ net405 _09353_ _09363_ VGND VGND VPWR VPWR _10205_ sky130_fd_sc_hd__and3_1
X_15434_ _07266_ _07280_ VGND VGND VPWR VPWR _07533_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18153_ _10044_ _10045_ _10136_ VGND VGND VPWR VPWR _10137_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15365_ _07442_ _07463_ VGND VGND VPWR VPWR _07464_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17104_ net826 _09114_ _09128_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14316_ _06523_ _06525_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18084_ top0.pid_d.curr_int\[2\] _09981_ _09982_ top0.pid_d.out\[2\] VGND VGND VPWR
+ VPWR _10068_ sky130_fd_sc_hd__a31o_1
X_15296_ _07393_ _07394_ VGND VGND VPWR VPWR _07395_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold308 top0.cordic0.cos\[6\] VGND VGND VPWR VPWR net1008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17035_ _09084_ _09086_ VGND VGND VPWR VPWR _09087_ sky130_fd_sc_hd__nand2_1
X_14247_ _06453_ _06457_ VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__xor2_1
XFILLER_0_150_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14178_ _06358_ _06366_ _06388_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_194_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18986_ _10954_ _10959_ VGND VGND VPWR VPWR _10960_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17937_ _09919_ _09922_ VGND VGND VPWR VPWR _09923_ sky130_fd_sc_hd__xnor2_2
X_17868_ _09851_ _09854_ VGND VGND VPWR VPWR _09855_ sky130_fd_sc_hd__xor2_1
XFILLER_0_139_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19607_ _11486_ _11490_ VGND VGND VPWR VPWR _11496_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16819_ top0.pid_q.prev_error\[0\] top0.pid_q.curr_error\[0\] VGND VGND VPWR VPWR
+ _08886_ sky130_fd_sc_hd__xor2_1
X_17799_ _09666_ _09785_ VGND VGND VPWR VPWR _09786_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_191_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19538_ net186 net190 _11427_ VGND VGND VPWR VPWR _11428_ sky130_fd_sc_hd__or3_2
XFILLER_0_88_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19469_ _10834_ _11364_ VGND VGND VPWR VPWR _11365_ sky130_fd_sc_hd__nor2_1
X_21500_ net97 VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22480_ _01953_ _01976_ _01971_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21431_ _00996_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24150_ _03506_ _03507_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21362_ _00929_ _13182_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23101_ top0.svm0.delta\[1\] net555 _02443_ _02598_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__o211a_1
X_20313_ _12086_ _12088_ _12091_ _12097_ VGND VGND VPWR VPWR _12162_ sky130_fd_sc_hd__o2bb2a_1
X_24081_ _03346_ _03348_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__nand2_1
X_21293_ _13112_ _13135_ VGND VGND VPWR VPWR _13136_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_47_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23032_ top0.svm0.counter\[15\] _02531_ _02532_ _02533_ VGND VGND VPWR VPWR _02534_
+ sky130_fd_sc_hd__a22o_1
X_20244_ _12086_ _12088_ _12091_ VGND VGND VPWR VPWR _12093_ sky130_fd_sc_hd__a21o_1
X_20175_ net209 _12008_ _12026_ VGND VGND VPWR VPWR _12027_ sky130_fd_sc_hd__mux2_1
X_24983_ _04315_ _04316_ _04332_ _04170_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26722_ clknet_leaf_78_clk_sys _00339_ net633 VGND VGND VPWR VPWR top0.pid_d.curr_int\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_23934_ _03270_ _03271_ _03287_ _03290_ _03291_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__o311a_1
X_26653_ clknet_leaf_75_clk_sys _00270_ net636 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_23865_ _03213_ _03222_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_168_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25604_ net836 _00000_ _04893_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_41_clk_sys clknet_3_7__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_41_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_196_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22816_ top0.svm0.counter\[9\] top0.svm0.tA\[9\] VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__or2_1
X_26584_ clknet_leaf_53_clk_sys _00207_ net674 VGND VGND VPWR VPWR top0.pid_q.prev_error\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_23796_ _03144_ _03153_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25535_ top0.matmul0.b\[7\] top0.matmul0.matmul_stage_inst.f\[7\] _04846_ VGND VGND
+ VPWR VPWR _04854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22747_ net186 _11558_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25466_ _04808_ _04750_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__and2_1
XFILLER_0_176_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13480_ _05681_ _05692_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22678_ _02186_ _02227_ _02229_ net210 VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__o211a_1
XFILLER_0_192_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27205_ clknet_leaf_92_clk_sys _00819_ net599 VGND VGND VPWR VPWR top0.cordic0.slte0.opB\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24417_ _03767_ _03772_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21629_ _01062_ _01067_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__or2_1
X_25397_ _04685_ _04688_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27136_ clknet_leaf_13_clk_sys _00750_ net616 VGND VGND VPWR VPWR top0.b_in_matmul\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_15150_ net521 net480 VGND VGND VPWR VPWR _07249_ sky130_fd_sc_hd__nand2_1
X_24348_ _03210_ _03211_ _03209_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14101_ _06206_ _06207_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__and2_1
X_27067_ clknet_leaf_2_clk_sys _00684_ net582 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.c\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15081_ net540 _07178_ _07179_ net464 VGND VGND VPWR VPWR _07180_ sky130_fd_sc_hd__o22a_1
XFILLER_0_200_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24279_ _03626_ _03630_ _03631_ VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14032_ net64 _06135_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__nand2_1
X_26018_ top0.b_in_matmul\[13\] _05214_ _05196_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18840_ _10809_ _10815_ VGND VGND VPWR VPWR _10816_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18771_ _10746_ _10744_ VGND VGND VPWR VPWR _10748_ sky130_fd_sc_hd__or2b_1
XFILLER_0_100_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15983_ top0.pid_q.curr_int\[3\] _07901_ _08077_ VGND VGND VPWR VPWR _08078_ sky130_fd_sc_hd__o21ba_1
X_17722_ net391 net381 net357 VGND VGND VPWR VPWR _09709_ sky130_fd_sc_hd__o21ai_1
X_14934_ _07088_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__clkbuf_1
X_17653_ _09637_ _09638_ _09639_ net378 VGND VGND VPWR VPWR _09640_ sky130_fd_sc_hd__a2bb2o_1
X_14865_ spi0.data_packed\[73\] top0.kpd\[9\] _07042_ VGND VGND VPWR VPWR _07052_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16604_ _08687_ _08688_ _08689_ _08677_ VGND VGND VPWR VPWR _08690_ sky130_fd_sc_hd__o211ai_4
X_13816_ _06027_ _06028_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__xnor2_2
X_17584_ net412 _09569_ _09570_ net415 VGND VGND VPWR VPWR _09571_ sky130_fd_sc_hd__a2bb2o_1
X_14796_ _06949_ _06993_ _06994_ _06935_ VGND VGND VPWR VPWR _06997_ sky130_fd_sc_hd__a22o_1
X_19323_ top0.matmul0.alpha_pass\[14\] _11245_ VGND VGND VPWR VPWR _11263_ sky130_fd_sc_hd__and2_1
XFILLER_0_161_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16535_ _08621_ _07703_ VGND VGND VPWR VPWR _08622_ sky130_fd_sc_hd__nor2_1
X_13747_ net62 _05472_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19254_ net438 _11198_ _11199_ VGND VGND VPWR VPWR _11200_ sky130_fd_sc_hd__and3_1
X_16466_ net455 net500 VGND VGND VPWR VPWR _08554_ sky130_fd_sc_hd__nand2_2
XFILLER_0_39_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13678_ _05869_ _05870_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__xor2_2
XFILLER_0_73_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18205_ net345 net370 VGND VGND VPWR VPWR _10188_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15417_ _07460_ _07465_ _07514_ _07515_ VGND VGND VPWR VPWR _07516_ sky130_fd_sc_hd__a211o_1
XFILLER_0_183_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19185_ _11135_ _11136_ VGND VGND VPWR VPWR _11137_ sky130_fd_sc_hd__or2_1
XFILLER_0_171_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16397_ _08406_ _08484_ _08485_ VGND VGND VPWR VPWR _08486_ sky130_fd_sc_hd__o21ai_2
X_18136_ _10025_ _10027_ _10026_ VGND VGND VPWR VPWR _10120_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15348_ net533 _07402_ VGND VGND VPWR VPWR _07447_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold105 top0.matmul0.matmul_stage_inst.c\[9\] VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__dlygate4sd3_1
X_18067_ _10050_ _10051_ VGND VGND VPWR VPWR _10052_ sky130_fd_sc_hd__nand2_1
Xhold116 _00132_ VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__dlygate4sd3_1
X_15279_ _07328_ _07334_ _07337_ _07342_ VGND VGND VPWR VPWR _07378_ sky130_fd_sc_hd__or4_1
XFILLER_0_110_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold127 top0.kpq\[8\] VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 top0.svm0.tB\[14\] VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 top0.pid_q.prev_error\[5\] VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ top0.pid_q.prev_error\[13\] top0.pid_q.curr_error\[13\] VGND VGND VPWR VPWR
+ _09071_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout607 net608 VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__clkbuf_4
Xfanout618 net619 VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__clkbuf_4
Xfanout629 net630 VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18969_ net376 net308 VGND VGND VPWR VPWR _10943_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21980_ _01468_ _01479_ _01539_ _01536_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__o2bb2a_1
X_20931_ _12777_ _12778_ VGND VGND VPWR VPWR _12779_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23650_ _03006_ _03007_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__nor2_2
X_20862_ _12701_ _12709_ _12710_ VGND VGND VPWR VPWR _12711_ sky130_fd_sc_hd__nand3_1
XFILLER_0_113_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22601_ _01213_ _01063_ net92 VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__or3_1
XFILLER_0_147_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23581_ _02957_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20793_ _12598_ _12641_ VGND VGND VPWR VPWR _12642_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_165_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25320_ _04521_ _04643_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22532_ _02003_ _02085_ _02087_ _02007_ net210 VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25251_ _04597_ _04527_ _04455_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22463_ net88 _01775_ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__xnor2_2
X_24202_ _03315_ _03323_ _03217_ _03337_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__a22o_1
X_21414_ _00979_ _00980_ VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__nand2_1
X_25182_ _04455_ _04526_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__nand2_1
X_22394_ _01921_ _01928_ _01916_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__a21o_1
X_24133_ _03036_ _03037_ _03027_ _03028_ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21345_ _13159_ _13186_ VGND VGND VPWR VPWR _13187_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24064_ _03413_ _03414_ _03420_ _03421_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__a211o_1
X_21276_ _13031_ _13113_ VGND VGND VPWR VPWR _13119_ sky130_fd_sc_hd__and2b_1
XFILLER_0_60_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23015_ net172 _02317_ _02518_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__o21ai_1
X_20227_ _11758_ _12074_ _12075_ VGND VGND VPWR VPWR _12076_ sky130_fd_sc_hd__nor3_1
XFILLER_0_200_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20158_ _12009_ net208 VGND VGND VPWR VPWR _12010_ sky130_fd_sc_hd__or2_1
XFILLER_0_200_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24966_ _04172_ _04178_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__and2_1
X_20089_ net194 net203 _11730_ _11947_ _11948_ VGND VGND VPWR VPWR _11949_ sky130_fd_sc_hd__a41o_1
X_26705_ clknet_leaf_84_clk_sys net904 net641 VGND VGND VPWR VPWR top0.pid_d.prev_error\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_23917_ _03273_ _03274_ _03272_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__a21o_1
XFILLER_0_197_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24897_ _03962_ _04059_ _04060_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__o21ai_1
X_14650_ _06755_ _06756_ _06753_ VGND VGND VPWR VPWR _06855_ sky130_fd_sc_hd__a21o_1
X_26636_ clknet_leaf_81_clk_sys _00253_ net636 VGND VGND VPWR VPWR top0.pid_d.out\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_23848_ _03199_ _03205_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__xor2_2
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13601_ _05811_ _05812_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14581_ _06714_ _06725_ VGND VGND VPWR VPWR _06787_ sky130_fd_sc_hd__or2_1
X_26567_ clknet_leaf_52_clk_sys _00190_ net672 VGND VGND VPWR VPWR top0.pid_q.curr_error\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_23779_ _03132_ _03133_ _03136_ _03087_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__a22o_1
X_16320_ _08316_ _08330_ _08394_ VGND VGND VPWR VPWR _08410_ sky130_fd_sc_hd__a21o_1
X_25518_ top0.matmul0.matmul_stage_inst.mult1\[15\] _04827_ _03148_ VGND VGND VPWR
+ VPWR _04845_ sky130_fd_sc_hd__mux2_1
X_13532_ _05672_ _05661_ _05669_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_82_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26498_ clknet_leaf_73_clk_sys _00121_ net655 VGND VGND VPWR VPWR top0.pid_d.prev_int\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16251_ net476 _08141_ _08341_ VGND VGND VPWR VPWR _08342_ sky130_fd_sc_hd__a21o_1
X_25449_ _04723_ _04724_ _04722_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__a21bo_1
X_13463_ _05653_ _05675_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15202_ _07251_ _07300_ VGND VGND VPWR VPWR _07301_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16182_ _08272_ _08273_ VGND VGND VPWR VPWR _08274_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13394_ net63 VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__inv_2
X_27119_ clknet_leaf_33_clk_sys _00733_ net665 VGND VGND VPWR VPWR top0.c_out_calc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_15133_ net520 _07162_ _07163_ VGND VGND VPWR VPWR _07232_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19941_ _11484_ _11504_ VGND VGND VPWR VPWR _11812_ sky130_fd_sc_hd__and2_1
X_15064_ net517 net493 VGND VGND VPWR VPWR _07163_ sky130_fd_sc_hd__nand2_2
XFILLER_0_120_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14015_ _06094_ _05822_ _06097_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__o21ai_1
X_19872_ _11519_ _11719_ _11732_ _11747_ VGND VGND VPWR VPWR _11748_ sky130_fd_sc_hd__o31ai_1
X_18823_ net373 net362 _10793_ net323 VGND VGND VPWR VPWR _10799_ sky130_fd_sc_hd__o22a_1
Xclkbuf_3_2__f_clk_mosi clknet_0_clk_mosi VGND VGND VPWR VPWR clknet_3_2__leaf_clk_mosi
+ sky130_fd_sc_hd__clkbuf_16
X_18754_ _10707_ _10730_ VGND VGND VPWR VPWR _10731_ sky130_fd_sc_hd__xnor2_4
X_15966_ _08039_ _08060_ VGND VGND VPWR VPWR _08061_ sky130_fd_sc_hd__xnor2_2
X_17705_ net385 net381 VGND VGND VPWR VPWR _09692_ sky130_fd_sc_hd__nand2_1
X_14917_ _07079_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__clkbuf_1
X_18685_ net401 _09433_ _10228_ VGND VGND VPWR VPWR _10663_ sky130_fd_sc_hd__or3_2
XFILLER_0_37_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15897_ top0.pid_q.out\[3\] VGND VGND VPWR VPWR _07993_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_159_Right_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17636_ _09621_ _09622_ VGND VGND VPWR VPWR _09623_ sky130_fd_sc_hd__xnor2_1
X_14848_ _07043_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17567_ _09551_ _09553_ VGND VGND VPWR VPWR _09554_ sky130_fd_sc_hd__nand2_1
X_14779_ _06974_ _06979_ VGND VGND VPWR VPWR _06980_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_187_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16518_ _08393_ _08410_ _08490_ VGND VGND VPWR VPWR _08606_ sky130_fd_sc_hd__a21o_1
X_19306_ _11119_ _11245_ _11246_ VGND VGND VPWR VPWR _11247_ sky130_fd_sc_hd__and3_1
XFILLER_0_184_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17498_ _09483_ _09484_ VGND VGND VPWR VPWR _09485_ sky130_fd_sc_hd__xor2_1
XFILLER_0_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16449_ _08533_ _08536_ VGND VGND VPWR VPWR _08538_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19237_ _11183_ _11175_ top0.pid_d.prev_error\[6\] VGND VGND VPWR VPWR _11184_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_183_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19168_ top0.pid_d.state\[0\] net433 _07136_ VGND VGND VPWR VPWR _11122_ sky130_fd_sc_hd__or3_1
XFILLER_0_147_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18119_ net307 VGND VGND VPWR VPWR _10103_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19099_ _10848_ _11069_ _11070_ VGND VGND VPWR VPWR _11071_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21130_ _12094_ _12917_ _12972_ net255 _12974_ VGND VGND VPWR VPWR _12975_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21061_ _12847_ _12900_ VGND VGND VPWR VPWR _12907_ sky130_fd_sc_hd__nand2_1
Xfanout404 top0.pid_d.mult0.a\[6\] VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout415 net417 VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__clkbuf_4
Xfanout426 net427 VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__clkbuf_4
X_20012_ _11876_ _11810_ _11877_ net195 _11512_ VGND VGND VPWR VPWR _11878_ sky130_fd_sc_hd__a221o_1
Xfanout437 net440 VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__buf_2
Xfanout448 top0.pid_q.mult0.b\[13\] VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkbuf_4
Xfanout459 net460 VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__buf_2
XFILLER_0_193_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24820_ _04078_ _04086_ _04171_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__a21oi_2
X_24751_ _04094_ _04103_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__xnor2_2
X_21963_ net160 net130 _01372_ net165 VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23702_ _03059_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20914_ net218 net232 VGND VGND VPWR VPWR _12762_ sky130_fd_sc_hd__or2b_1
XFILLER_0_179_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24682_ _03916_ _03917_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__nand2_1
X_21894_ _01411_ _01410_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__nor2_4
X_26421_ clknet_leaf_60_clk_sys _00062_ net650 VGND VGND VPWR VPWR top0.kpq\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23633_ _02990_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__clkbuf_4
X_20845_ net271 _12215_ _12691_ _12692_ _12693_ VGND VGND VPWR VPWR _12694_ sky130_fd_sc_hd__a41o_1
Xfanout11 net328 VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__buf_4
Xfanout22 net23 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout33 net35 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_4
X_26352_ spi0.data_packed\[74\] spi0.data_packed\[75\] net690 VGND VGND VPWR VPWR
+ _05408_ sky130_fd_sc_hd__mux2_1
Xfanout44 top0.periodTop_r\[8\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_4
X_23564_ net965 top0.matmul0.b\[5\] _02948_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__mux2_1
X_20776_ _11608_ _12611_ VGND VGND VPWR VPWR _12625_ sky130_fd_sc_hd__xnor2_1
Xfanout55 top0.periodTop_r\[4\] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
X_25303_ _04645_ _04648_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__xnor2_1
Xfanout66 net67 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout77 net78 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_4
X_22515_ _02053_ _02070_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__xnor2_1
X_26283_ _05373_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__clkbuf_1
Xfanout88 net89 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_4
Xfanout99 net101 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_4
X_23495_ _02912_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25234_ _04382_ _04580_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_190_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22446_ _01999_ _02002_ _01885_ VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_161_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25165_ _04510_ _04512_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22377_ _01832_ _01859_ _01935_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__a21oi_1
X_24116_ _02989_ _02991_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__nor2_4
X_21328_ net248 net227 VGND VGND VPWR VPWR _13170_ sky130_fd_sc_hd__xnor2_2
X_25096_ _04364_ _04366_ _04444_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24047_ _03250_ _03252_ _03363_ _03120_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__o211a_1
X_21259_ _13053_ _13098_ _13102_ VGND VGND VPWR VPWR _13103_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15820_ net488 net502 VGND VGND VPWR VPWR _07916_ sky130_fd_sc_hd__nand2_1
X_25998_ _05013_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15751_ _07753_ _07758_ VGND VGND VPWR VPWR _07848_ sky130_fd_sc_hd__nand2_1
X_24949_ _04287_ _04299_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__xor2_1
X_14702_ _06904_ _06905_ VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__nor2_2
X_18470_ net396 net312 VGND VGND VPWR VPWR _10450_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15682_ _07663_ _07667_ VGND VGND VPWR VPWR _07780_ sky130_fd_sc_hd__nand2_1
X_17421_ net419 net333 VGND VGND VPWR VPWR _09408_ sky130_fd_sc_hd__nand2_1
X_14633_ _06760_ _06762_ _06761_ VGND VGND VPWR VPWR _06838_ sky130_fd_sc_hd__o21a_1
X_26619_ clknet_leaf_28_clk_sys _00236_ net623 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17352_ _07141_ VGND VGND VPWR VPWR _09339_ sky130_fd_sc_hd__clkbuf_4
X_14564_ _06768_ _06769_ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16303_ _08392_ _08390_ VGND VGND VPWR VPWR _08394_ sky130_fd_sc_hd__and2b_1
X_13515_ net64 _05726_ _05727_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__and3_1
X_17283_ top0.matmul0.matmul_stage_inst.mult2\[5\] VGND VGND VPWR VPWR _09280_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14495_ net41 _05726_ _05727_ VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__and3_1
X_19022_ _10968_ _10969_ _10963_ VGND VGND VPWR VPWR _10995_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16234_ _08324_ _08245_ top0.pid_q.out\[7\] VGND VGND VPWR VPWR _08325_ sky130_fd_sc_hd__o21ba_1
X_13446_ _05536_ _05637_ _05638_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16165_ net523 net446 VGND VGND VPWR VPWR _08257_ sky130_fd_sc_hd__nand2_2
X_13377_ net61 _05551_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15116_ _07211_ _07212_ _07214_ VGND VGND VPWR VPWR _07215_ sky130_fd_sc_hd__nand3_1
X_16096_ _08185_ _08188_ VGND VGND VPWR VPWR _08189_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19924_ _11632_ net202 net184 VGND VGND VPWR VPWR _11796_ sky130_fd_sc_hd__or3_1
X_15047_ net517 net490 VGND VGND VPWR VPWR _07146_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19855_ _11731_ VGND VGND VPWR VPWR _11732_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_79_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18806_ net371 net366 _10780_ _10781_ _09364_ VGND VGND VPWR VPWR _10782_ sky130_fd_sc_hd__a32o_1
X_19786_ _11621_ _11665_ _11666_ _11667_ VGND VGND VPWR VPWR _11668_ sky130_fd_sc_hd__a31o_1
X_16998_ top0.pid_q.prev_error\[12\] top0.pid_q.curr_error\[12\] _09049_ VGND VGND
+ VPWR VPWR _09052_ sky130_fd_sc_hd__o21ba_1
X_18737_ _10710_ _10713_ VGND VGND VPWR VPWR _10714_ sky130_fd_sc_hd__xnor2_2
X_15949_ _08042_ _08043_ VGND VGND VPWR VPWR _08044_ sky130_fd_sc_hd__xor2_1
X_18668_ _10642_ _10645_ VGND VGND VPWR VPWR _10646_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17619_ net417 net331 VGND VGND VPWR VPWR _09606_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18599_ _10575_ _10577_ VGND VGND VPWR VPWR _10578_ sky130_fd_sc_hd__xor2_2
Xclkbuf_leaf_88_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_88_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20630_ net287 _12478_ VGND VGND VPWR VPWR _12479_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_88_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20561_ _12084_ _12116_ VGND VGND VPWR VPWR _12410_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22300_ _01832_ _01859_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__xor2_2
XFILLER_0_27_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20492_ _12330_ _12332_ _12340_ VGND VGND VPWR VPWR _12341_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23280_ net182 _02727_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22231_ _11674_ _01775_ _01776_ _01783_ _01791_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__o41a_1
XFILLER_0_48_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22162_ _01229_ _01242_ _01723_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21113_ _12878_ _12958_ VGND VGND VPWR VPWR _12959_ sky130_fd_sc_hd__nor2_1
X_26970_ clknet_leaf_29_clk_sys _00587_ net623 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_22093_ _01619_ _01628_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__and2_1
Xfanout201 net203 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout212 top0.cordic0.slte0.opA\[15\] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__buf_2
X_25921_ _05102_ _05126_ _05135_ _05130_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__a31o_1
X_21044_ _12863_ _12835_ VGND VGND VPWR VPWR _12890_ sky130_fd_sc_hd__or2b_1
Xfanout223 net224 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_4
Xfanout234 net235 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_201_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout245 top0.cordic0.vec\[0\]\[11\] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__buf_4
Xfanout256 net257 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__clkbuf_4
Xfanout267 net268 VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_4
X_25852_ top0.matmul0.beta_pass\[6\] _05065_ _05072_ top0.matmul0.alpha_pass\[6\]
+ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__a22oi_2
Xfanout278 net279 VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__buf_4
XFILLER_0_119_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout289 net293 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__clkbuf_4
X_24803_ _04155_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25783_ net208 net205 VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__or2b_2
XFILLER_0_202_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22995_ net169 _02483_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24734_ _04081_ _04086_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__xnor2_2
X_21946_ net165 net137 _01356_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24665_ _03252_ _03826_ _03875_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21877_ _01412_ _01438_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26404_ clknet_leaf_98_clk_sys _00045_ net589 VGND VGND VPWR VPWR top0.kpd\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23616_ top0.matmul0.alpha_pass\[15\] _09337_ net561 VGND VGND VPWR VPWR _02975_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20828_ _12230_ _12240_ _12676_ VGND VGND VPWR VPWR _12677_ sky130_fd_sc_hd__o21a_1
X_24596_ _03833_ _03837_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26335_ _05399_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__clkbuf_1
X_23547_ top0.a_in_matmul\[13\] top0.matmul0.a\[13\] _02937_ VGND VGND VPWR VPWR _02940_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20759_ _11408_ _12264_ _12326_ _12607_ VGND VGND VPWR VPWR _12608_ sky130_fd_sc_hd__o31a_2
XFILLER_0_52_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13300_ net42 _05489_ _05491_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14280_ net48 _05726_ _05727_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__and3_1
X_26266_ spi0.data_packed\[31\] spi0.data_packed\[32\] net690 VGND VGND VPWR VPWR
+ _05365_ sky130_fd_sc_hd__mux2_1
X_23478_ _02903_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25217_ _04558_ _04563_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__xor2_1
X_13231_ _05451_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__clkbuf_1
X_22429_ _01985_ _01986_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__or2b_1
X_26197_ _05329_ top0.cordic0.slte0.opB\[15\] _12003_ VGND VGND VPWR VPWR _05330_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25148_ _04494_ _04495_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25079_ net1017 _04097_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__nor2_2
X_17970_ _09948_ _09955_ VGND VGND VPWR VPWR _09956_ sky130_fd_sc_hd__xnor2_1
X_16921_ net550 _08979_ _08980_ VGND VGND VPWR VPWR _08981_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19640_ _11443_ _11445_ _11449_ _11450_ _11451_ VGND VGND VPWR VPWR _11528_ sky130_fd_sc_hd__a32o_1
X_16852_ top0.currT_r\[2\] _08903_ VGND VGND VPWR VPWR _08916_ sky130_fd_sc_hd__or2_1
X_15803_ top0.pid_q.out\[2\] top0.pid_q.curr_int\[2\] _07802_ _07803_ VGND VGND VPWR
+ VPWR _07899_ sky130_fd_sc_hd__a22oi_2
X_19571_ top0.cordic0.slte0.opB\[5\] top0.cordic0.slte0.opA\[5\] VGND VGND VPWR VPWR
+ _11460_ sky130_fd_sc_hd__nand2_1
X_16783_ net539 _08856_ _08859_ net757 _08864_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__a221o_1
XFILLER_0_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13995_ _06206_ _06207_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__xor2_2
X_18522_ _10493_ _10501_ VGND VGND VPWR VPWR _10502_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15734_ _07828_ _07830_ VGND VGND VPWR VPWR _07831_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18453_ _10331_ _10343_ _10420_ VGND VGND VPWR VPWR _10433_ sky130_fd_sc_hd__or3_2
X_15665_ _07738_ _07762_ VGND VGND VPWR VPWR _07763_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14616_ _06775_ _06782_ VGND VGND VPWR VPWR _06821_ sky130_fd_sc_hd__and2b_1
X_17404_ _09386_ _09390_ VGND VGND VPWR VPWR _09391_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18384_ net338 net369 VGND VGND VPWR VPWR _10365_ sky130_fd_sc_hd__nand2_2
XFILLER_0_157_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15596_ _07690_ _07692_ _07693_ _07688_ VGND VGND VPWR VPWR _07695_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_29_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17335_ _09323_ _09324_ VGND VGND VPWR VPWR _09325_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_157_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14547_ _06649_ _06725_ _06752_ VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__o21a_2
XFILLER_0_44_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17266_ top0.matmul0.matmul_stage_inst.mult1\[3\] top0.matmul0.matmul_stage_inst.mult2\[3\]
+ VGND VGND VPWR VPWR _09266_ sky130_fd_sc_hd__xnor2_1
X_14478_ _06672_ _06673_ _06683_ _06684_ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16217_ _08307_ _08308_ VGND VGND VPWR VPWR _08309_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19005_ _10976_ _10978_ VGND VGND VPWR VPWR _10979_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13429_ _05605_ _05640_ _05641_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17197_ top0.pid_q.curr_int\[9\] _09141_ _09206_ _09136_ VGND VGND VPWR VPWR _00222_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16148_ top0.pid_q.out\[6\] _08237_ _08240_ VGND VGND VPWR VPWR _08241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16079_ _08168_ _08171_ VGND VGND VPWR VPWR _08172_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19907_ _11779_ _11780_ VGND VGND VPWR VPWR _11781_ sky130_fd_sc_hd__nor2_1
X_19838_ _11632_ net83 _11575_ _11715_ VGND VGND VPWR VPWR _11716_ sky130_fd_sc_hd__o22a_1
XFILLER_0_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 cs VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
X_19769_ _11650_ _11646_ net1020 VGND VGND VPWR VPWR _11652_ sky130_fd_sc_hd__a21oi_1
X_21800_ _01355_ _01361_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_79_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22780_ top0.svm0.counter\[13\] top0.svm0.counter\[14\] top0.svm0.counter\[15\] _02303_
+ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__or4_1
XFILLER_0_79_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21731_ _01291_ _01292_ net139 VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_78_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24450_ net566 net558 top0.matmul0.matmul_stage_inst.e\[15\] VGND VGND VPWR VPWR
+ _03806_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21662_ net111 net107 VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_164_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23401_ net111 _02827_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20613_ _12440_ _12454_ VGND VGND VPWR VPWR _12462_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24381_ _03192_ _03174_ _03737_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__a21o_2
XFILLER_0_47_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21593_ net141 net148 VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26120_ spi0.data_packed\[17\] _05279_ _05280_ net919 VGND VGND VPWR VPWR _00798_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23332_ _02774_ _02776_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20544_ _12360_ _12387_ _12372_ VGND VGND VPWR VPWR _12393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26051_ _05240_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23263_ net215 _11633_ _02711_ _11409_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20475_ _12283_ _12323_ VGND VGND VPWR VPWR _12324_ sky130_fd_sc_hd__xnor2_4
X_25002_ _04348_ _04351_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22214_ net98 net94 VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_132_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23194_ _05719_ _07000_ _02648_ net809 VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22145_ _01105_ net127 VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__nand2_1
X_26953_ clknet_leaf_16_clk_sys _00570_ net613 VGND VGND VPWR VPWR top0.matmul0.b\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_22076_ _01610_ _01612_ _01637_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_199_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25904_ net429 _05104_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__nor2_1
X_21027_ _12868_ _12873_ VGND VGND VPWR VPWR _12874_ sky130_fd_sc_hd__xnor2_2
X_26884_ clknet_leaf_38_clk_sys _00501_ net677 VGND VGND VPWR VPWR top0.svm0.tB\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25835_ _05052_ _05054_ _05057_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_96_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13780_ _05991_ _05989_ _05987_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__o21ai_1
X_25766_ top0.matmul0.matmul_stage_inst.a\[11\] _04900_ _05457_ VGND VGND VPWR VPWR
+ _05004_ sky130_fd_sc_hd__mux2_1
X_22978_ _02485_ _02480_ _02486_ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__a21o_1
X_24717_ _03502_ _03687_ _03985_ _03986_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__a22o_1
X_21929_ _01489_ _01490_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__or2_1
X_25697_ _04962_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__clkbuf_1
X_15450_ _07273_ _07271_ _07548_ VGND VGND VPWR VPWR _07549_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24648_ _03883_ _03884_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14401_ _06608_ _06609_ VGND VGND VPWR VPWR _06610_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15381_ net538 net486 VGND VGND VPWR VPWR _07480_ sky130_fd_sc_hd__nand2_1
X_24579_ _03774_ _03932_ _03933_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17120_ net553 _09137_ _09138_ _08887_ VGND VGND VPWR VPWR _09139_ sky130_fd_sc_hd__a211o_1
XFILLER_0_182_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14332_ _06532_ _06541_ VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26318_ spi0.data_packed\[57\] spi0.data_packed\[58\] net699 VGND VGND VPWR VPWR
+ _05391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27298_ clknet_3_1__leaf_clk_mosi _00912_ VGND VGND VPWR VPWR spi0.opcode\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17051_ net551 _00008_ _08854_ VGND VGND VPWR VPWR _09101_ sky130_fd_sc_hd__and3b_1
XFILLER_0_80_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14263_ net853 _06280_ _06473_ _06381_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26249_ _05356_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__clkbuf_1
X_16002_ _08094_ _08095_ VGND VGND VPWR VPWR _08096_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13214_ net997 _05432_ _05439_ VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__a21o_1
X_14194_ _06403_ _06404_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_36_clk_sys clknet_3_7__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_36_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17953_ _09935_ _09938_ VGND VGND VPWR VPWR _09939_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16904_ _08963_ _08964_ VGND VGND VPWR VPWR _08965_ sky130_fd_sc_hd__and2_1
X_17884_ net424 net315 VGND VGND VPWR VPWR _09871_ sky130_fd_sc_hd__nand2_1
X_19623_ _11511_ VGND VGND VPWR VPWR _11512_ sky130_fd_sc_hd__buf_6
X_16835_ _08899_ VGND VGND VPWR VPWR _08900_ sky130_fd_sc_hd__buf_4
XFILLER_0_189_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19554_ _11420_ net179 _11442_ VGND VGND VPWR VPWR _11443_ sky130_fd_sc_hd__or3_2
X_13978_ _06190_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__clkbuf_2
X_16766_ top0.pid_q.out\[15\] _05442_ _07704_ VGND VGND VPWR VPWR _08850_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18505_ _10483_ _10484_ VGND VGND VPWR VPWR _10485_ sky130_fd_sc_hd__xnor2_2
X_15717_ net469 net515 VGND VGND VPWR VPWR _07814_ sky130_fd_sc_hd__nand2_1
XFILLER_0_198_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16697_ _08749_ _08781_ VGND VGND VPWR VPWR _08782_ sky130_fd_sc_hd__xnor2_2
X_19485_ _11368_ _11377_ _11378_ VGND VGND VPWR VPWR _11379_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18436_ _10415_ _10416_ VGND VGND VPWR VPWR _10417_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15648_ _07638_ _07639_ _07640_ VGND VGND VPWR VPWR _07746_ sky130_fd_sc_hd__o21a_1
XFILLER_0_173_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18367_ _10260_ _10265_ _10347_ _10255_ VGND VGND VPWR VPWR _10348_ sky130_fd_sc_hd__a2bb2o_1
X_15579_ _07296_ VGND VGND VPWR VPWR _07678_ sky130_fd_sc_hd__inv_2
X_17318_ top0.matmul0.matmul_stage_inst.mult2\[10\] VGND VGND VPWR VPWR _09310_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18298_ net325 net386 VGND VGND VPWR VPWR _10280_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17249_ top0.matmul0.beta_pass\[0\] _09251_ net563 VGND VGND VPWR VPWR _09252_ sky130_fd_sc_hd__mux2_1
X_20260_ net305 net290 VGND VGND VPWR VPWR _12109_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20191_ net252 _12039_ VGND VGND VPWR VPWR _12040_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_12_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23950_ _03302_ _03303_ _03307_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__o21a_2
X_22901_ top0.svm0.tC\[7\] _02418_ top0.svm0.counter\[7\] VGND VGND VPWR VPWR _02419_
+ sky130_fd_sc_hd__o21ba_1
X_23881_ _03024_ _03025_ _03027_ _03028_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__o22a_1
X_25620_ top0.matmul0.op\[1\] top0.matmul0.cos\[13\] VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22832_ top0.svm0.counter\[1\] VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25551_ _04862_ VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22763_ net976 _02292_ _02295_ top0.pid_q.curr_int\[7\] VGND VGND VPWR VPWR _00426_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24502_ _03654_ _03657_ _03847_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21714_ _01265_ _01275_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__nor2_1
X_25482_ _04821_ _04756_ _04764_ _04824_ _04661_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__a32o_1
XFILLER_0_17_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22694_ net90 _01849_ _01948_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27221_ clknet_3_5__leaf_clk_mosi _00835_ VGND VGND VPWR VPWR spi0.data_packed\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_24433_ _03786_ _03787_ _03784_ _03785_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__a211oi_2
X_21645_ _01139_ _01206_ net155 VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__mux2_2
XFILLER_0_81_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27152_ clknet_leaf_11_clk_sys _00766_ net601 VGND VGND VPWR VPWR top0.a_in_matmul\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_24364_ _03195_ _03719_ _03720_ _03324_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__o211a_1
X_21576_ net131 net126 VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__nor2_1
X_26103_ top0.periodTop\[2\] _05276_ _05278_ net59 VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23315_ net140 _02744_ _02758_ _02760_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__a22o_1
X_27083_ clknet_leaf_20_clk_sys _00700_ net609 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_20527_ _12372_ _12375_ VGND VGND VPWR VPWR _12376_ sky130_fd_sc_hd__xnor2_1
X_24295_ _03646_ _03651_ _03450_ _03618_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__a211o_2
XFILLER_0_127_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26034_ top0.a_in_matmul\[1\] _05226_ _05196_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__mux2_1
X_23246_ _02686_ _02695_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__xnor2_1
X_20458_ net287 _12302_ VGND VGND VPWR VPWR _12307_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23177_ _05717_ _07038_ _02644_ net800 VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20389_ net235 net226 VGND VGND VPWR VPWR _12238_ sky130_fd_sc_hd__nand2_2
X_22128_ net96 _01225_ _11674_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__a21oi_1
X_14950_ _07096_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__clkbuf_1
X_22059_ _01549_ _01553_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__or2_1
X_26936_ clknet_leaf_8_clk_sys _00553_ net595 VGND VGND VPWR VPWR top0.matmul0.a\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13901_ net37 _05475_ _05476_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__and3_1
X_14881_ _07060_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__clkbuf_1
X_26867_ clknet_leaf_39_clk_sys _00484_ net683 VGND VGND VPWR VPWR top0.svm0.tA\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_16620_ _08700_ _08705_ VGND VGND VPWR VPWR _08706_ sky130_fd_sc_hd__xor2_1
X_13832_ net59 _05497_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_199_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25818_ _05042_ _05039_ _05035_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__o21bai_2
X_26798_ clknet_leaf_102_clk_sys _00415_ net589 VGND VGND VPWR VPWR top0.cordic0.gm0.iter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16551_ net450 net503 VGND VGND VPWR VPWR _08638_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13763_ _05974_ _05975_ net58 _05495_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__o211a_1
X_25749_ _04995_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15502_ _07599_ VGND VGND VPWR VPWR _07601_ sky130_fd_sc_hd__inv_2
X_16482_ _08497_ _08498_ _08496_ VGND VGND VPWR VPWR _08570_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19270_ top0.pid_d.curr_error\[9\] VGND VGND VPWR VPWR _11214_ sky130_fd_sc_hd__inv_2
X_13694_ _05875_ _05878_ _05906_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18221_ net405 _10203_ _09363_ VGND VGND VPWR VPWR _10204_ sky130_fd_sc_hd__o21ai_1
X_15433_ _07527_ _07528_ _07531_ VGND VGND VPWR VPWR _07532_ sky130_fd_sc_hd__a21o_1
XFILLER_0_183_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18152_ _10044_ _10045_ _10046_ VGND VGND VPWR VPWR _10136_ sky130_fd_sc_hd__a21o_1
X_15364_ _07443_ _07462_ VGND VGND VPWR VPWR _07463_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14315_ _06421_ _06423_ _06524_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__a21oi_2
X_17103_ top0.pid_q.curr_error\[10\] _08860_ _09116_ VGND VGND VPWR VPWR _09128_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18083_ top0.pid_d.out\[2\] _09339_ _10066_ _10067_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15295_ _07354_ _07364_ VGND VGND VPWR VPWR _07394_ sky130_fd_sc_hd__xor2_1
XFILLER_0_180_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17034_ _09081_ top0.currT_r\[14\] _08900_ _09085_ VGND VGND VPWR VPWR _09086_ sky130_fd_sc_hd__o31a_1
X_14246_ _06455_ _06456_ VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__xor2_1
Xhold309 top0.b_in_matmul\[14\] VGND VGND VPWR VPWR net1009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14177_ _06239_ _06251_ _06252_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_180_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18985_ _10845_ _10958_ VGND VGND VPWR VPWR _10959_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17936_ _09920_ _09921_ VGND VGND VPWR VPWR _09922_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17867_ _09778_ _09852_ _09853_ VGND VGND VPWR VPWR _09854_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_84_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19606_ _11494_ _11492_ VGND VGND VPWR VPWR _11495_ sky130_fd_sc_hd__or2_1
XFILLER_0_178_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16818_ net547 _08884_ VGND VGND VPWR VPWR _08885_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17798_ _09783_ _09784_ VGND VGND VPWR VPWR _09785_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19537_ net194 net203 VGND VGND VPWR VPWR _11427_ sky130_fd_sc_hd__or2_2
X_16749_ _08721_ _08753_ _08832_ VGND VGND VPWR VPWR _08833_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_202_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19468_ _11289_ VGND VGND VPWR VPWR _11364_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18419_ _10270_ _10302_ _10301_ VGND VGND VPWR VPWR _10400_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_173_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19399_ _11301_ _11302_ VGND VGND VPWR VPWR _11303_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21430_ _00966_ _00995_ _00987_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21361_ _13161_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__inv_2
XFILLER_0_185_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23100_ top0.svm0.delta\[1\] net555 _02440_ _02596_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_47_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20312_ _12154_ _12159_ _12160_ VGND VGND VPWR VPWR _12161_ sky130_fd_sc_hd__o21a_4
X_24080_ _03437_ _03332_ _03329_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_31_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21292_ _13036_ _13134_ VGND VGND VPWR VPWR _13135_ sky130_fd_sc_hd__xor2_2
XFILLER_0_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23031_ _07115_ top0.svm0.counter\[15\] VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__nor2_1
X_20243_ _12086_ _12088_ _12091_ VGND VGND VPWR VPWR _12092_ sky130_fd_sc_hd__nand3_1
XFILLER_0_40_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20174_ _12010_ _12011_ _12014_ _05439_ _12025_ VGND VGND VPWR VPWR _12026_ sky130_fd_sc_hd__o221a_2
XFILLER_0_196_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24982_ _04315_ _04317_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__or2_1
X_23933_ _03276_ _03284_ _03285_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__o21a_1
X_26721_ clknet_leaf_81_clk_sys _00338_ net636 VGND VGND VPWR VPWR top0.pid_d.curr_int\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_192_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26652_ clknet_leaf_75_clk_sys _00269_ net639 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_23864_ _03220_ _03221_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25603_ _04886_ top0.matmul0.cos\[5\] _04878_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__or3_1
X_22815_ top0.svm0.counter\[8\] top0.svm0.tA\[8\] VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__or2_1
XFILLER_0_169_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26583_ clknet_leaf_53_clk_sys _00206_ net674 VGND VGND VPWR VPWR top0.pid_q.prev_error\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23795_ _03149_ _03152_ VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25534_ _04853_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__clkbuf_1
X_22746_ net186 _02288_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25465_ _04748_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22677_ _02207_ _02228_ _02180_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__or3b_1
XFILLER_0_165_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27204_ clknet_leaf_92_clk_sys _00818_ net599 VGND VGND VPWR VPWR top0.cordic0.slte0.opB\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_24416_ _03768_ _03771_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21628_ _01188_ _01189_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_106_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25396_ _04685_ _04688_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_33_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27135_ clknet_leaf_12_clk_sys _00749_ net616 VGND VGND VPWR VPWR top0.b_in_matmul\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_24347_ _03202_ _03203_ _03060_ _03124_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21559_ _01117_ _01120_ VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14100_ _06222_ _06224_ _06223_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27066_ clknet_leaf_8_clk_sys _00683_ net592 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.c\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_15080_ net540 net460 VGND VGND VPWR VPWR _07179_ sky130_fd_sc_hd__nand2_1
X_24278_ _03627_ _03635_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14031_ _06148_ _06149_ _06243_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__o21a_1
X_26017_ top0.matmul0.beta_pass\[13\] _05203_ _05213_ VGND VGND VPWR VPWR _05214_
+ sky130_fd_sc_hd__a21o_1
X_23229_ _11425_ _02667_ _02668_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_129_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_1__f_clk_mosi clknet_0_clk_mosi VGND VGND VPWR VPWR clknet_3_1__leaf_clk_mosi
+ sky130_fd_sc_hd__clkbuf_16
X_18770_ _10744_ _10746_ VGND VGND VPWR VPWR _10747_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_42_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15982_ _08076_ _07899_ _07900_ _07993_ VGND VGND VPWR VPWR _08077_ sky130_fd_sc_hd__o31a_1
X_17721_ net385 net352 VGND VGND VPWR VPWR _09708_ sky130_fd_sc_hd__nand2_1
X_14933_ spi0.data_packed\[41\] top0.kid\[9\] _07086_ VGND VGND VPWR VPWR _07088_
+ sky130_fd_sc_hd__mux2_1
X_26919_ clknet_leaf_1_clk_sys _00536_ net582 VGND VGND VPWR VPWR top0.matmul0.sin\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17652_ net388 net359 _09637_ VGND VGND VPWR VPWR _09639_ sky130_fd_sc_hd__mux2_1
X_14864_ _07051_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16603_ _08601_ _08676_ VGND VGND VPWR VPWR _08689_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13815_ _05996_ _05997_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__xor2_2
X_14795_ _06992_ _06994_ _06995_ _06910_ _06991_ VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__o221a_1
X_17583_ net412 net418 _09395_ VGND VGND VPWR VPWR _09570_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19322_ top0.matmul0.alpha_pass\[14\] _11245_ VGND VGND VPWR VPWR _11262_ sky130_fd_sc_hd__nor2_1
X_13746_ _05924_ _05958_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__xnor2_1
X_16534_ top0.pid_q.curr_int\[12\] VGND VGND VPWR VPWR _08621_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19253_ _11196_ _11197_ VGND VGND VPWR VPWR _11199_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13677_ net58 _05517_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__nand2_1
X_16465_ _08553_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_51_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18204_ top0.pid_d.mult0.b\[4\] net372 VGND VGND VPWR VPWR _10187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15416_ _07432_ _07453_ VGND VGND VPWR VPWR _07515_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19184_ top0.pid_d.prev_error\[2\] top0.pid_d.curr_error\[2\] VGND VGND VPWR VPWR
+ _11136_ sky130_fd_sc_hd__xor2_1
X_16396_ top0.pid_q.out\[9\] top0.pid_q.curr_int\[9\] VGND VGND VPWR VPWR _08485_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18135_ _10115_ _10118_ VGND VGND VPWR VPWR _10119_ sky130_fd_sc_hd__xnor2_2
X_15347_ _07444_ _07445_ net534 VGND VGND VPWR VPWR _07446_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_0_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold106 top0.svm0.tA\[11\] VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__dlygate4sd3_1
X_18066_ _10040_ _10049_ VGND VGND VPWR VPWR _10051_ sky130_fd_sc_hd__or2_1
X_15278_ _07376_ VGND VGND VPWR VPWR _07377_ sky130_fd_sc_hd__inv_2
Xhold117 top0.svm0.tC\[9\] VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold128 top0.pid_d.curr_int\[10\] VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 top0.svm0.tB\[15\] VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ _06435_ _06439_ VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__xnor2_4
X_17017_ top0.currT_r\[14\] _09069_ VGND VGND VPWR VPWR _09070_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout608 net630 VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout619 net620 VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_60_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18968_ _10940_ _10941_ VGND VGND VPWR VPWR _10942_ sky130_fd_sc_hd__or2b_1
XFILLER_0_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17919_ net332 net399 VGND VGND VPWR VPWR _09905_ sky130_fd_sc_hd__nand2_1
X_18899_ _10772_ _10873_ VGND VGND VPWR VPWR _10874_ sky130_fd_sc_hd__xnor2_2
X_20930_ net276 net256 VGND VGND VPWR VPWR _12778_ sky130_fd_sc_hd__xor2_2
XFILLER_0_152_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20861_ _12704_ _12706_ _12708_ VGND VGND VPWR VPWR _12710_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22600_ net101 net97 net87 _11674_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__a31o_1
X_23580_ top0.b_in_matmul\[13\] top0.matmul0.b\[13\] _02948_ VGND VGND VPWR VPWR _02957_
+ sky130_fd_sc_hd__mux2_1
X_20792_ _12587_ _12640_ VGND VGND VPWR VPWR _12641_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22531_ _02003_ _02084_ _02085_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__o21a_1
XFILLER_0_187_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25250_ _04525_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22462_ _01224_ _02018_ net125 VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24201_ _03540_ _03546_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__xor2_2
X_21413_ _00977_ _00978_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__nand2_1
X_25181_ _04306_ _04455_ _04527_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__or3_1
XFILLER_0_162_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22393_ _01936_ _01949_ _01950_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24132_ _03473_ _03475_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__xnor2_2
X_21344_ _13184_ _13185_ VGND VGND VPWR VPWR _13186_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24063_ _03400_ _03407_ _03408_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21275_ _13114_ _13117_ VGND VGND VPWR VPWR _13118_ sky130_fd_sc_hd__or2_1
X_23014_ top0.svm0.counter\[13\] _02439_ _02517_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__or3_1
X_20226_ net252 net240 VGND VGND VPWR VPWR _12075_ sky130_fd_sc_hd__nand2_2
XFILLER_0_21_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20157_ net207 VGND VGND VPWR VPWR _12009_ sky130_fd_sc_hd__inv_2
X_24965_ _04172_ _04178_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__or2_1
X_20088_ _11714_ _11629_ _11936_ _11428_ VGND VGND VPWR VPWR _11948_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26704_ clknet_leaf_84_clk_sys _00321_ net646 VGND VGND VPWR VPWR top0.pid_d.prev_error\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_23916_ _03237_ _03242_ _03246_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24896_ _04166_ _04241_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23847_ _03201_ _03204_ VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__xnor2_2
X_26635_ clknet_leaf_75_clk_sys _00252_ net637 VGND VGND VPWR VPWR top0.pid_d.out\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_170_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13600_ _05811_ _05812_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14580_ _06714_ _06725_ VGND VGND VPWR VPWR _06786_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26566_ clknet_leaf_53_clk_sys _00189_ net672 VGND VGND VPWR VPWR top0.pid_q.curr_error\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_23778_ _03110_ _03135_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__nor2_1
XFILLER_0_178_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13531_ _05700_ _05703_ _05706_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__a21oi_1
X_25517_ _04844_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22729_ _02277_ _02278_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26497_ clknet_leaf_72_clk_sys _00120_ net655 VGND VGND VPWR VPWR top0.pid_d.prev_int\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_137_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16250_ net476 _08141_ net473 VGND VGND VPWR VPWR _08341_ sky130_fd_sc_hd__o21a_1
X_13462_ _05655_ _05674_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__xnor2_1
X_25448_ _04789_ _04790_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__or2b_1
XFILLER_0_152_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15201_ _07263_ _07299_ VGND VGND VPWR VPWR _07300_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16181_ net463 net507 VGND VGND VPWR VPWR _08273_ sky130_fd_sc_hd__nand2_1
X_13393_ net61 _05605_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__nand2_2
X_25379_ _04272_ _04131_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__nor2_2
XFILLER_0_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15132_ net522 _07227_ _07229_ _07230_ VGND VGND VPWR VPWR _07231_ sky130_fd_sc_hd__a31o_1
X_27118_ clknet_leaf_33_clk_sys _00732_ net665 VGND VGND VPWR VPWR top0.c_out_calc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27049_ clknet_leaf_22_clk_sys _00666_ net607 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.d\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_19940_ net183 _11509_ VGND VGND VPWR VPWR _11811_ sky130_fd_sc_hd__or2_1
X_15063_ net522 net484 VGND VGND VPWR VPWR _07162_ sky130_fd_sc_hd__nand2_2
X_14014_ _06094_ _05822_ _06097_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__nor3_1
XFILLER_0_31_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19871_ _11719_ _11732_ net237 VGND VGND VPWR VPWR _11747_ sky130_fd_sc_hd__a21o_1
X_18822_ net320 net368 VGND VGND VPWR VPWR _10798_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18753_ _10728_ _10729_ VGND VGND VPWR VPWR _10730_ sky130_fd_sc_hd__nor2_2
X_15965_ _08040_ _08059_ VGND VGND VPWR VPWR _08060_ sky130_fd_sc_hd__xor2_1
X_17704_ net386 net381 VGND VGND VPWR VPWR _09691_ sky130_fd_sc_hd__or2_1
X_14916_ spi0.data_packed\[33\] top0.kid\[1\] _07075_ VGND VGND VPWR VPWR _07079_
+ sky130_fd_sc_hd__mux2_1
X_18684_ net396 _10660_ _10661_ VGND VGND VPWR VPWR _10662_ sky130_fd_sc_hd__o21ai_2
X_15896_ net545 _07903_ _07904_ net548 _07991_ VGND VGND VPWR VPWR _07992_ sky130_fd_sc_hd__a32o_1
XFILLER_0_187_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17635_ net398 net345 VGND VGND VPWR VPWR _09622_ sky130_fd_sc_hd__nand2_1
X_14847_ spi0.data_packed\[64\] top0.kpd\[0\] _07042_ VGND VGND VPWR VPWR _07043_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17566_ net412 _09531_ _09552_ VGND VGND VPWR VPWR _09553_ sky130_fd_sc_hd__or3_1
X_14778_ _06977_ _06978_ VGND VGND VPWR VPWR _06979_ sky130_fd_sc_hd__xor2_1
X_19305_ top0.matmul0.alpha_pass\[13\] _11241_ VGND VGND VPWR VPWR _11246_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16517_ _08546_ _08604_ VGND VGND VPWR VPWR _08605_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13729_ _05931_ _05935_ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17497_ net419 net330 VGND VGND VPWR VPWR _09484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19236_ top0.pid_d.curr_error\[6\] VGND VGND VPWR VPWR _11183_ sky130_fd_sc_hd__inv_2
X_16448_ _08533_ _08536_ VGND VGND VPWR VPWR _08537_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19167_ _11120_ VGND VGND VPWR VPWR _11121_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_182_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16379_ _08383_ _08381_ VGND VGND VPWR VPWR _08469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18118_ _10098_ _10101_ VGND VGND VPWR VPWR _10102_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19098_ _10772_ _11003_ _11010_ VGND VGND VPWR VPWR _11070_ sky130_fd_sc_hd__or3_1
XFILLER_0_83_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18049_ _10031_ _10033_ VGND VGND VPWR VPWR _10034_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_197_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_84_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_84_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21060_ _12902_ _12905_ _11673_ VGND VGND VPWR VPWR _12906_ sky130_fd_sc_hd__a21o_1
Xfanout405 top0.pid_d.mult0.a\[5\] VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkbuf_4
Xfanout416 net417 VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__buf_2
Xfanout427 top0.pid_d.mult0.a\[0\] VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__clkbuf_4
X_20011_ _11410_ top0.cordic0.gm0.iter\[2\] net183 VGND VGND VPWR VPWR _11877_ sky130_fd_sc_hd__a21oi_1
Xfanout438 net440 VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout449 net451 VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__buf_4
XFILLER_0_20_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24750_ _04096_ _04102_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21962_ net155 _01105_ net160 VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23701_ _03057_ _03058_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__or2_1
X_20913_ net229 net226 VGND VGND VPWR VPWR _12761_ sky130_fd_sc_hd__nor2b_4
X_24681_ _03899_ _04033_ _04034_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_178_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21893_ net148 _01392_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__xor2_4
XFILLER_0_49_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23632_ net570 top0.matmul0.matmul_stage_inst.b\[7\] top0.matmul0.matmul_stage_inst.a\[7\]
+ net566 VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__a22o_1
X_26420_ clknet_leaf_58_clk_sys _00061_ net650 VGND VGND VPWR VPWR top0.kpq\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_194_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20844_ net271 _12040_ _12215_ VGND VGND VPWR VPWR _12693_ sky130_fd_sc_hd__nor3_1
XFILLER_0_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout12 net321 VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__buf_4
X_26351_ _05407_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__clkbuf_1
Xfanout23 net24 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
X_23563_ _05460_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout34 net35 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
X_20775_ net303 _12623_ VGND VGND VPWR VPWR _12624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_175_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout45 top0.periodTop_r\[7\] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25302_ _04522_ _04647_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__xnor2_1
Xfanout56 net58 VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout67 net68 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_2
X_22514_ _02026_ _02069_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__xnor2_1
X_26282_ net967 net946 net688 VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout78 net81 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_4
X_23494_ top0.cordic0.cos\[2\] top0.matmul0.cos\[2\] _02904_ VGND VGND VPWR VPWR _02912_
+ sky130_fd_sc_hd__mux2_1
Xfanout89 top0.cordic0.vec\[1\]\[16\] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_4
X_25233_ _04516_ _04512_ _04571_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_190_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22445_ _01998_ _02001_ _01895_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25164_ _04443_ _04445_ _04511_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_107_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22376_ _01832_ _01859_ _01818_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24115_ _03458_ _03457_ _03472_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21327_ net257 _13165_ _13168_ VGND VGND VPWR VPWR _13169_ sky130_fd_sc_hd__a21oi_2
X_25095_ _04364_ _04366_ _04365_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_202_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24046_ _03195_ _03254_ _03324_ _03056_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__o211a_1
X_21258_ _13099_ _13100_ _13101_ VGND VGND VPWR VPWR _13102_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20209_ net299 _12056_ VGND VGND VPWR VPWR _12058_ sky130_fd_sc_hd__xnor2_1
X_21189_ _13028_ _13032_ VGND VGND VPWR VPWR _13033_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25997_ _12031_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15750_ _07837_ _07846_ VGND VGND VPWR VPWR _07847_ sky130_fd_sc_hd__xnor2_1
X_24948_ _04293_ _04298_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__xnor2_2
X_14701_ _06865_ _06903_ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__nor2_1
X_15681_ _07665_ VGND VGND VPWR VPWR _07779_ sky130_fd_sc_hd__inv_2
X_24879_ _04111_ _04229_ _04230_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__a21o_2
XFILLER_0_200_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17420_ net417 net337 VGND VGND VPWR VPWR _09407_ sky130_fd_sc_hd__and2_2
X_14632_ _06833_ _06836_ VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__xnor2_2
X_26618_ clknet_leaf_29_clk_sys _00235_ net623 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_142_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14563_ net39 _05726_ _05727_ VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__and3_1
X_17351_ _09338_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26549_ clknet_leaf_50_clk_sys _00172_ net675 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16302_ _08390_ _08392_ VGND VGND VPWR VPWR _08393_ sky130_fd_sc_hd__or2b_1
X_13514_ _05664_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14494_ net39 _05723_ _05724_ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__and3_1
XFILLER_0_165_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17282_ _09279_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19021_ _10935_ _10972_ _10973_ VGND VGND VPWR VPWR _10994_ sky130_fd_sc_hd__a21oi_2
X_13445_ _05657_ _05608_ _05609_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__or3_1
XFILLER_0_64_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16233_ top0.pid_q.curr_int\[7\] VGND VGND VPWR VPWR _08324_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13376_ net54 _05586_ _05588_ net57 VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16164_ net447 net521 VGND VGND VPWR VPWR _08256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15115_ net540 net538 _07181_ _07213_ VGND VGND VPWR VPWR _07214_ sky130_fd_sc_hd__nand4_2
X_16095_ _08186_ _08187_ VGND VGND VPWR VPWR _08188_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_192_Right_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19923_ _11789_ _11794_ _11795_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__o21ai_1
X_15046_ net520 net485 VGND VGND VPWR VPWR _07145_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19854_ net82 _11440_ _11730_ VGND VGND VPWR VPWR _11731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18805_ _10690_ net371 VGND VGND VPWR VPWR _10781_ sky130_fd_sc_hd__nor2_1
X_19785_ net266 _11643_ VGND VGND VPWR VPWR _11667_ sky130_fd_sc_hd__and2_1
X_16997_ net449 _08861_ _09045_ _09051_ _08889_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__o221a_1
X_18736_ _10711_ _10712_ VGND VGND VPWR VPWR _10713_ sky130_fd_sc_hd__xnor2_1
X_15948_ net474 net506 VGND VGND VPWR VPWR _08043_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18667_ _10484_ _10644_ VGND VGND VPWR VPWR _10645_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15879_ _07967_ _07974_ VGND VGND VPWR VPWR _07975_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17618_ net413 net335 VGND VGND VPWR VPWR _09605_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18598_ _10499_ _10500_ _10576_ VGND VGND VPWR VPWR _10577_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17549_ _09518_ _09519_ _09534_ VGND VGND VPWR VPWR _09536_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_47_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20560_ _12401_ _12402_ _12408_ VGND VGND VPWR VPWR _12409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19219_ _11166_ _11167_ VGND VGND VPWR VPWR _11168_ sky130_fd_sc_hd__nand2_1
X_20491_ _11438_ _12335_ _12336_ _12339_ VGND VGND VPWR VPWR _12340_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_41_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22230_ _01782_ _01786_ _01789_ _01781_ _01790_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__o32a_1
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22161_ _01229_ _01242_ _01245_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21112_ _12880_ _12955_ _12943_ VGND VGND VPWR VPWR _12958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22092_ _01619_ _01628_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout202 net203 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlymetal6s2s_1
X_25920_ _05436_ _05129_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__nand2_1
Xfanout213 net214 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_4
X_21043_ net756 _12034_ _12037_ _12889_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__a31o_1
Xfanout224 top0.cordic0.vec\[0\]\[16\] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__buf_2
Xfanout235 net236 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_4
Xfanout246 net247 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__buf_2
Xfanout257 top0.cordic0.vec\[0\]\[9\] VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__buf_4
X_25851_ top0.matmul0.beta_pass\[6\] _05071_ _05065_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__a21o_1
Xfanout268 top0.cordic0.vec\[0\]\[7\] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__buf_2
XFILLER_0_199_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout279 top0.cordic0.vec\[0\]\[5\] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__buf_2
XFILLER_0_158_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24802_ top0.matmul0.matmul_stage_inst.mult2\[5\] _04154_ _03642_ VGND VGND VPWR
+ VPWR _04155_ sky130_fd_sc_hd__mux2_1
X_22994_ _06277_ _02500_ net172 VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__o21ai_1
X_25782_ _05013_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_198_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24733_ _04000_ _04084_ _04085_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__a21o_2
XFILLER_0_9_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21945_ net165 _01503_ _01504_ net145 _01506_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_69_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24664_ _03252_ _03825_ _03875_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__a21o_1
X_21876_ net151 _01122_ _01299_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23615_ _02974_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__clkbuf_1
X_26403_ clknet_leaf_98_clk_sys _00044_ net588 VGND VGND VPWR VPWR top0.kpd\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20827_ _12228_ _12229_ _12240_ _12233_ VGND VGND VPWR VPWR _12676_ sky130_fd_sc_hd__a31o_1
X_24595_ _03820_ _03838_ _03949_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_181_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23546_ _02939_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__clkbuf_1
X_26334_ spi0.data_packed\[65\] spi0.data_packed\[66\] net695 VGND VGND VPWR VPWR
+ _05399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20758_ net300 net285 _12554_ net302 VGND VGND VPWR VPWR _12607_ sky130_fd_sc_hd__a211o_1
XFILLER_0_135_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26265_ _05364_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23477_ net1001 top0.matmul0.sin\[8\] _05461_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__mux2_1
X_20689_ _12427_ _12457_ VGND VGND VPWR VPWR _12538_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25216_ _04371_ _04560_ _04562_ _04518_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13230_ top0.pid_q.state\[0\] top0.pid_d.iterate_enable net1019 VGND VGND VPWR VPWR
+ _05451_ sky130_fd_sc_hd__and3_1
X_22428_ _01951_ _01984_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26196_ spi0.data_packed\[13\] _05328_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__xor2_1
XFILLER_0_165_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25147_ _04371_ _04174_ _04039_ _04493_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22359_ _01217_ net114 VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25078_ _04349_ _04425_ _04426_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__a21o_1
X_24029_ _03385_ _03386_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__xnor2_2
X_16920_ _08977_ _08978_ VGND VGND VPWR VPWR _08980_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16851_ top0.currT_r\[2\] _08903_ top0.matmul0.beta_pass\[2\] VGND VGND VPWR VPWR
+ _08915_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_102_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15802_ _07898_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__clkbuf_1
X_19570_ top0.cordic0.slte0.opB\[5\] top0.cordic0.slte0.opA\[5\] VGND VGND VPWR VPWR
+ _11459_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16782_ top0.kiq\[1\] _08863_ _08861_ VGND VGND VPWR VPWR _08864_ sky130_fd_sc_hd__and3_1
X_13994_ net33 _05475_ _05476_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18521_ _10499_ _10500_ VGND VGND VPWR VPWR _10501_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15733_ _07725_ _07730_ _07829_ VGND VGND VPWR VPWR _07830_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_32_clk_sys clknet_3_6__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_32_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18452_ _10429_ _10430_ VGND VGND VPWR VPWR _10432_ sky130_fd_sc_hd__or2_1
X_15664_ _07656_ _07761_ VGND VGND VPWR VPWR _07762_ sky130_fd_sc_hd__xor2_1
XFILLER_0_197_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17403_ _09344_ _09349_ _09389_ VGND VGND VPWR VPWR _09390_ sky130_fd_sc_hd__a21oi_1
X_14615_ _06759_ _06784_ VGND VGND VPWR VPWR _06820_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18383_ _10348_ _10363_ VGND VGND VPWR VPWR _10364_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15595_ _07688_ _07690_ _07692_ _07693_ VGND VGND VPWR VPWR _07694_ sky130_fd_sc_hd__and4_2
XFILLER_0_200_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17334_ top0.matmul0.matmul_stage_inst.mult1\[13\] top0.matmul0.matmul_stage_inst.mult2\[13\]
+ VGND VGND VPWR VPWR _09324_ sky130_fd_sc_hd__xor2_1
XFILLER_0_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14546_ _06649_ _06725_ _06713_ VGND VGND VPWR VPWR _06752_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_139_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17265_ _09263_ _09259_ _09264_ VGND VGND VPWR VPWR _09265_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_71_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14477_ _06672_ _06673_ _06608_ VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__o21a_1
XFILLER_0_125_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19004_ _10854_ _10855_ _10977_ VGND VGND VPWR VPWR _10978_ sky130_fd_sc_hd__o21a_1
X_16216_ _08220_ _08180_ _08306_ VGND VGND VPWR VPWR _08308_ sky130_fd_sc_hd__or3_1
X_13428_ net61 _05625_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__xnor2_1
X_17196_ top0.pid_q.state\[5\] _08479_ _09205_ net554 _09009_ VGND VGND VPWR VPWR
+ _09206_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13359_ net42 _05484_ _05486_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16147_ top0.pid_q.curr_int\[6\] _08239_ VGND VGND VPWR VPWR _08240_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16078_ _08169_ _08170_ VGND VGND VPWR VPWR _08171_ sky130_fd_sc_hd__xnor2_1
X_19906_ _11778_ _11771_ _11772_ VGND VGND VPWR VPWR _11780_ sky130_fd_sc_hd__and3_1
X_15029_ _07143_ VGND VGND VPWR VPWR _07144_ sky130_fd_sc_hd__clkbuf_4
X_19837_ _11632_ _11560_ VGND VGND VPWR VPWR _11715_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput2 rstb VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19768_ _11433_ VGND VGND VPWR VPWR _11651_ sky130_fd_sc_hd__buf_1
XFILLER_0_78_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18719_ net377 net314 VGND VGND VPWR VPWR _10696_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19699_ _11584_ VGND VGND VPWR VPWR _11585_ sky130_fd_sc_hd__inv_2
X_21730_ net123 net108 VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__xor2_2
XFILLER_0_148_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21661_ _01221_ _01222_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__nand2_4
XFILLER_0_46_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23400_ _01065_ _02810_ _02815_ _02817_ _02839_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__o2111a_1
X_20612_ _12458_ _12459_ _12427_ VGND VGND VPWR VPWR _12461_ sky130_fd_sc_hd__a21o_1
X_24380_ _03170_ _03171_ _03192_ _03174_ VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_47_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21592_ _01088_ _01090_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__xor2_2
XFILLER_0_188_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23331_ _02755_ _02764_ _02775_ VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__a21oi_1
X_20543_ _12389_ _12391_ _12280_ VGND VGND VPWR VPWR _12392_ sky130_fd_sc_hd__mux2_1
X_26050_ top0.a_in_matmul\[4\] _05239_ _05230_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__mux2_1
X_23262_ net228 net223 net203 VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__mux2_1
X_20474_ _12314_ _12322_ VGND VGND VPWR VPWR _12323_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25001_ _04349_ _04350_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__xnor2_1
X_22213_ _01755_ _01773_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23193_ _05719_ _06971_ _02648_ net790 VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__a22o_1
XFILLER_0_160_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22144_ net155 _01701_ _01704_ _01705_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__a211o_2
XFILLER_0_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26952_ clknet_leaf_16_clk_sys _00569_ net613 VGND VGND VPWR VPWR top0.matmul0.b\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_22075_ _01629_ _01636_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__xnor2_4
X_25903_ top0.matmul0.alpha_pass\[10\] VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__inv_2
X_21026_ _12683_ _12871_ _12872_ _11789_ VGND VGND VPWR VPWR _12873_ sky130_fd_sc_hd__a211oi_4
X_26883_ clknet_leaf_39_clk_sys _00500_ net683 VGND VGND VPWR VPWR top0.svm0.tB\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25834_ _05050_ _05051_ _05054_ _05053_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22977_ _02485_ _02480_ net170 VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__o21ba_1
X_25765_ _05003_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__clkbuf_1
X_24716_ _04068_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__clkbuf_8
X_21928_ net130 _01487_ _01488_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__and3_1
X_25696_ top0.matmul0.matmul_stage_inst.c\[15\] _04896_ _04960_ VGND VGND VPWR VPWR
+ _04962_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24647_ _03883_ _03884_ _03885_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__a21o_1
X_21859_ _01418_ _01409_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14400_ _06603_ _06607_ VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15380_ _07476_ _07459_ _07478_ VGND VGND VPWR VPWR _07479_ sky130_fd_sc_hd__nor3b_1
X_24578_ _03713_ _03708_ _03775_ _03776_ _03778_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_92_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14331_ _06536_ _06540_ VGND VGND VPWR VPWR _06541_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26317_ _05390_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23529_ _02930_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__clkbuf_1
X_27297_ clknet_3_1__leaf_clk_mosi _00911_ VGND VGND VPWR VPWR spi0.opcode\[3\] sky130_fd_sc_hd__dfxtp_1
X_14262_ _06387_ _06472_ VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__xnor2_2
X_17050_ _09099_ VGND VGND VPWR VPWR _09100_ sky130_fd_sc_hd__clkbuf_4
X_26248_ spi0.data_packed\[22\] spi0.data_packed\[23\] net698 VGND VGND VPWR VPWR
+ _05356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13213_ _05438_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__buf_4
X_16001_ net529 net446 VGND VGND VPWR VPWR _08095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14193_ net51 _05726_ _05727_ VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__and3_1
X_26179_ spi0.data_packed\[9\] _05315_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17952_ _09936_ _09937_ VGND VGND VPWR VPWR _09938_ sky130_fd_sc_hd__xnor2_1
X_16903_ top0.pid_q.curr_error\[5\] _08951_ top0.pid_q.prev_error\[5\] VGND VGND VPWR
+ VPWR _08964_ sky130_fd_sc_hd__a21o_1
X_17883_ net426 net313 VGND VGND VPWR VPWR _09870_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19622_ _11510_ VGND VGND VPWR VPWR _11511_ sky130_fd_sc_hd__buf_6
X_16834_ _05601_ VGND VGND VPWR VPWR _08899_ sky130_fd_sc_hd__buf_2
XFILLER_0_73_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19553_ _11440_ _11441_ _11419_ VGND VGND VPWR VPWR _11442_ sky130_fd_sc_hd__mux2_1
X_16765_ _08789_ _08787_ _08839_ VGND VGND VPWR VPWR _08849_ sky130_fd_sc_hd__mux2_2
X_13977_ net1025 _05723_ _05724_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__and3_1
X_18504_ net341 _10458_ _10388_ VGND VGND VPWR VPWR _10484_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_87_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15716_ net474 net512 VGND VGND VPWR VPWR _07813_ sky130_fd_sc_hd__nand2_2
X_19484_ top0.pid_d.curr_int\[11\] top0.pid_d.prev_int\[11\] VGND VGND VPWR VPWR _11378_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16696_ _08755_ _08780_ VGND VGND VPWR VPWR _08781_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18435_ _10411_ _10414_ VGND VGND VPWR VPWR _10416_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15647_ _07650_ _07651_ _07744_ VGND VGND VPWR VPWR _07745_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_158_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18366_ net396 _09518_ _09399_ _10074_ VGND VGND VPWR VPWR _10347_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15578_ _07660_ _07676_ VGND VGND VPWR VPWR _07677_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17317_ _09309_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__clkbuf_1
X_14529_ _06727_ _06735_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18297_ net1023 net391 VGND VGND VPWR VPWR _10279_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17248_ top0.matmul0.matmul_stage_inst.mult1\[0\] top0.matmul0.matmul_stage_inst.mult2\[0\]
+ VGND VGND VPWR VPWR _09251_ sky130_fd_sc_hd__xor2_1
XFILLER_0_141_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17179_ top0.pid_q.curr_int\[7\] _09141_ _09190_ _09136_ VGND VGND VPWR VPWR _00220_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20190_ net259 net255 VGND VGND VPWR VPWR _12039_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_45_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22900_ _02324_ top0.svm0.tC\[6\] _02417_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23880_ _02981_ _03017_ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__nor2_2
X_22831_ _02346_ _02348_ _02349_ _02350_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__or4_1
XFILLER_0_155_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25550_ top0.matmul0.b\[14\] top0.matmul0.matmul_stage_inst.f\[14\] _04856_ VGND
+ VGND VPWR VPWR _04862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22762_ top0.pid_q.prev_int\[6\] _02292_ _02295_ top0.pid_q.curr_int\[6\] VGND VGND
+ VPWR VPWR _00425_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24501_ _03856_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__clkbuf_1
X_21713_ _01267_ _01271_ _01272_ _01274_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__a31o_1
X_25481_ _04821_ _04755_ _04764_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22693_ net78 net99 net91 _01221_ _01937_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__o32a_1
XFILLER_0_13_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27220_ clknet_3_5__leaf_clk_mosi _00834_ VGND VGND VPWR VPWR spi0.data_packed\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_24432_ _03784_ _03785_ _03786_ _03787_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21644_ net138 _01105_ VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24363_ _03196_ _03197_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__or2_2
X_27151_ clknet_leaf_11_clk_sys _00765_ net601 VGND VGND VPWR VPWR top0.a_in_matmul\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_40 top0.c_out_calc\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21575_ net139 _01135_ _01136_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26102_ top0.periodTop\[1\] _05276_ _05278_ net62 VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__a22o_1
X_23314_ net150 _02717_ _02718_ net145 VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27082_ clknet_leaf_20_clk_sys _00699_ net609 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_20526_ _12373_ _12374_ VGND VGND VPWR VPWR _12375_ sky130_fd_sc_hd__xnor2_1
X_24294_ _03647_ _03648_ _03649_ _03650_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23245_ _02692_ _02694_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__xnor2_2
X_26033_ top0.matmul0.alpha_pass\[1\] _05203_ _05225_ VGND VGND VPWR VPWR _05226_
+ sky130_fd_sc_hd__a21o_1
X_20457_ net280 _12287_ _12300_ _12304_ _12305_ VGND VGND VPWR VPWR _12306_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23176_ _05717_ _07034_ _02644_ net908 VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__a22o_1
X_20388_ net214 _12165_ VGND VGND VPWR VPWR _12237_ sky130_fd_sc_hd__nand2_1
Xclkbuf_3_0__f_clk_mosi clknet_0_clk_mosi VGND VGND VPWR VPWR clknet_3_0__leaf_clk_mosi
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_112_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22127_ _11444_ _01687_ _01688_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22058_ _01558_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__inv_2
X_26935_ clknet_leaf_3_clk_sys _00552_ net583 VGND VGND VPWR VPWR top0.matmul0.cos\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13900_ net33 _05478_ _05479_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__and3_1
X_21009_ net229 _12852_ _12854_ _12855_ VGND VGND VPWR VPWR _12856_ sky130_fd_sc_hd__a31o_1
X_26866_ clknet_leaf_41_clk_sys _00483_ net683 VGND VGND VPWR VPWR top0.svm0.tA\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_14880_ spi0.data_packed\[48\] top0.kpq\[0\] _07053_ VGND VGND VPWR VPWR _07060_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25817_ top0.matmul0.alpha_pass\[1\] top0.matmul0.beta_pass\[1\] VGND VGND VPWR VPWR
+ _05042_ sky130_fd_sc_hd__and2_1
X_13831_ _06041_ _06043_ _06036_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__o21a_1
XFILLER_0_173_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26797_ clknet_leaf_105_clk_sys _00414_ net576 VGND VGND VPWR VPWR top0.cordic0.gm0.iter\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_98_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16550_ net456 net497 VGND VGND VPWR VPWR _08637_ sky130_fd_sc_hd__nand2_2
XFILLER_0_97_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13762_ net1027 _05484_ _05486_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__and3_1
X_25748_ top0.matmul0.matmul_stage_inst.a\[2\] _04889_ _05458_ VGND VGND VPWR VPWR
+ _04995_ sky130_fd_sc_hd__mux2_1
X_15501_ _07298_ _07599_ VGND VGND VPWR VPWR _07600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16481_ _08500_ _08505_ _08568_ VGND VGND VPWR VPWR _08569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13693_ _05881_ _05904_ _05905_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__a21bo_1
X_25679_ top0.matmul0.sin\[10\] _04942_ _04884_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__o21a_1
X_18220_ net354 net358 VGND VGND VPWR VPWR _10203_ sky130_fd_sc_hd__nor2_2
XFILLER_0_66_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15432_ _07240_ _07529_ _07530_ VGND VGND VPWR VPWR _07531_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_150_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18151_ _10001_ _10005_ _10134_ VGND VGND VPWR VPWR _10135_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15363_ net482 _07461_ VGND VGND VPWR VPWR _07462_ sky130_fd_sc_hd__nand2_1
X_17102_ net820 _09115_ _09127_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__a21o_1
X_14314_ _06421_ _06423_ _06422_ VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__o21ba_1
X_18082_ net1019 VGND VGND VPWR VPWR _10067_ sky130_fd_sc_hd__clkbuf_4
X_15294_ net542 net464 VGND VGND VPWR VPWR _07393_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17033_ _09081_ top0.currT_r\[14\] _08900_ top0.currT_r\[13\] _05662_ VGND VGND VPWR
+ VPWR _09085_ sky130_fd_sc_hd__a2111o_1
X_14245_ net56 _06135_ VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14176_ _06178_ _06384_ _06386_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_0_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18984_ _10955_ _10957_ VGND VGND VPWR VPWR _10958_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17935_ net342 net383 VGND VGND VPWR VPWR _09921_ sky130_fd_sc_hd__nand2_1
XFILLER_0_178_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17866_ net404 net336 net399 net339 VGND VGND VPWR VPWR _09853_ sky130_fd_sc_hd__a22oi_1
X_16817_ top0.currT_r\[0\] _08883_ VGND VGND VPWR VPWR _08884_ sky130_fd_sc_hd__xnor2_1
X_19605_ top0.cordic0.slte0.opA\[9\] VGND VGND VPWR VPWR _11494_ sky130_fd_sc_hd__inv_2
X_17797_ top0.pid_d.mult0.a\[3\] net326 VGND VGND VPWR VPWR _09784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19536_ _11425_ VGND VGND VPWR VPWR _11426_ sky130_fd_sc_hd__buf_4
X_16748_ _08142_ _08721_ _08753_ VGND VGND VPWR VPWR _08832_ sky130_fd_sc_hd__nor3_1
XFILLER_0_88_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19467_ net441 _11361_ _11362_ _11220_ VGND VGND VPWR VPWR _11363_ sky130_fd_sc_hd__a31o_1
XFILLER_0_186_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16679_ _08701_ _08702_ _08763_ VGND VGND VPWR VPWR _08764_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_124_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18418_ _10364_ _10398_ VGND VGND VPWR VPWR _10399_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19398_ top0.pid_d.curr_int\[1\] top0.pid_d.prev_int\[1\] top0.pid_d.prev_int\[0\]
+ top0.pid_d.curr_int\[0\] VGND VGND VPWR VPWR _11302_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_174_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18349_ _10325_ _10328_ VGND VGND VPWR VPWR _10331_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21360_ _00916_ _00927_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20311_ _12155_ _12158_ VGND VGND VPWR VPWR _12160_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21291_ _13121_ _13133_ VGND VGND VPWR VPWR _13134_ sky130_fd_sc_hd__xnor2_2
X_23030_ _02526_ _02530_ top0.svm0.delta\[15\] VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20242_ net264 _12066_ _12089_ _12065_ _12090_ VGND VGND VPWR VPWR _12091_ sky130_fd_sc_hd__a221o_2
XFILLER_0_3_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20173_ top0.pid_d.out_valid _12016_ _12018_ _12020_ _12024_ VGND VGND VPWR VPWR
+ _12025_ sky130_fd_sc_hd__o221a_1
XFILLER_0_110_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24981_ _04251_ _04325_ _04330_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26720_ clknet_leaf_82_clk_sys _00337_ net638 VGND VGND VPWR VPWR top0.pid_d.curr_int\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_23932_ _03087_ _03289_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_157_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26651_ clknet_leaf_75_clk_sys _00268_ net639 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_23863_ _03218_ _03219_ _03214_ _03215_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25602_ net747 _00000_ _04892_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__o21a_1
X_22814_ top0.svm0.counter\[8\] top0.svm0.tA\[8\] VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__nand2_1
X_26582_ clknet_leaf_53_clk_sys _00205_ net674 VGND VGND VPWR VPWR top0.pid_q.prev_error\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_23794_ _03150_ _03151_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__nor2_2
XFILLER_0_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25533_ top0.matmul0.b\[6\] top0.matmul0.matmul_stage_inst.f\[6\] _04846_ VGND VGND
+ VPWR VPWR _04853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22745_ net176 _11558_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_79_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_79_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_181_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25464_ _04801_ _04806_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__xnor2_2
X_22676_ _02182_ _02183_ _02171_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27203_ clknet_leaf_91_clk_sys _00817_ net599 VGND VGND VPWR VPWR top0.cordic0.slte0.opB\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_24415_ _03769_ _03770_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__xor2_1
X_21627_ _01154_ _01146_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__xor2_1
XFILLER_0_191_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25395_ _04732_ _04738_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_152_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27134_ clknet_leaf_11_clk_sys _00748_ net601 VGND VGND VPWR VPWR top0.matmul0.op_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24346_ _03202_ _03203_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21558_ _01118_ _01119_ net119 VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20509_ _12261_ _12324_ VGND VGND VPWR VPWR _12358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24277_ _03290_ _03629_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__xor2_1
X_27065_ clknet_leaf_0_clk_sys _00682_ net586 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.c\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_21489_ _01023_ _01049_ _01051_ _01052_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__o31a_1
XFILLER_0_160_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14030_ net64 _06131_ _06148_ _06149_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26016_ top0.pid_q.out\[13\] _05198_ _05199_ spi0.data_packed\[61\] VGND VGND VPWR
+ VPWR _05213_ sky130_fd_sc_hd__a22o_1
X_23228_ _02676_ _02677_ net1016 VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23159_ _07115_ _02308_ _02642_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15981_ top0.pid_q.curr_int\[3\] VGND VGND VPWR VPWR _08076_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17720_ net385 _09706_ _09362_ _09433_ VGND VGND VPWR VPWR _09707_ sky130_fd_sc_hd__or4_1
X_14932_ _07087_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__clkbuf_1
X_26918_ clknet_leaf_1_clk_sys _00535_ net582 VGND VGND VPWR VPWR top0.matmul0.sin\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_145_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17651_ net388 net378 net359 VGND VGND VPWR VPWR _09638_ sky130_fd_sc_hd__o21a_1
X_26849_ clknet_leaf_44_clk_sys _00466_ net686 VGND VGND VPWR VPWR top0.svm0.delta\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_14863_ spi0.data_packed\[72\] top0.kpd\[8\] _07042_ VGND VGND VPWR VPWR _07051_
+ sky130_fd_sc_hd__mux2_1
X_16602_ _08599_ _08676_ VGND VGND VPWR VPWR _08688_ sky130_fd_sc_hd__nand2_1
X_13814_ net59 _05496_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__nand2_1
X_17582_ net415 _09567_ _09568_ VGND VGND VPWR VPWR _09569_ sky130_fd_sc_hd__a21oi_1
X_14794_ _06943_ _06994_ VGND VGND VPWR VPWR _06995_ sky130_fd_sc_hd__or2_1
XFILLER_0_159_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19321_ _11259_ _11260_ net437 VGND VGND VPWR VPWR _11261_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_35_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16533_ net13 _08618_ _08619_ VGND VGND VPWR VPWR _08620_ sky130_fd_sc_hd__a21bo_1
X_13745_ _05956_ _05957_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19252_ _11196_ _11197_ VGND VGND VPWR VPWR _11198_ sky130_fd_sc_hd__nand2_1
X_16464_ net1018 _08552_ VGND VGND VPWR VPWR _08553_ sky130_fd_sc_hd__and2_1
X_13676_ _05887_ _05888_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18203_ net350 net366 VGND VGND VPWR VPWR _10186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15415_ _07472_ _07510_ _07460_ _07465_ _07513_ VGND VGND VPWR VPWR _07514_ sky130_fd_sc_hd__o221a_1
XFILLER_0_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19183_ _11133_ _11134_ VGND VGND VPWR VPWR _11135_ sky130_fd_sc_hd__and2_1
X_16395_ top0.pid_q.out\[9\] top0.pid_q.curr_int\[9\] VGND VGND VPWR VPWR _08484_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18134_ _10116_ _10117_ VGND VGND VPWR VPWR _10118_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15346_ _07436_ _07437_ _07366_ VGND VGND VPWR VPWR _07445_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18065_ _10040_ _10049_ VGND VGND VPWR VPWR _10050_ sky130_fd_sc_hd__nand2_1
X_15277_ net479 _07371_ _07374_ _07375_ VGND VGND VPWR VPWR _07376_ sky130_fd_sc_hd__a31oi_4
Xhold107 top0.svm0.tC\[10\] VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold118 top0.pid_q.prev_error\[7\] VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__dlygate4sd3_1
X_17016_ _09065_ _09066_ _09067_ _09068_ VGND VGND VPWR VPWR _09069_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_22_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold129 _00127_ VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__dlygate4sd3_1
X_14228_ _06437_ _06438_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14159_ _06255_ _06272_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout609 net630 VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18967_ net373 net311 _10384_ _09965_ VGND VGND VPWR VPWR _10941_ sky130_fd_sc_hd__a211o_1
X_17918_ net336 net393 VGND VGND VPWR VPWR _09904_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18898_ _10864_ _10872_ VGND VGND VPWR VPWR _10873_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_179_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17849_ net332 net404 VGND VGND VPWR VPWR _09836_ sky130_fd_sc_hd__nand2_1
X_20860_ _12704_ _12706_ _12708_ VGND VGND VPWR VPWR _12709_ sky130_fd_sc_hd__nand3_1
XFILLER_0_88_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19519_ net196 VGND VGND VPWR VPWR _11409_ sky130_fd_sc_hd__inv_2
X_20791_ _12588_ _12639_ VGND VGND VPWR VPWR _12640_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_80_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_80_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22530_ _02007_ _02085_ _02084_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__a21o_1
XFILLER_0_158_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22461_ net111 _01211_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24200_ _03555_ _03557_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__xor2_1
XFILLER_0_161_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21412_ _00977_ _00978_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__or2_1
X_25180_ _04455_ _04526_ _04527_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__o21ai_1
X_22392_ _01939_ _01934_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__and2b_1
XFILLER_0_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24131_ _03482_ _03484_ _03486_ _03487_ _03488_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__o221a_2
X_21343_ _11789_ _13035_ VGND VGND VPWR VPWR _13185_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24062_ _03419_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21274_ net247 _13028_ VGND VGND VPWR VPWR _13117_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23013_ top0.svm0.delta\[13\] _02516_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__xor2_1
X_20225_ _12072_ _12073_ VGND VGND VPWR VPWR _12074_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20156_ net207 net206 net209 VGND VGND VPWR VPWR _12008_ sky130_fd_sc_hd__a21oi_1
X_24964_ _04303_ _04314_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__xnor2_2
X_20087_ _11426_ _11514_ VGND VGND VPWR VPWR _11947_ sky130_fd_sc_hd__nand2_1
X_26703_ clknet_leaf_83_clk_sys net875 net646 VGND VGND VPWR VPWR top0.pid_d.prev_error\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23915_ _03237_ _03242_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__nand2_1
X_24895_ _03959_ _04061_ _04245_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__nor3_1
XFILLER_0_170_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26634_ clknet_leaf_74_clk_sys _00251_ net637 VGND VGND VPWR VPWR top0.pid_d.out\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_23846_ _03202_ _03203_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26565_ clknet_leaf_53_clk_sys _00188_ net672 VGND VGND VPWR VPWR top0.pid_q.curr_error\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23777_ _03098_ _03134_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__nor2_1
X_20989_ net262 _12135_ VGND VGND VPWR VPWR _12836_ sky130_fd_sc_hd__nor2_1
XFILLER_0_178_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25516_ top0.matmul0.matmul_stage_inst.mult1\[14\] _04767_ _03148_ VGND VGND VPWR
+ VPWR _04844_ sky130_fd_sc_hd__mux2_1
X_13530_ _05700_ _05703_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__nor2_1
XFILLER_0_193_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22728_ _02257_ _02267_ _01877_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26496_ clknet_leaf_73_clk_sys _00119_ net655 VGND VGND VPWR VPWR top0.pid_d.prev_int\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13461_ _05661_ _05673_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__xor2_1
X_25447_ _04288_ _03936_ _04787_ _04788_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__a22o_1
X_22659_ _02181_ _02211_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_173_Right_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15200_ _07220_ _07298_ VGND VGND VPWR VPWR _07299_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_164_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16180_ net466 net503 VGND VGND VPWR VPWR _08272_ sky130_fd_sc_hd__nand2_1
X_25378_ _03900_ _03936_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__nand2_2
X_13392_ _05604_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__buf_4
XFILLER_0_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27117_ clknet_leaf_33_clk_sys _00731_ net665 VGND VGND VPWR VPWR top0.c_out_calc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_15131_ net521 VGND VGND VPWR VPWR _07230_ sky130_fd_sc_hd__inv_2
X_24329_ _03177_ _03179_ _03685_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__o21ai_2
X_27048_ clknet_leaf_17_clk_sys _00665_ net611 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.d\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_15062_ _07149_ _07160_ VGND VGND VPWR VPWR _07161_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14013_ _06222_ _06225_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__xnor2_2
X_19870_ net243 _11729_ _11745_ VGND VGND VPWR VPWR _11746_ sky130_fd_sc_hd__o21ai_1
X_18821_ net323 _10792_ _10793_ _10794_ _10796_ VGND VGND VPWR VPWR _10797_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18752_ _10725_ _10726_ VGND VGND VPWR VPWR _10729_ sky130_fd_sc_hd__and2_1
X_15964_ _08053_ _08058_ VGND VGND VPWR VPWR _08059_ sky130_fd_sc_hd__xnor2_2
X_17703_ net385 _09687_ _09689_ net352 VGND VGND VPWR VPWR _09690_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14915_ _07078_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18683_ net309 _10526_ _10659_ _09351_ VGND VGND VPWR VPWR _10661_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_198_Left_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15895_ _07905_ _07990_ VGND VGND VPWR VPWR _07991_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17634_ net403 net342 VGND VGND VPWR VPWR _09621_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14846_ _07041_ VGND VGND VPWR VPWR _07042_ sky130_fd_sc_hd__buf_4
XFILLER_0_59_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17565_ net418 net354 VGND VGND VPWR VPWR _09552_ sky130_fd_sc_hd__nand2_1
X_14777_ net31 _06867_ VGND VGND VPWR VPWR _06978_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19304_ top0.matmul0.alpha_pass\[13\] _11241_ VGND VGND VPWR VPWR _11245_ sky130_fd_sc_hd__or2_1
X_16516_ _08489_ _08603_ _08490_ VGND VGND VPWR VPWR _08604_ sky130_fd_sc_hd__a21oi_1
X_13728_ _05937_ _05940_ VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17496_ net417 net333 VGND VGND VPWR VPWR _09483_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19235_ net336 _11117_ _11179_ _11182_ _08889_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__o221a_1
X_16447_ _08220_ _08535_ VGND VGND VPWR VPWR _08536_ sky130_fd_sc_hd__xnor2_1
X_13659_ _05869_ _05870_ _05871_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19166_ _11119_ VGND VGND VPWR VPWR _11120_ sky130_fd_sc_hd__buf_2
X_16378_ _08386_ VGND VGND VPWR VPWR _08468_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18117_ _10099_ _10100_ VGND VGND VPWR VPWR _10101_ sky130_fd_sc_hd__xnor2_1
X_15329_ _07391_ _07395_ VGND VGND VPWR VPWR _07428_ sky130_fd_sc_hd__xor2_1
XFILLER_0_147_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19097_ _11003_ _11010_ VGND VGND VPWR VPWR _11069_ sky130_fd_sc_hd__nand2_1
X_18048_ _09903_ _09904_ _10032_ VGND VGND VPWR VPWR _10033_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_112_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_27_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_27_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout406 top0.pid_d.mult0.a\[5\] VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__dlymetal6s2s_1
X_20010_ _11612_ net190 VGND VGND VPWR VPWR _11876_ sky130_fd_sc_hd__nor2_1
Xfanout417 top0.pid_d.mult0.a\[3\] VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__buf_4
Xfanout428 top0.matmul0.beta_pass\[14\] VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__clkbuf_4
Xfanout439 net440 VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__buf_2
X_19999_ top0.cordic0.slte0.opA\[4\] net10 VGND VGND VPWR VPWR _11866_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21961_ _01521_ _01522_ _01518_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__o21a_1
X_23700_ net556 top0.matmul0.matmul_stage_inst.c\[3\] top0.matmul0.matmul_stage_inst.b\[3\]
+ net568 VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__a22o_2
X_20912_ net291 _12756_ _12759_ VGND VGND VPWR VPWR _12760_ sky130_fd_sc_hd__a21oi_2
X_24680_ _03921_ _03922_ _03924_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__a21boi_2
X_21892_ _01432_ _01453_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23631_ _02988_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__clkbuf_4
X_20843_ _11593_ _12040_ VGND VGND VPWR VPWR _12692_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_202_Left_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout13 net75 VGND VGND VPWR VPWR net1024 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26350_ spi0.data_packed\[73\] spi0.data_packed\[74\] net690 VGND VGND VPWR VPWR
+ _05407_ sky130_fd_sc_hd__mux2_1
X_23562_ _02947_ VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__clkbuf_1
X_20774_ net295 net278 VGND VGND VPWR VPWR _12623_ sky130_fd_sc_hd__and2_1
Xfanout24 top0.periodTop_r\[15\] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
Xfanout35 top0.periodTop_r\[12\] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25301_ _04411_ _04573_ _04646_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__o21a_1
Xfanout46 net47 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout57 net58 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22513_ _02060_ _02068_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__xor2_2
Xfanout68 top0.periodTop_r\[0\] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_4
X_26281_ net954 VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__clkbuf_1
X_23493_ _02911_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout79 net80 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25232_ _04508_ _04577_ _04578_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__a21oi_1
X_22444_ _01809_ _01891_ _02000_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25163_ _04443_ _04445_ _04441_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__a21o_1
X_22375_ _01899_ _01933_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24114_ _03458_ _03457_ _03459_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__o21a_1
X_21326_ _13162_ _13167_ _13125_ VGND VGND VPWR VPWR _13168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25094_ _04355_ _04357_ _04442_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24045_ _03384_ _03401_ _03402_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__o21ba_1
X_21257_ _12965_ _13007_ VGND VGND VPWR VPWR _13101_ sky130_fd_sc_hd__nor2_1
X_20208_ net296 net289 VGND VGND VPWR VPWR _12057_ sky130_fd_sc_hd__nand2b_2
X_21188_ _13030_ _13031_ VGND VGND VPWR VPWR _13032_ sky130_fd_sc_hd__xor2_1
X_20139_ _11967_ _11968_ top0.cordic0.slte0.opA\[14\] VGND VGND VPWR VPWR _11995_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25996_ _05197_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__clkbuf_1
X_24947_ _04295_ _04297_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__xnor2_1
X_14700_ _06865_ _06903_ VGND VGND VPWR VPWR _06904_ sky130_fd_sc_hd__and2_1
X_15680_ _07718_ _07777_ VGND VGND VPWR VPWR _07778_ sky130_fd_sc_hd__xnor2_1
X_24878_ _04114_ _04115_ _04227_ _04228_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__o22a_1
XFILLER_0_169_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14631_ _06834_ _06835_ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__or2b_1
X_26617_ clknet_leaf_28_clk_sys _00234_ net621 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_23829_ _03015_ _03016_ _03029_ _03030_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__o22a_1
XFILLER_0_157_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17350_ top0.matmul0.beta_pass\[15\] _09337_ net562 VGND VGND VPWR VPWR _09338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14562_ net36 _05723_ _05724_ VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__and3_1
X_26548_ clknet_leaf_49_clk_sys _00171_ net675 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16301_ _08254_ _08311_ _08391_ VGND VGND VPWR VPWR _08392_ sky130_fd_sc_hd__o21ai_1
X_13513_ _05663_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__clkbuf_4
X_17281_ top0.matmul0.beta_pass\[5\] _09278_ net562 VGND VGND VPWR VPWR _09279_ sky130_fd_sc_hd__mux2_1
X_14493_ net44 _06131_ VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__nand2_1
X_26479_ clknet_leaf_11_clk_sys _00110_ net604 VGND VGND VPWR VPWR top0.periodTop\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_19020_ _10930_ _10979_ _10980_ VGND VGND VPWR VPWR _10993_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_125_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16232_ _08323_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__clkbuf_1
X_13444_ net60 VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16163_ _07320_ net444 VGND VGND VPWR VPWR _08255_ sky130_fd_sc_hd__nand2_2
X_13375_ _05587_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15114_ net462 net464 VGND VGND VPWR VPWR _07213_ sky130_fd_sc_hd__and2_4
X_16094_ net526 net446 VGND VGND VPWR VPWR _08187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15045_ net815 _07139_ _07143_ top0.pid_d.curr_int\[15\] VGND VGND VPWR VPWR _00132_
+ sky130_fd_sc_hd__a22o_1
X_19922_ net220 _11784_ _11793_ VGND VGND VPWR VPWR _11795_ sky130_fd_sc_hd__or3_1
X_19853_ _11451_ VGND VGND VPWR VPWR _11730_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18804_ _10690_ net360 _10779_ VGND VGND VPWR VPWR _10780_ sky130_fd_sc_hd__a21o_1
X_16996_ net551 _09050_ _08881_ VGND VGND VPWR VPWR _09051_ sky130_fd_sc_hd__a21o_1
X_19784_ net266 _11643_ VGND VGND VPWR VPWR _11666_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15947_ net477 net505 VGND VGND VPWR VPWR _08042_ sky130_fd_sc_hd__nand2_1
X_18735_ net323 net368 VGND VGND VPWR VPWR _10712_ sky130_fd_sc_hd__nand2_2
XFILLER_0_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18666_ _09377_ _10643_ net364 VGND VGND VPWR VPWR _10644_ sky130_fd_sc_hd__o21a_1
X_15878_ _07969_ _07973_ VGND VGND VPWR VPWR _07974_ sky130_fd_sc_hd__xor2_1
XFILLER_0_153_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14829_ net851 _06279_ _07028_ _05465_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17617_ net408 net337 VGND VGND VPWR VPWR _09604_ sky130_fd_sc_hd__nand2_1
X_18597_ _10499_ _10500_ _10493_ VGND VGND VPWR VPWR _10576_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17548_ _09518_ _09519_ _09528_ _09534_ VGND VGND VPWR VPWR _09535_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17479_ _09357_ _09428_ VGND VGND VPWR VPWR _09466_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19218_ top0.pid_d.prev_error\[5\] top0.pid_d.curr_error\[5\] VGND VGND VPWR VPWR
+ _11167_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20490_ net289 _12061_ _12338_ net304 net301 VGND VGND VPWR VPWR _12339_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19149_ top0.kid\[9\] _11098_ _11100_ top0.kpd\[9\] VGND VGND VPWR VPWR _11110_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22160_ _01695_ _01721_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21111_ _12943_ _12878_ _12955_ _12956_ VGND VGND VPWR VPWR _12957_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_160_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22091_ _01650_ _01651_ _01652_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__a21o_1
Xfanout203 net204 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_4
X_21042_ _12740_ _12888_ VGND VGND VPWR VPWR _12889_ sky130_fd_sc_hd__nor2_1
Xfanout214 top0.cordic0.vec\[0\]\[17\] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__buf_4
XFILLER_0_10_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout225 net226 VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_4
Xfanout236 net237 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_4
Xfanout247 net248 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_2
X_25850_ top0.matmul0.alpha_pass\[4\] top0.matmul0.alpha_pass\[5\] top0.matmul0.beta_pass\[4\]
+ _05063_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__or4_1
Xfanout258 net261 VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__buf_4
XFILLER_0_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout269 net270 VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__buf_4
XFILLER_0_157_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24801_ _04064_ _04153_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_199_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25781_ net205 _12019_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__nor2_2
XFILLER_0_198_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22993_ top0.svm0.delta\[10\] _02499_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__xor2_1
X_24732_ _04003_ _04004_ _04082_ _04083_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__o22a_1
X_21944_ _01311_ _01505_ _01267_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24663_ _04013_ _04016_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__xnor2_1
X_21875_ _01412_ _01436_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__xnor2_1
X_26402_ clknet_leaf_98_clk_sys _00043_ net589 VGND VGND VPWR VPWR top0.kpd\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23614_ top0.matmul0.alpha_pass\[14\] _09331_ net561 VGND VGND VPWR VPWR _02974_
+ sky130_fd_sc_hd__mux2_1
X_20826_ _12244_ _12674_ VGND VGND VPWR VPWR _12675_ sky130_fd_sc_hd__and2_2
X_24594_ _03820_ _03838_ _03816_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__a21o_1
XFILLER_0_166_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26333_ _05398_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__clkbuf_1
X_23545_ top0.a_in_matmul\[12\] top0.matmul0.a\[12\] _02937_ VGND VGND VPWR VPWR _02939_
+ sky130_fd_sc_hd__mux2_1
X_20757_ _12583_ _12605_ VGND VGND VPWR VPWR _12606_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26264_ spi0.data_packed\[30\] spi0.data_packed\[31\] net696 VGND VGND VPWR VPWR
+ _05364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20688_ _12427_ _12457_ VGND VGND VPWR VPWR _12537_ sky130_fd_sc_hd__or2_1
X_23476_ _02902_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25215_ _04371_ _04561_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__nor2_1
X_22427_ _01951_ _01984_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26195_ spi0.data_packed\[11\] spi0.data_packed\[12\] _05321_ net18 VGND VGND VPWR
+ VPWR _05328_ sky130_fd_sc_hd__a31o_1
X_25146_ _04039_ _04493_ _04371_ _04174_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22358_ _01062_ _01777_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_14_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21309_ net738 _12034_ _12037_ _13151_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__a31o_1
X_25077_ _03496_ _03826_ _04350_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__and3_1
X_22289_ net90 net86 VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__nand2_1
X_24028_ _03380_ _03381_ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__xnor2_1
Xhold290 top0.pid_d.prev_int\[9\] VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__dlygate4sd3_1
X_16850_ _08882_ _08907_ _08913_ _08914_ _08889_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__o311a_1
XFILLER_0_102_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15801_ _07800_ _07897_ VGND VGND VPWR VPWR _07898_ sky130_fd_sc_hd__and2_1
X_16781_ _05448_ VGND VGND VPWR VPWR _08863_ sky130_fd_sc_hd__clkbuf_2
X_13993_ net30 _05478_ _05479_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__and3_1
X_25979_ _05184_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18520_ net410 _09460_ _10228_ VGND VGND VPWR VPWR _10500_ sky130_fd_sc_hd__or3_1
XFILLER_0_137_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15732_ _07725_ _07730_ _07723_ VGND VGND VPWR VPWR _07829_ sky130_fd_sc_hd__o21a_1
X_18451_ _10429_ _10430_ VGND VGND VPWR VPWR _10431_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15663_ _07749_ _07760_ VGND VGND VPWR VPWR _07761_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_158_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17402_ _09387_ _09388_ VGND VGND VPWR VPWR _09389_ sky130_fd_sc_hd__xnor2_1
X_14614_ _06751_ _06790_ _06818_ VGND VGND VPWR VPWR _06819_ sky130_fd_sc_hd__a21o_1
XFILLER_0_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18382_ _10361_ _10362_ VGND VGND VPWR VPWR _10363_ sky130_fd_sc_hd__or2b_1
X_15594_ _07596_ _07691_ VGND VGND VPWR VPWR _07693_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17333_ top0.matmul0.matmul_stage_inst.mult2\[12\] _09318_ _09322_ VGND VGND VPWR
+ VPWR _09323_ sky130_fd_sc_hd__o21ai_2
X_14545_ _06729_ _06732_ _06750_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__o21a_2
XFILLER_0_173_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17264_ top0.matmul0.matmul_stage_inst.mult2\[2\] _09257_ _09258_ top0.matmul0.matmul_stage_inst.mult1\[2\]
+ VGND VGND VPWR VPWR _09264_ sky130_fd_sc_hd__a31o_1
X_14476_ _06554_ _06677_ _06603_ _06607_ _06672_ VGND VGND VPWR VPWR _06683_ sky130_fd_sc_hd__o221a_1
X_19003_ _10854_ _10855_ _10850_ VGND VGND VPWR VPWR _10977_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_141_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16215_ _08180_ _08306_ _08220_ VGND VGND VPWR VPWR _08307_ sky130_fd_sc_hd__o21ai_1
X_13427_ _05639_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17195_ _09203_ _09204_ VGND VGND VPWR VPWR _09205_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16146_ top0.pid_q.curr_int\[5\] _08083_ _08238_ VGND VGND VPWR VPWR _08239_ sky130_fd_sc_hd__o21ai_2
X_13358_ net43 _05489_ _05491_ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16077_ net473 net500 VGND VGND VPWR VPWR _08170_ sky130_fd_sc_hd__nand2_2
X_13289_ _05500_ _05501_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__nor2_1
X_19905_ _11771_ _11772_ _11778_ VGND VGND VPWR VPWR _11779_ sky130_fd_sc_hd__a21oi_1
X_15028_ _07142_ VGND VGND VPWR VPWR _07143_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_126_Left_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19836_ _11654_ _11560_ VGND VGND VPWR VPWR _11714_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19767_ _11649_ VGND VGND VPWR VPWR _11650_ sky130_fd_sc_hd__buf_4
X_16979_ top0.currT_r\[11\] _09034_ VGND VGND VPWR VPWR _09035_ sky130_fd_sc_hd__xnor2_1
Xinput3 spi_mosi VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
X_18718_ net381 net312 VGND VGND VPWR VPWR _10695_ sky130_fd_sc_hd__nand2_1
X_19698_ _11581_ _11583_ VGND VGND VPWR VPWR _11584_ sky130_fd_sc_hd__xor2_4
XFILLER_0_189_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18649_ _10621_ _10624_ VGND VGND VPWR VPWR _10627_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21660_ net81 net96 VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_135_Left_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20611_ _12427_ _12458_ _12459_ VGND VGND VPWR VPWR _12460_ sky130_fd_sc_hd__nand3_2
XFILLER_0_15_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21591_ _01150_ _01152_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20542_ _12360_ _12390_ _12372_ VGND VGND VPWR VPWR _12391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23330_ _02755_ _02764_ net133 VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20473_ _12316_ _12321_ VGND VGND VPWR VPWR _12322_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23261_ net291 net286 net278 net272 net198 net192 VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__mux4_1
XFILLER_0_85_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25000_ _03474_ _03719_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22212_ _01765_ _01772_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__xnor2_2
X_23192_ _05719_ _06945_ _02648_ net774 VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22143_ net133 _01076_ _01208_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_144_Left_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26951_ clknet_leaf_9_clk_sys _00568_ net596 VGND VGND VPWR VPWR top0.matmul0.a\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_22074_ _01632_ _01635_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_168_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25902_ _08900_ _05110_ _05115_ _05118_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__o31a_1
X_21025_ _12869_ _12795_ _11759_ VGND VGND VPWR VPWR _12872_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26882_ clknet_leaf_41_clk_sys _00499_ net683 VGND VGND VPWR VPWR top0.svm0.tB\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25833_ top0.c_out_calc\[4\] _05029_ _05031_ _05056_ VGND VGND VPWR VPWR _00735_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25764_ top0.matmul0.matmul_stage_inst.a\[10\] _04899_ _05457_ VGND VGND VPWR VPWR
+ _05003_ sky130_fd_sc_hd__mux2_1
X_22976_ top0.svm0.delta\[7\] VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24715_ _03908_ _04067_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__or2_1
XFILLER_0_201_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21927_ top0.cordic0.vec\[1\]\[6\] _01487_ _01488_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_153_Left_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25695_ _04961_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24646_ _03996_ _03999_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21858_ net145 net129 VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20809_ net254 _12559_ _12657_ net285 VGND VGND VPWR VPWR _12658_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24577_ _03775_ _03776_ _03779_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_194_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21789_ _01337_ _01340_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14330_ _06461_ _06538_ _06539_ VGND VGND VPWR VPWR _06540_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26316_ spi0.data_packed\[56\] spi0.data_packed\[57\] net698 VGND VGND VPWR VPWR
+ _05390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23528_ top0.a_in_matmul\[4\] top0.matmul0.a\[4\] _02926_ VGND VGND VPWR VPWR _02930_
+ sky130_fd_sc_hd__mux2_1
X_27296_ clknet_3_0__leaf_clk_mosi _00910_ VGND VGND VPWR VPWR spi0.opcode\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14261_ _06470_ _06471_ VGND VGND VPWR VPWR _06472_ sky130_fd_sc_hd__nor2_2
X_26247_ _05355_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23459_ net85 _11649_ _02892_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__and3_1
X_16000_ net448 net526 VGND VGND VPWR VPWR _08094_ sky130_fd_sc_hd__nand2_1
X_13212_ _05437_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14192_ net48 _05723_ _05724_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__and3_1
X_26178_ net19 _05314_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_162_Left_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25129_ net1017 _04272_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17951_ net416 net319 VGND VGND VPWR VPWR _09937_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16902_ top0.pid_q.curr_error\[5\] _08951_ VGND VGND VPWR VPWR _08963_ sky130_fd_sc_hd__or2_1
X_17882_ _09757_ _09867_ _09868_ VGND VGND VPWR VPWR _09869_ sky130_fd_sc_hd__a21oi_2
X_19621_ _11484_ _11504_ _11509_ VGND VGND VPWR VPWR _11510_ sky130_fd_sc_hd__a21oi_4
X_16833_ net492 _08890_ _08898_ _07710_ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19552_ net121 net1031 net113 net108 net198 net191 VGND VGND VPWR VPWR _11441_ sky130_fd_sc_hd__mux4_1
X_16764_ top0.pid_q.out\[15\] _08843_ _08847_ VGND VGND VPWR VPWR _08848_ sky130_fd_sc_hd__mux2_1
X_13976_ _06187_ _06141_ _06188_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_171_Left_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18503_ _10365_ _10367_ _10482_ VGND VGND VPWR VPWR _10483_ sky130_fd_sc_hd__a21oi_2
X_15715_ _07786_ _07789_ _07811_ VGND VGND VPWR VPWR _07812_ sky130_fd_sc_hd__a21oi_1
X_16695_ _08777_ _08779_ VGND VGND VPWR VPWR _08780_ sky130_fd_sc_hd__nand2_1
X_19483_ top0.pid_d.curr_int\[11\] top0.pid_d.prev_int\[11\] VGND VGND VPWR VPWR _11377_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18434_ _10411_ _10414_ VGND VGND VPWR VPWR _10415_ sky130_fd_sc_hd__or2_1
X_15646_ _07650_ _07651_ _07652_ VGND VGND VPWR VPWR _07744_ sky130_fd_sc_hd__o21a_1
XFILLER_0_186_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_186_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18365_ _10306_ _10316_ _10345_ VGND VGND VPWR VPWR _10346_ sky130_fd_sc_hd__o21a_1
XFILLER_0_185_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15577_ _07671_ _07675_ VGND VGND VPWR VPWR _07676_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17316_ net430 _09308_ net562 VGND VGND VPWR VPWR _09309_ sky130_fd_sc_hd__mux2_1
X_14528_ _06729_ _06734_ VGND VGND VPWR VPWR _06735_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18296_ net329 net382 VGND VGND VPWR VPWR _10278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17247_ _09094_ _09135_ _09192_ _08842_ _09250_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__a221o_1
X_14459_ _06596_ _06664_ _06662_ _06560_ VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_180_Left_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17178_ net543 _08320_ _09189_ net554 _08981_ VGND VGND VPWR VPWR _09190_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16129_ _08132_ _08133_ _08221_ VGND VGND VPWR VPWR _08222_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19819_ net1013 _11697_ _11689_ VGND VGND VPWR VPWR _11699_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22830_ _02345_ top0.svm0.tA\[11\] VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22761_ top0.pid_q.prev_int\[5\] _02292_ _02295_ top0.pid_q.curr_int\[5\] VGND VGND
+ VPWR VPWR _00424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24500_ top0.matmul0.matmul_stage_inst.mult2\[2\] _03855_ _03642_ VGND VGND VPWR
+ VPWR _03856_ sky130_fd_sc_hd__mux2_1
X_21712_ net149 _01149_ _01273_ net164 net158 VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__o221a_1
X_25480_ _04762_ _04664_ _04821_ _04755_ _04822_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__a32o_1
XFILLER_0_52_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22692_ net97 net87 net91 net79 VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__a211o_1
XFILLER_0_192_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24431_ _03709_ _03710_ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21643_ _01108_ _01198_ _01202_ net160 _01204_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__a221o_4
XFILLER_0_164_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27150_ clknet_leaf_12_clk_sys _00764_ net618 VGND VGND VPWR VPWR top0.b_in_matmul\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_24362_ _03717_ _03718_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__nor2_2
X_21574_ net154 net149 VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__and2_2
XANTENNA_30 net1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_41 top0.matmul0.matmul_stage_inst.e\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_26101_ top0.periodTop\[0\] _05276_ _05278_ net68 VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23313_ net150 _02719_ _02758_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__o21a_1
X_27081_ clknet_leaf_0_clk_sys _00698_ net586 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_20525_ _12069_ _12060_ VGND VGND VPWR VPWR _12374_ sky130_fd_sc_hd__xor2_1
X_24293_ _03299_ _03300_ _03631_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__or3_1
XFILLER_0_104_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26032_ top0.pid_d.out\[1\] _05198_ _05199_ spi0.data_packed\[65\] VGND VGND VPWR
+ VPWR _05225_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20456_ _12284_ _12285_ VGND VGND VPWR VPWR _12305_ sky130_fd_sc_hd__nor2_1
X_23244_ _11484_ _11504_ _11509_ _02693_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__a211o_1
XFILLER_0_162_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23175_ _05717_ _07028_ _02644_ net777 VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__a22o_1
X_20387_ _12137_ _12234_ _12235_ VGND VGND VPWR VPWR _12236_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_75_clk_sys clknet_3_4__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_75_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_22126_ _01063_ _01225_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26934_ clknet_leaf_7_clk_sys _00551_ net593 VGND VGND VPWR VPWR top0.matmul0.cos\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_22057_ _01614_ _01618_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__xnor2_4
X_21008_ _12697_ _12853_ _11739_ VGND VGND VPWR VPWR _12855_ sky130_fd_sc_hd__o21a_1
XFILLER_0_199_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26865_ clknet_leaf_41_clk_sys _00482_ net683 VGND VGND VPWR VPWR top0.svm0.tA\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25816_ net798 _05029_ _05031_ _05041_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__a22o_1
X_13830_ _06002_ _06042_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__xnor2_1
X_26796_ clknet_leaf_104_clk_sys _00413_ net576 VGND VGND VPWR VPWR top0.cordic0.gm0.iter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap10 net1012 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
XFILLER_0_98_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13761_ net54 _05489_ _05491_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__and3_1
X_25747_ net768 _04925_ _04994_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22959_ _02440_ _02469_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15500_ net480 _07258_ _07259_ _07598_ VGND VGND VPWR VPWR _07599_ sky130_fd_sc_hd__o22a_2
X_16480_ _08500_ _08505_ _08495_ VGND VGND VPWR VPWR _08568_ sky130_fd_sc_hd__o21ba_1
X_13692_ _05883_ _05903_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__nand2_1
X_25678_ net854 _04904_ _04936_ _04948_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15431_ _07251_ _07300_ VGND VGND VPWR VPWR _07530_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24629_ _03902_ _03903_ _03982_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__a21o_1
X_18150_ _10001_ _10005_ _10003_ VGND VGND VPWR VPWR _10134_ sky130_fd_sc_hd__o21a_1
X_15362_ net533 _07446_ VGND VGND VPWR VPWR _07461_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17101_ top0.pid_q.curr_error\[9\] _08860_ _09117_ VGND VGND VPWR VPWR _09127_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14313_ _06437_ _06438_ _06522_ VGND VGND VPWR VPWR _06523_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18081_ net434 _09985_ _10065_ net439 _07138_ VGND VGND VPWR VPWR _10066_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15293_ _07390_ _07391_ VGND VGND VPWR VPWR _07392_ sky130_fd_sc_hd__nand2_1
X_27279_ clknet_3_4__leaf_clk_mosi _00893_ VGND VGND VPWR VPWR spi0.data_packed\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17032_ _09079_ _09080_ _09082_ _09083_ _09059_ VGND VGND VPWR VPWR _09084_ sky130_fd_sc_hd__a41o_1
X_14244_ _06282_ _06283_ _06454_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14175_ _06256_ _06370_ _06371_ _06385_ VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18983_ net363 _10877_ _10956_ VGND VGND VPWR VPWR _10957_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17934_ net346 net380 VGND VGND VPWR VPWR _09920_ sky130_fd_sc_hd__nand2_1
XFILLER_0_178_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17865_ net404 net336 net399 net339 VGND VGND VPWR VPWR _09852_ sky130_fd_sc_hd__nand4_1
X_19604_ top0.cordic0.slte0.opB\[9\] _11492_ VGND VGND VPWR VPWR _11493_ sky130_fd_sc_hd__or2_1
X_16816_ top0.matmul0.beta_pass\[0\] _05438_ VGND VGND VPWR VPWR _08883_ sky130_fd_sc_hd__nand2_1
X_17796_ net413 net329 VGND VGND VPWR VPWR _09783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19535_ _11422_ VGND VGND VPWR VPWR _11425_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_187_Right_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13959_ _05786_ _05787_ _05796_ _05794_ _05789_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__o32a_1
X_16747_ _08808_ _08830_ VGND VGND VPWR VPWR _08831_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16678_ _08701_ _08702_ _08703_ VGND VGND VPWR VPWR _08763_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19466_ _11359_ _11360_ VGND VGND VPWR VPWR _11362_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_185_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18417_ _10394_ _10397_ VGND VGND VPWR VPWR _10398_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15629_ net506 net488 VGND VGND VPWR VPWR _07727_ sky130_fd_sc_hd__nand2_1
X_19397_ top0.pid_d.curr_int\[1\] top0.pid_d.prev_int\[1\] VGND VGND VPWR VPWR _11301_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18348_ _10326_ _10329_ VGND VGND VPWR VPWR _10330_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18279_ net406 net312 VGND VGND VPWR VPWR _10261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20310_ _12155_ _12158_ VGND VGND VPWR VPWR _12159_ sky130_fd_sc_hd__nor2_1
X_21290_ _13127_ _13132_ VGND VGND VPWR VPWR _13133_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20241_ net270 net264 VGND VGND VPWR VPWR _12090_ sky130_fd_sc_hd__nor2_1
X_20172_ _12015_ _12023_ VGND VGND VPWR VPWR _12024_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24980_ _04322_ _04324_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23931_ _03130_ _03288_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__xor2_2
X_26650_ clknet_leaf_76_clk_sys _00267_ net639 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_23862_ _03214_ _03215_ _03218_ _03219_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25601_ _04886_ top0.matmul0.cos\[4\] _04878_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__or3_1
X_22813_ _02331_ top0.svm0.tA\[5\] top0.svm0.tA\[4\] _02332_ VGND VGND VPWR VPWR _02333_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26581_ clknet_leaf_53_clk_sys _00204_ net674 VGND VGND VPWR VPWR top0.pid_q.prev_error\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_23793_ net572 top0.matmul0.matmul_stage_inst.d\[12\] top0.matmul0.matmul_stage_inst.c\[12\]
+ net556 VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__a22o_2
XFILLER_0_196_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25532_ _04852_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__clkbuf_1
X_22744_ _11654_ _02287_ VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_177_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25463_ _04802_ _04803_ _04804_ _04805_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__or4b_2
XFILLER_0_177_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22675_ _02180_ _02225_ _02226_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_176_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27202_ clknet_leaf_92_clk_sys _00816_ net599 VGND VGND VPWR VPWR top0.cordic0.slte0.opB\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_24414_ _03045_ _03046_ _03150_ _03151_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__o22a_1
XFILLER_0_164_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21626_ net149 _01186_ _01187_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__a21oi_1
X_25394_ _04733_ _04737_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27133_ clknet_leaf_11_clk_sys _00747_ net601 VGND VGND VPWR VPWR top0.matmul0.op_in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24345_ _03206_ _03223_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__and2_1
X_21557_ net115 net110 VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20508_ _12341_ _12343_ _12356_ VGND VGND VPWR VPWR _12357_ sky130_fd_sc_hd__a21oi_2
X_27064_ clknet_leaf_110_clk_sys _00681_ net578 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.c\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_24276_ _03450_ _03618_ _03627_ _03633_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_50_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21488_ _01023_ _01037_ _01038_ _01049_ _01022_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_200_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26015_ _05212_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__clkbuf_1
X_23227_ net161 _02669_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__nand2_1
X_20439_ _11571_ _12287_ _12108_ net296 VGND VGND VPWR VPWR _12288_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23158_ top0.svm0.state\[1\] VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22109_ _01637_ _01605_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__nand2_1
X_15980_ _07998_ _08074_ VGND VGND VPWR VPWR _08075_ sky130_fd_sc_hd__xor2_1
X_23089_ net40 net169 VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14931_ spi0.data_packed\[40\] top0.kid\[8\] _07086_ VGND VGND VPWR VPWR _07087_
+ sky130_fd_sc_hd__mux2_1
X_26917_ clknet_leaf_3_clk_sys _00534_ net583 VGND VGND VPWR VPWR top0.matmul0.sin\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_17650_ net382 net355 VGND VGND VPWR VPWR _09637_ sky130_fd_sc_hd__nand2_1
X_14862_ _07050_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__clkbuf_1
X_26848_ clknet_leaf_44_clk_sys _00465_ net686 VGND VGND VPWR VPWR top0.svm0.delta\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_202_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13813_ net68 _06025_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__nand2_1
X_16601_ _08491_ _08548_ _08547_ VGND VGND VPWR VPWR _08687_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17581_ net415 net418 net423 net358 VGND VGND VPWR VPWR _09568_ sky130_fd_sc_hd__and4b_1
X_14793_ _06949_ _06993_ _06990_ VGND VGND VPWR VPWR _06994_ sky130_fd_sc_hd__o21a_1
X_26779_ clknet_leaf_6_clk_sys _00396_ net590 VGND VGND VPWR VPWR top0.cordic0.cos\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19320_ _11258_ _11254_ _11255_ VGND VGND VPWR VPWR _11260_ sky130_fd_sc_hd__or3_1
X_16532_ top0.pid_q.out\[12\] top0.pid_q.curr_int\[12\] VGND VGND VPWR VPWR _08619_
+ sky130_fd_sc_hd__nand2_1
X_13744_ _05947_ _05926_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19251_ top0.pid_d.prev_error\[8\] top0.pid_d.curr_error\[8\] VGND VGND VPWR VPWR
+ _11197_ sky130_fd_sc_hd__xnor2_1
X_16463_ top0.pid_q.out\[10\] _08551_ net13 VGND VGND VPWR VPWR _08552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13675_ _05839_ _05840_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__xor2_1
XFILLER_0_156_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18202_ _10105_ _10110_ _10184_ VGND VGND VPWR VPWR _10185_ sky130_fd_sc_hd__a21o_1
X_15414_ _07511_ _07512_ _07501_ VGND VGND VPWR VPWR _07513_ sky130_fd_sc_hd__a21o_1
X_19182_ top0.pid_d.prev_error\[0\] top0.pid_d.curr_error\[0\] top0.pid_d.prev_error\[1\]
+ top0.pid_d.curr_error\[1\] VGND VGND VPWR VPWR _11134_ sky130_fd_sc_hd__a22o_1
X_16394_ top0.pid_q.out\[10\] top0.pid_q.curr_int\[10\] VGND VGND VPWR VPWR _08483_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_38_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18133_ net346 net372 VGND VGND VPWR VPWR _10117_ sky130_fd_sc_hd__nand2_1
X_15345_ _07436_ _07437_ VGND VGND VPWR VPWR _07444_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18064_ _10042_ _10048_ VGND VGND VPWR VPWR _10049_ sky130_fd_sc_hd__xnor2_1
X_15276_ _07365_ _07370_ VGND VGND VPWR VPWR _07375_ sky130_fd_sc_hd__nor2_1
Xhold108 top0.matmul0.matmul_stage_inst.b\[10\] VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__dlygate4sd3_1
X_17015_ _05662_ net428 top0.currT_r\[13\] _08899_ VGND VGND VPWR VPWR _09068_ sky130_fd_sc_hd__or4_1
XFILLER_0_110_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14227_ net22 _05523_ _05524_ VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__and3_2
Xhold119 top0.matmul0.matmul_stage_inst.b\[3\] VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14158_ _06358_ _06369_ VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__xor2_4
XFILLER_0_81_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14089_ _06296_ _06297_ _06298_ _06299_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__o22a_1
X_18966_ _09965_ _10384_ net311 net373 VGND VGND VPWR VPWR _10940_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17917_ net339 net388 VGND VGND VPWR VPWR _09903_ sky130_fd_sc_hd__nand2_2
X_18897_ _10869_ _10871_ VGND VGND VPWR VPWR _10872_ sky130_fd_sc_hd__xor2_1
X_17848_ net336 net399 VGND VGND VPWR VPWR _09835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17779_ _09764_ _09765_ VGND VGND VPWR VPWR _09766_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19518_ _11407_ VGND VGND VPWR VPWR _11408_ sky130_fd_sc_hd__buf_4
XFILLER_0_53_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_23_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_23_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20790_ _11653_ _12273_ VGND VGND VPWR VPWR _12639_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19449_ _11345_ _11346_ VGND VGND VPWR VPWR _11347_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22460_ net109 _02014_ _02016_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_134_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21411_ net218 _12765_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22391_ _01948_ _01934_ _01938_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__or3_1
XFILLER_0_173_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24130_ _03485_ _03487_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21342_ _13161_ _13183_ VGND VGND VPWR VPWR _13184_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_142_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24061_ _03402_ _03384_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__and2b_1
X_21273_ _12207_ _13031_ _13113_ net247 _13115_ VGND VGND VPWR VPWR _13116_ sky130_fd_sc_hd__a221o_1
Xclkbuf_3_5__f_clk_sys clknet_0_clk_sys VGND VGND VPWR VPWR clknet_3_5__leaf_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23012_ _02514_ _02510_ _02515_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20224_ net247 net234 VGND VGND VPWR VPWR _12073_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20155_ _12007_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24963_ _04305_ _04313_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__xnor2_1
X_20086_ top0.cordic0.slte0.opA\[11\] _11945_ _11946_ _11944_ VGND VGND VPWR VPWR
+ _00371_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23914_ _03256_ _03259_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__nand2_1
X_26702_ clknet_leaf_82_clk_sys net890 net646 VGND VGND VPWR VPWR top0.pid_d.prev_error\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_24894_ _04166_ _04241_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26633_ clknet_leaf_82_clk_sys _00250_ net638 VGND VGND VPWR VPWR top0.pid_d.out\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_23845_ _03076_ _03077_ _03090_ _03091_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__o22a_1
XFILLER_0_197_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26564_ clknet_leaf_53_clk_sys _00187_ net671 VGND VGND VPWR VPWR top0.pid_q.curr_error\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23776_ _03075_ _03082_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__xnor2_4
X_20988_ _12818_ _12825_ _12831_ net213 _12834_ VGND VGND VPWR VPWR _12835_ sky130_fd_sc_hd__a221o_2
XFILLER_0_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25515_ _04843_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22727_ _02272_ _02276_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26495_ clknet_leaf_71_clk_sys _00118_ net657 VGND VGND VPWR VPWR top0.pid_d.prev_int\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_149_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13460_ _05669_ _05672_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__xnor2_1
X_25446_ _04288_ _03936_ _04787_ _04788_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__and4_1
XFILLER_0_193_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22658_ _02184_ _02210_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21609_ _01160_ _01170_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__xnor2_1
X_25377_ _04691_ _04690_ _04720_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__a21o_1
X_13391_ _05602_ _05603_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22589_ _02142_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__inv_2
X_15130_ net517 net493 _07228_ VGND VGND VPWR VPWR _07229_ sky130_fd_sc_hd__a21o_1
X_27116_ clknet_leaf_90_clk_sys _00730_ net600 VGND VGND VPWR VPWR top0.cordic_done
+ sky130_fd_sc_hd__dfrtp_1
X_24328_ _03177_ _03179_ _03178_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27047_ clknet_leaf_8_clk_sys _00664_ net592 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_15061_ _07154_ _07159_ VGND VGND VPWR VPWR _07160_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24259_ _03454_ _03616_ _03423_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_160_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14012_ _06223_ _06224_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__xor2_1
X_18820_ _10712_ _10795_ net320 VGND VGND VPWR VPWR _10796_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18751_ _10727_ VGND VGND VPWR VPWR _10728_ sky130_fd_sc_hd__inv_2
X_15963_ _08055_ _08057_ VGND VGND VPWR VPWR _08058_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17702_ _09688_ net381 VGND VGND VPWR VPWR _09689_ sky130_fd_sc_hd__nor2_1
X_14914_ spi0.data_packed\[32\] top0.kid\[0\] _07075_ VGND VGND VPWR VPWR _07078_
+ sky130_fd_sc_hd__mux2_1
X_18682_ _10494_ _10659_ VGND VGND VPWR VPWR _10660_ sky130_fd_sc_hd__xnor2_1
X_15894_ _07987_ _07989_ VGND VGND VPWR VPWR _07990_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17633_ net392 net349 VGND VGND VPWR VPWR _09620_ sky130_fd_sc_hd__nand2_1
X_14845_ state\[0\] net17 VGND VGND VPWR VPWR _07041_ sky130_fd_sc_hd__nand2_4
XFILLER_0_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14776_ _06975_ _06976_ VGND VGND VPWR VPWR _06977_ sky130_fd_sc_hd__xor2_2
X_17564_ _09549_ _09550_ net347 _09524_ VGND VGND VPWR VPWR _09551_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_147_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19303_ net315 _11117_ _11244_ _10067_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13727_ _05938_ _05939_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__xor2_1
X_16515_ _08316_ _08330_ _08393_ _08394_ VGND VGND VPWR VPWR _08603_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17495_ net413 net337 VGND VGND VPWR VPWR _09482_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19234_ _11121_ _11180_ _11181_ _11123_ VGND VGND VPWR VPWR _11182_ sky130_fd_sc_hd__a31o_1
X_13658_ _05869_ _05870_ net57 _05472_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__o211a_1
X_16446_ _08446_ _08534_ _08451_ VGND VGND VPWR VPWR _08535_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16377_ _08413_ _08466_ VGND VGND VPWR VPWR _08467_ sky130_fd_sc_hd__xnor2_2
X_19165_ top0.matmul0.done_pass top0.matmul0.state\[1\] top0.pid_d.state\[3\] VGND
+ VGND VPWR VPWR _11119_ sky130_fd_sc_hd__and3_1
X_13589_ _05559_ _05598_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__xor2_1
XFILLER_0_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18116_ net334 net383 VGND VGND VPWR VPWR _10100_ sky130_fd_sc_hd__nand2_1
X_15328_ _07374_ _07405_ _07406_ _07424_ _07426_ VGND VGND VPWR VPWR _07427_ sky130_fd_sc_hd__o32a_1
XFILLER_0_170_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19096_ _11062_ _11067_ VGND VGND VPWR VPWR _11068_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18047_ _09903_ _09904_ _09905_ VGND VGND VPWR VPWR _10032_ sky130_fd_sc_hd__o21a_1
X_15259_ _07356_ _07357_ VGND VGND VPWR VPWR _07358_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout407 net408 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout418 net420 VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__buf_2
Xfanout429 net430 VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__clkbuf_4
X_19998_ _11860_ _11864_ top0.cordic0.gm0.iter\[4\] VGND VGND VPWR VPWR _11865_ sky130_fd_sc_hd__a21oi_2
X_18949_ _10829_ _10841_ VGND VGND VPWR VPWR _10923_ sky130_fd_sc_hd__or2b_1
XFILLER_0_193_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21960_ _01325_ _01515_ _01517_ net137 VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_146_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20911_ net265 _12715_ _12757_ _12758_ VGND VGND VPWR VPWR _12759_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21891_ _01444_ _01435_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23630_ net574 top0.matmul0.matmul_stage_inst.d\[7\] top0.matmul0.matmul_stage_inst.c\[7\]
+ net558 VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__a22o_1
X_20842_ _11593_ _12040_ VGND VGND VPWR VPWR _12691_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23561_ top0.b_in_matmul\[4\] top0.matmul0.b\[4\] _02937_ VGND VGND VPWR VPWR _02947_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout14 net55 VGND VGND VPWR VPWR net1025 sky130_fd_sc_hd__buf_4
X_20773_ _12614_ _12621_ VGND VGND VPWR VPWR _12622_ sky130_fd_sc_hd__xor2_2
XFILLER_0_18_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout25 net27 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25300_ _04069_ _04339_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__nand2_1
Xfanout36 net37 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_4
Xfanout47 top0.periodTop_r\[7\] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_4
X_22512_ _02064_ _02067_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__xor2_2
Xfanout58 top0.periodTop_r\[3\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_4
X_26280_ net953 spi0.data_packed\[39\] net688 VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23492_ top0.cordic0.cos\[1\] top0.matmul0.cos\[1\] _02904_ VGND VGND VPWR VPWR _02911_
+ sky130_fd_sc_hd__mux2_1
Xfanout69 top0.matmul0.op\[1\] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_2
XFILLER_0_135_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25231_ _04508_ _04577_ _04506_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_29_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22443_ _01943_ _01942_ _01987_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25162_ _04069_ _04509_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_17_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22374_ _01931_ _01932_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__and2b_1
X_24113_ _03468_ _03470_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__nand2_2
XFILLER_0_115_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21325_ _13163_ _13166_ net235 VGND VGND VPWR VPWR _13167_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25093_ _04355_ _04357_ _04356_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24044_ _03342_ _03344_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_13_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21256_ _12939_ _12950_ _12938_ VGND VGND VPWR VPWR _13100_ sky130_fd_sc_hd__a21o_1
XFILLER_0_187_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20207_ net269 _12049_ VGND VGND VPWR VPWR _12056_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21187_ net257 net234 VGND VGND VPWR VPWR _13031_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_198_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20138_ _11967_ _11968_ VGND VGND VPWR VPWR _11994_ sky130_fd_sc_hd__or2_1
X_25995_ top0.b_in_matmul\[8\] _05195_ _05196_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__mux2_1
X_24946_ _04199_ _04200_ _04296_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__o21a_1
X_20069_ _11924_ _11925_ _11930_ VGND VGND VPWR VPWR _11931_ sky130_fd_sc_hd__o21a_1
XFILLER_0_197_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24877_ _04114_ _04115_ _04227_ _04228_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__or4_1
X_14630_ net20 _05640_ _05629_ _06106_ VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__a211o_1
XFILLER_0_158_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26616_ clknet_leaf_29_clk_sys _00233_ net623 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_23828_ _03185_ _03152_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__nor2_2
XFILLER_0_200_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14561_ net41 _06131_ VGND VGND VPWR VPWR _06767_ sky130_fd_sc_hd__nand2_1
X_26547_ clknet_leaf_49_clk_sys _00170_ net675 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_166_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23759_ _03004_ _03005_ _03054_ _03055_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__o22a_1
XFILLER_0_95_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13512_ net60 _05723_ _05724_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__and3_1
XFILLER_0_166_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16300_ _08254_ _08311_ _08313_ VGND VGND VPWR VPWR _08391_ sky130_fd_sc_hd__a21o_1
X_17280_ _09276_ _09277_ VGND VGND VPWR VPWR _09278_ sky130_fd_sc_hd__xnor2_1
X_14492_ _06636_ _06650_ _06698_ VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_138_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26478_ clknet_leaf_11_clk_sys _00109_ net604 VGND VGND VPWR VPWR top0.periodTop\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16231_ _07800_ _08322_ VGND VGND VPWR VPWR _08323_ sky130_fd_sc_hd__and2_1
X_25429_ _04516_ _04771_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__nand2_1
X_13443_ net56 _05602_ _05603_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16162_ _08219_ _08223_ _08253_ VGND VGND VPWR VPWR _08254_ sky130_fd_sc_hd__o21ai_2
X_13374_ _05543_ _05545_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__nor2_2
XFILLER_0_24_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15113_ _07149_ _07159_ VGND VGND VPWR VPWR _07212_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16093_ top0.pid_q.mult0.b\[13\] net523 VGND VGND VPWR VPWR _08186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_39_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15044_ net941 _07139_ _07143_ top0.pid_d.curr_int\[14\] VGND VGND VPWR VPWR _00131_
+ sky130_fd_sc_hd__a22o_1
X_19921_ _11650_ _11793_ net1020 VGND VGND VPWR VPWR _11794_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19852_ _11514_ _11728_ VGND VGND VPWR VPWR _11729_ sky130_fd_sc_hd__and2_1
X_18803_ net374 _09395_ _09356_ VGND VGND VPWR VPWR _10779_ sky130_fd_sc_hd__a21oi_1
X_19783_ net272 _11644_ VGND VGND VPWR VPWR _11665_ sky130_fd_sc_hd__or2_1
X_16995_ _09046_ _09049_ VGND VGND VPWR VPWR _09050_ sky130_fd_sc_hd__xnor2_1
X_18734_ net320 net373 VGND VGND VPWR VPWR _10711_ sky130_fd_sc_hd__nand2_1
X_15946_ net468 net509 VGND VGND VPWR VPWR _08041_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18665_ net334 net338 net369 net331 VGND VGND VPWR VPWR _10643_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_48_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15877_ _07970_ _07972_ VGND VGND VPWR VPWR _07973_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17616_ _09535_ _09547_ _09602_ VGND VGND VPWR VPWR _09603_ sky130_fd_sc_hd__o21ai_1
X_14828_ _07008_ _07027_ VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_188_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18596_ _10490_ _10502_ _10574_ VGND VGND VPWR VPWR _10575_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17547_ net403 net358 _09529_ _09533_ net354 VGND VGND VPWR VPWR _09534_ sky130_fd_sc_hd__a32o_1
X_14759_ _06921_ _06922_ VGND VGND VPWR VPWR _06961_ sky130_fd_sc_hd__nand2_1
XFILLER_0_175_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17478_ net354 _09464_ VGND VGND VPWR VPWR _09465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19217_ _11164_ _11156_ _11165_ VGND VGND VPWR VPWR _11166_ sky130_fd_sc_hd__a21o_1
X_16429_ _08515_ _08517_ VGND VGND VPWR VPWR _08518_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19148_ net393 _11096_ _11109_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19079_ _10690_ net370 _10495_ _10790_ VGND VGND VPWR VPWR _11051_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21110_ _12805_ _12880_ _12878_ VGND VGND VPWR VPWR _12956_ sky130_fd_sc_hd__or3b_1
X_22090_ _01650_ _01651_ _01614_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21041_ _12878_ _12887_ VGND VGND VPWR VPWR _12888_ sky130_fd_sc_hd__xor2_2
XFILLER_0_160_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout204 top0.cordic0.gm0.iter\[0\] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_4
Xfanout215 net217 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_4
Xfanout226 top0.cordic0.vec\[0\]\[15\] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__buf_2
XFILLER_0_201_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout237 top0.cordic0.vec\[0\]\[13\] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_4
Xfanout248 top0.cordic0.vec\[0\]\[11\] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__buf_4
Xfanout259 net261 VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_4
X_24800_ _04066_ _04152_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__xor2_1
X_25780_ _12030_ _12023_ _05011_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__o21ai_1
X_22992_ _02497_ _02493_ _02498_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_158_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24731_ _04003_ _04004_ _04082_ _04083_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__or4_1
X_21943_ _01320_ net154 VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24662_ _04014_ _04015_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__xor2_1
X_21874_ net151 _01122_ _01338_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__a21o_1
X_26401_ clknet_leaf_98_clk_sys _00042_ net588 VGND VGND VPWR VPWR top0.kpd\[6\] sky130_fd_sc_hd__dfrtp_1
X_23613_ _02973_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20825_ _12420_ _12668_ _12673_ VGND VGND VPWR VPWR _12674_ sky130_fd_sc_hd__a21o_1
XFILLER_0_194_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24593_ _03928_ _03947_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_148_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26332_ spi0.data_packed\[64\] spi0.data_packed\[65\] net693 VGND VGND VPWR VPWR
+ _05398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23544_ _02938_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__clkbuf_1
X_20756_ _11593_ net258 _12589_ _12600_ _12604_ VGND VGND VPWR VPWR _12605_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26263_ _05363_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23475_ net1000 top0.matmul0.sin\[7\] _05461_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20687_ _12487_ _12489_ _12533_ _12535_ VGND VGND VPWR VPWR _12536_ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25214_ _03325_ _03254_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__nand2_2
XFILLER_0_163_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22426_ _01978_ _01983_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26194_ _05327_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25145_ _03325_ _03254_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22357_ _01217_ _01913_ _01915_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_131_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21308_ _12036_ _13150_ VGND VGND VPWR VPWR _13151_ sky130_fd_sc_hd__nor2_1
X_25076_ _03474_ _04182_ _04348_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__o21ai_1
X_22288_ _01846_ _01847_ net81 VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__mux2_1
X_24027_ _03010_ _03157_ VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__nand2_1
Xhold280 top0.b_in_matmul\[11\] VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__dlygate4sd3_1
X_21239_ _12610_ _13082_ _12642_ VGND VGND VPWR VPWR _13083_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold291 top0.pid_q.prev_int\[0\] VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__dlygate4sd3_1
X_15800_ top0.pid_q.out\[2\] _07704_ _07806_ net544 _07896_ VGND VGND VPWR VPWR _07897_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_176_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13992_ net37 net1015 VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__nand2_2
X_16780_ net542 _08856_ _08859_ net843 _08862_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__a221o_1
X_25978_ top0.b_in_matmul\[4\] _05183_ _05165_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15731_ _07745_ _07747_ _07827_ VGND VGND VPWR VPWR _07828_ sky130_fd_sc_hd__o21ai_2
X_24929_ net1017 _03200_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18450_ top0.pid_d.out\[7\] top0.pid_d.curr_int\[7\] VGND VGND VPWR VPWR _10430_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15662_ _07750_ _07759_ VGND VGND VPWR VPWR _07760_ sky130_fd_sc_hd__xor2_1
X_17401_ net338 net423 VGND VGND VPWR VPWR _09388_ sky130_fd_sc_hd__nand2_1
X_14613_ _06751_ _06790_ _06749_ VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__o21a_1
XFILLER_0_200_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18381_ _10358_ _10360_ VGND VGND VPWR VPWR _10362_ sky130_fd_sc_hd__nand2_1
X_15593_ _07599_ _07606_ _07691_ _07596_ VGND VGND VPWR VPWR _07692_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14544_ _06729_ _06732_ _06733_ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__a21bo_1
X_17332_ top0.matmul0.matmul_stage_inst.mult2\[12\] _09318_ top0.matmul0.matmul_stage_inst.mult1\[12\]
+ VGND VGND VPWR VPWR _09322_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14475_ net864 _06280_ _06682_ _06381_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17263_ top0.matmul0.matmul_stage_inst.mult2\[2\] VGND VGND VPWR VPWR _09263_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19002_ _10935_ _10975_ VGND VGND VPWR VPWR _10976_ sky130_fd_sc_hd__xnor2_1
X_13426_ _05637_ _05638_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__nor2_4
X_16214_ _08174_ _08179_ VGND VGND VPWR VPWR _08306_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17194_ top0.pid_q.curr_int\[9\] top0.pid_q.prev_int\[9\] VGND VGND VPWR VPWR _09204_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16145_ top0.pid_q.curr_int\[5\] _08083_ top0.pid_q.out\[5\] VGND VGND VPWR VPWR
+ _08238_ sky130_fd_sc_hd__a21o_1
X_13357_ _05568_ _05569_ VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16076_ net468 net503 VGND VGND VPWR VPWR _08169_ sky130_fd_sc_hd__nand2_1
X_13288_ _05484_ _05486_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__nand2_1
X_19904_ _11773_ _11777_ VGND VGND VPWR VPWR _11778_ sky130_fd_sc_hd__xnor2_1
X_15027_ net437 net432 _05442_ _07141_ VGND VGND VPWR VPWR _07142_ sky130_fd_sc_hd__and4b_1
XFILLER_0_20_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19835_ _11706_ _11711_ _11712_ VGND VGND VPWR VPWR _11713_ sky130_fd_sc_hd__a21o_1
X_19766_ _11648_ VGND VGND VPWR VPWR _11649_ sky130_fd_sc_hd__clkbuf_4
X_16978_ top0.matmul0.beta_pass\[11\] _05438_ VGND VGND VPWR VPWR _09034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18717_ net317 _10692_ _10693_ _10208_ VGND VGND VPWR VPWR _10694_ sky130_fd_sc_hd__a22o_1
X_15929_ _08020_ _08023_ VGND VGND VPWR VPWR _08024_ sky130_fd_sc_hd__xnor2_2
X_19697_ _11511_ _11582_ VGND VGND VPWR VPWR _11583_ sky130_fd_sc_hd__nand2_2
XFILLER_0_190_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18648_ _10625_ VGND VGND VPWR VPWR _10626_ sky130_fd_sc_hd__inv_2
X_18579_ _10555_ _10557_ VGND VGND VPWR VPWR _10558_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_143_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20610_ _12457_ _12446_ _12455_ VGND VGND VPWR VPWR _12459_ sky130_fd_sc_hd__nand3_1
XFILLER_0_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21590_ _01136_ _01151_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20541_ _12271_ _12275_ VGND VGND VPWR VPWR _12390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23260_ net268 net259 net254 net251 net204 net196 VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__mux4_1
XFILLER_0_172_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20472_ _12319_ _12320_ VGND VGND VPWR VPWR _12321_ sky130_fd_sc_hd__or2b_1
XFILLER_0_43_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22211_ _01768_ _01771_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23191_ _02646_ _06907_ _02649_ net797 VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22142_ net133 _01208_ _01702_ _01703_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__and4_1
XFILLER_0_112_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26950_ clknet_leaf_13_clk_sys _00567_ net616 VGND VGND VPWR VPWR top0.matmul0.a\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_22073_ _01560_ _01633_ _01634_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_26_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25901_ _05110_ _05117_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__nand2_1
X_21024_ _12869_ _12783_ _12870_ net225 VGND VGND VPWR VPWR _12871_ sky130_fd_sc_hd__a211o_1
XFILLER_0_199_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26881_ clknet_leaf_41_clk_sys _00498_ net685 VGND VGND VPWR VPWR top0.svm0.tB\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25832_ _05052_ _05055_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22975_ net170 _02482_ _02484_ _02481_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__a22o_1
X_25763_ _05002_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24714_ _03315_ _03974_ VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__xnor2_2
X_21926_ net151 net129 VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__nand2_1
X_25694_ top0.matmul0.matmul_stage_inst.c\[14\] _04896_ _04960_ VGND VGND VPWR VPWR
+ _04961_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_85_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24645_ _03997_ _03998_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21857_ _01408_ _01409_ _01418_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_71_clk_sys clknet_3_5__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_71_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20808_ net254 _12559_ _12650_ _12652_ _12654_ VGND VGND VPWR VPWR _12657_ sky130_fd_sc_hd__o2111a_1
X_24576_ _03781_ _03929_ _03930_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__o21bai_2
X_21788_ _01342_ _01349_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__xor2_1
XFILLER_0_182_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26315_ _05389_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__clkbuf_1
X_23527_ _02929_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20739_ net294 net282 net264 VGND VGND VPWR VPWR _12588_ sky130_fd_sc_hd__and3_1
X_27295_ clknet_3_0__leaf_clk_mosi _00909_ VGND VGND VPWR VPWR spi0.opcode\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14260_ _06389_ _06390_ _06469_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__and3_1
XFILLER_0_151_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26246_ spi0.data_packed\[21\] spi0.data_packed\[22\] net698 VGND VGND VPWR VPWR
+ _05355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23458_ net85 _11857_ _02892_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__nor3_1
XFILLER_0_163_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13211_ _05436_ VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22409_ _01131_ _01759_ _01761_ _01762_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__a211o_2
X_14191_ net1025 _05721_ VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26177_ spi0.data_packed\[8\] _05310_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__and2_1
X_23389_ _02827_ _02829_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25128_ _02982_ _03936_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25059_ _04391_ _04407_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__or2_1
X_17950_ net355 net372 VGND VGND VPWR VPWR _09936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16901_ _08959_ _08961_ VGND VGND VPWR VPWR _08962_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_168_Right_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17881_ net378 net355 net375 net359 VGND VGND VPWR VPWR _09868_ sky130_fd_sc_hd__a22oi_1
X_19620_ _11483_ _11508_ top0.cordic0.slte0.opA\[17\] VGND VGND VPWR VPWR _11509_
+ sky130_fd_sc_hd__o21bai_4
X_16832_ net547 _08894_ _08897_ net550 _08881_ VGND VGND VPWR VPWR _08898_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout590 net598 VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__clkbuf_4
X_19551_ net103 net98 net94 net88 net199 top0.cordic0.gm0.iter\[1\] VGND VGND VPWR
+ VPWR _11440_ sky130_fd_sc_hd__mux4_2
X_16763_ top0.pid_q.curr_int\[15\] _08846_ VGND VGND VPWR VPWR _08847_ sky130_fd_sc_hd__xnor2_1
X_13975_ net48 _05639_ _06139_ _05625_ net1025 VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_38_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18502_ _10365_ _10367_ _10366_ VGND VGND VPWR VPWR _10482_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15714_ _07786_ _07789_ _07778_ VGND VGND VPWR VPWR _07811_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19482_ top0.pid_d.curr_int\[12\] top0.pid_d.prev_int\[12\] VGND VGND VPWR VPWR _11376_
+ sky130_fd_sc_hd__xor2_1
X_16694_ _08778_ VGND VGND VPWR VPWR _08779_ sky130_fd_sc_hd__inv_2
XFILLER_0_198_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18433_ _10308_ _10412_ _10413_ VGND VGND VPWR VPWR _10414_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_185_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15645_ _07739_ _07742_ VGND VGND VPWR VPWR _07743_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18364_ _10306_ _10316_ _10304_ VGND VGND VPWR VPWR _10345_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15576_ _07564_ _07661_ _07673_ _07674_ VGND VGND VPWR VPWR _07675_ sky130_fd_sc_hd__o211a_1
X_17315_ _09306_ _09307_ VGND VGND VPWR VPWR _09308_ sky130_fd_sc_hd__xnor2_1
X_14527_ _06732_ _06733_ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__xnor2_1
X_18295_ _10175_ _10177_ _10276_ VGND VGND VPWR VPWR _10277_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_44_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17246_ net554 _05443_ _09134_ _09248_ _09249_ VGND VGND VPWR VPWR _09250_ sky130_fd_sc_hd__a41o_1
X_14458_ _06663_ _06664_ _06665_ _06662_ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__o22a_1
XFILLER_0_189_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13409_ net60 _05611_ _05612_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__and3_2
X_14389_ _06596_ _06597_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17177_ _09187_ _09188_ VGND VGND VPWR VPWR _09189_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16128_ _08132_ _08133_ _08130_ VGND VGND VPWR VPWR _08221_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16059_ _08090_ _08152_ VGND VGND VPWR VPWR _08153_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_110_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19818_ _11430_ _11697_ VGND VGND VPWR VPWR _11698_ sky130_fd_sc_hd__or2_1
XFILLER_0_194_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19749_ _11409_ VGND VGND VPWR VPWR _11632_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_194_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22760_ net982 _02292_ _02295_ top0.pid_q.curr_int\[4\] VGND VGND VPWR VPWR _00423_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21711_ _01091_ _01102_ net154 VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22691_ net100 _01924_ _01821_ _01762_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24430_ _03709_ _03710_ _03711_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21642_ _01200_ _01203_ net138 _01199_ VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24361_ net566 net560 top0.matmul0.matmul_stage_inst.e\[14\] VGND VGND VPWR VPWR
+ _03718_ sky130_fd_sc_hd__o21a_2
XFILLER_0_74_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_20 net1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21573_ _01071_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_31 net606 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26100_ _05277_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__buf_2
X_23312_ _01311_ _02757_ _02734_ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__a21oi_1
XANTENNA_42 net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27080_ clknet_leaf_22_clk_sys _00697_ net607 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_20524_ _12054_ _12055_ VGND VGND VPWR VPWR _12373_ sky130_fd_sc_hd__nand2_1
X_24292_ _03299_ _03300_ _03623_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_133_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26031_ _05224_ VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23243_ _02660_ _02669_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__nor2_1
X_20455_ net287 _12108_ _12303_ VGND VGND VPWR VPWR _12304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23174_ _05717_ _07000_ _02644_ net882 VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__a22o_1
X_20386_ _12137_ _12234_ _12145_ VGND VGND VPWR VPWR _12235_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_18_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_18_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_22125_ _01063_ _01225_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22056_ _01615_ _01617_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__xor2_4
X_26933_ clknet_leaf_3_clk_sys _00550_ net583 VGND VGND VPWR VPWR top0.matmul0.cos\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21007_ _12697_ _12853_ net234 VGND VGND VPWR VPWR _12854_ sky130_fd_sc_hd__o21ai_1
X_26864_ clknet_leaf_41_clk_sys _00481_ net683 VGND VGND VPWR VPWR top0.svm0.tA\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_25815_ _05039_ _05040_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_199_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26795_ clknet_leaf_88_clk_sys _00412_ net642 VGND VGND VPWR VPWR top0.start_svm
+ sky130_fd_sc_hd__dfrtp_4
Xmax_cap11 net12 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
XFILLER_0_202_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13760_ _05971_ _05972_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__xnor2_2
X_22958_ _02306_ _02469_ _02309_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__a21o_1
X_25746_ net69 top0.matmul0.cos\[1\] _05458_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__and3_1
XFILLER_0_186_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21909_ _01412_ _01470_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__xnor2_2
X_13691_ _05883_ _05903_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__or2_1
X_22889_ _02313_ top0.svm0.tB\[15\] _02407_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__o21ai_1
X_25677_ top0.matmul0.sin\[10\] _04947_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15430_ _07251_ _07300_ VGND VGND VPWR VPWR _07529_ sky130_fd_sc_hd__and2_1
X_24628_ _03902_ _03903_ _03502_ _03981_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15361_ net534 _07444_ _07446_ _07459_ net479 VGND VGND VPWR VPWR _07460_ sky130_fd_sc_hd__o2111a_1
X_24559_ _03907_ _03913_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17100_ net812 _09115_ _09126_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__a21o_1
X_14312_ _06437_ _06438_ net30 net1015 VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18080_ _10063_ _10064_ VGND VGND VPWR VPWR _10065_ sky130_fd_sc_hd__and2b_1
X_15292_ _07344_ _07345_ VGND VGND VPWR VPWR _07391_ sky130_fd_sc_hd__xnor2_2
X_27278_ clknet_3_4__leaf_clk_mosi _00892_ VGND VGND VPWR VPWR spi0.data_packed\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14243_ net56 _06131_ _06282_ _06283_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__a22o_1
X_17031_ _05662_ _09081_ _08899_ VGND VGND VPWR VPWR _09083_ sky130_fd_sc_hd__or3_1
XFILLER_0_123_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26229_ _05346_ VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14174_ _06374_ _06370_ _06266_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18982_ net320 _10632_ VGND VGND VPWR VPWR _10956_ sky130_fd_sc_hd__and2_1
X_17933_ net351 net375 VGND VGND VPWR VPWR _09919_ sky130_fd_sc_hd__nand2_2
X_17864_ _09793_ _09849_ _09850_ VGND VGND VPWR VPWR _09851_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_178_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19603_ _11468_ _11473_ _11477_ VGND VGND VPWR VPWR _11492_ sky130_fd_sc_hd__or3_1
XFILLER_0_108_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16815_ _08881_ VGND VGND VPWR VPWR _08882_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17795_ _09649_ _09650_ _09781_ VGND VGND VPWR VPWR _09782_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_75_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19534_ _11423_ VGND VGND VPWR VPWR _11424_ sky130_fd_sc_hd__clkbuf_4
X_16746_ _08820_ _08829_ VGND VGND VPWR VPWR _08830_ sky130_fd_sc_hd__xnor2_1
X_13958_ _05790_ _05792_ VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__nor2_2
XFILLER_0_177_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19465_ _11359_ _11360_ VGND VGND VPWR VPWR _11361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16677_ _08758_ _08761_ VGND VGND VPWR VPWR _08762_ sky130_fd_sc_hd__xnor2_2
X_13889_ _06086_ _06087_ _06100_ _06101_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_158_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18416_ _10395_ _10297_ _10396_ VGND VGND VPWR VPWR _10397_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15628_ net496 net502 VGND VGND VPWR VPWR _07726_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19396_ top0.pid_d.curr_int\[1\] _11290_ _11293_ _11300_ VGND VGND VPWR VPWR _00327_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18347_ _10328_ VGND VGND VPWR VPWR _10329_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15559_ _07656_ _07657_ VGND VGND VPWR VPWR _07658_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18278_ net317 _10258_ _10259_ _10208_ VGND VGND VPWR VPWR _10260_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17229_ top0.pid_q.curr_int\[13\] _09140_ _09234_ _09135_ VGND VGND VPWR VPWR _09235_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20240_ net264 net279 VGND VGND VPWR VPWR _12089_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20171_ _12021_ _12022_ net207 VGND VGND VPWR VPWR _12023_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_161_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23930_ _03110_ _03100_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23861_ _03102_ _03105_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22812_ top0.svm0.counter\[4\] VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__inv_2
X_25600_ net750 _00000_ _04889_ _04891_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__o22a_1
XFILLER_0_196_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26580_ clknet_leaf_53_clk_sys _00203_ net672 VGND VGND VPWR VPWR top0.pid_q.prev_error\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_23792_ net568 top0.matmul0.matmul_stage_inst.b\[12\] top0.matmul0.matmul_stage_inst.a\[12\]
+ net564 VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__a22o_2
XFILLER_0_79_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25531_ top0.matmul0.b\[5\] top0.matmul0.matmul_stage_inst.f\[5\] _04846_ VGND VGND
+ VPWR VPWR _04852_ sky130_fd_sc_hd__mux2_1
X_22743_ _11954_ _11629_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25462_ _04572_ _04739_ _04742_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__or3b_1
XFILLER_0_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22674_ _02175_ _02176_ _02225_ _02184_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__o31a_1
XFILLER_0_192_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24413_ _03015_ _03016_ _03162_ _03163_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__o22a_1
X_27201_ clknet_leaf_91_clk_sys _00815_ net600 VGND VGND VPWR VPWR top0.cordic0.slte0.opB\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21625_ _01148_ _01156_ _01151_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__mux2_1
X_25393_ _04633_ _04736_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27132_ clknet_leaf_32_clk_sys _00746_ net664 VGND VGND VPWR VPWR top0.c_out_calc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_24344_ _03694_ _03700_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__xnor2_2
X_21556_ net105 net86 VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__xor2_2
XFILLER_0_106_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27063_ clknet_leaf_110_clk_sys _00680_ net578 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.c\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_20507_ _12341_ _12343_ _12355_ VGND VGND VPWR VPWR _12356_ sky130_fd_sc_hd__o21a_1
X_24275_ _03630_ _03632_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__nand2_1
X_21487_ _01022_ _01036_ _01050_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26014_ top0.b_in_matmul\[12\] _05211_ _05196_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__mux2_1
X_23226_ _01267_ _02669_ _02660_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__or3b_1
XFILLER_0_105_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20438_ net294 net287 VGND VGND VPWR VPWR _12287_ sky130_fd_sc_hd__and2b_2
XFILLER_0_31_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23157_ _05717_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__clkbuf_4
X_20369_ _12210_ _12211_ _12217_ VGND VGND VPWR VPWR _12218_ sky130_fd_sc_hd__or3b_1
X_22108_ _01637_ _01611_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__nor2b_1
X_23088_ _02542_ _02588_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__xnor2_1
X_22039_ net146 _01081_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__or2_1
X_14930_ _07041_ VGND VGND VPWR VPWR _07086_ sky130_fd_sc_hd__buf_4
X_26916_ clknet_leaf_2_clk_sys _00533_ net583 VGND VGND VPWR VPWR top0.matmul0.sin\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_26847_ clknet_leaf_43_clk_sys _00464_ net681 VGND VGND VPWR VPWR top0.svm0.delta\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_14861_ spi0.data_packed\[71\] top0.kpd\[7\] _07042_ VGND VGND VPWR VPWR _07050_
+ sky130_fd_sc_hd__mux2_1
X_16600_ _08681_ _08686_ _07710_ VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__o21a_1
XFILLER_0_199_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13812_ _05520_ _05521_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_11_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17580_ net420 VGND VGND VPWR VPWR _09567_ sky130_fd_sc_hd__inv_2
XFILLER_0_202_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14792_ _06951_ _06967_ VGND VGND VPWR VPWR _06993_ sky130_fd_sc_hd__nor2_1
X_26778_ clknet_leaf_6_clk_sys _00395_ net591 VGND VGND VPWR VPWR top0.cordic0.cos\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16531_ top0.pid_q.out\[12\] top0.pid_q.curr_int\[12\] VGND VGND VPWR VPWR _08618_
+ sky130_fd_sc_hd__nor2_1
X_13743_ _05947_ _05926_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__nand2_1
X_25729_ top0.matmul0.sin\[10\] _04983_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19250_ _11194_ _11185_ _11195_ VGND VGND VPWR VPWR _11196_ sky130_fd_sc_hd__a21o_1
X_16462_ net545 _08487_ _08488_ net549 _08550_ VGND VGND VPWR VPWR _08551_ sky130_fd_sc_hd__a32o_1
X_13674_ net50 _05496_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18201_ _10105_ _10110_ _10102_ VGND VGND VPWR VPWR _10184_ sky130_fd_sc_hd__o21a_1
X_15413_ _07489_ _07490_ _07508_ VGND VGND VPWR VPWR _07512_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19181_ top0.pid_d.prev_error\[1\] top0.pid_d.curr_error\[1\] VGND VGND VPWR VPWR
+ _11133_ sky130_fd_sc_hd__or2_1
X_16393_ _08482_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18132_ net342 net375 VGND VGND VPWR VPWR _10116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15344_ _07402_ _07412_ _07401_ VGND VGND VPWR VPWR _07443_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18063_ _10044_ _10047_ VGND VGND VPWR VPWR _10048_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_20_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15275_ net487 _07372_ _07373_ net1026 VGND VGND VPWR VPWR _07374_ sky130_fd_sc_hd__o211a_2
XFILLER_0_41_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold109 top0.svm0.tB\[12\] VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__dlygate4sd3_1
X_17014_ _05662_ top0.currT_r\[13\] _08899_ _09059_ net428 VGND VGND VPWR VPWR _09067_
+ sky130_fd_sc_hd__a2111o_1
X_14226_ _06436_ VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__buf_2
XFILLER_0_145_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14157_ _06359_ _06364_ _06367_ _06368_ VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__o22a_2
XFILLER_0_46_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14088_ _06296_ _06297_ _06298_ _06299_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__nor4_1
X_18965_ _10880_ _10886_ _10937_ _10938_ VGND VGND VPWR VPWR _10939_ sky130_fd_sc_hd__o211a_1
XFILLER_0_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17916_ _09826_ _09890_ VGND VGND VPWR VPWR _09902_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18896_ _10075_ _10870_ VGND VGND VPWR VPWR _10871_ sky130_fd_sc_hd__xor2_2
X_17847_ net339 net393 VGND VGND VPWR VPWR _09834_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17778_ net426 net315 VGND VGND VPWR VPWR _09765_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19517_ net303 VGND VGND VPWR VPWR _11407_ sky130_fd_sc_hd__inv_2
X_16729_ net452 net455 _08772_ VGND VGND VPWR VPWR _08813_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_202_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19448_ top0.pid_d.curr_int\[8\] top0.pid_d.prev_int\[8\] VGND VGND VPWR VPWR _11346_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19379_ net903 _11284_ _11287_ top0.pid_d.curr_error\[12\] VGND VGND VPWR VPWR _00322_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21410_ net236 _00976_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__xnor2_2
X_22390_ _11674_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21341_ _13130_ _13182_ VGND VGND VPWR VPWR _13183_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24060_ _03384_ _03401_ _03403_ _03417_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__a211o_1
X_21272_ _13029_ _13114_ _13031_ VGND VGND VPWR VPWR _13115_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23011_ _02514_ _02510_ _02374_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__o21a_1
X_20223_ net221 VGND VGND VPWR VPWR _12072_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_200_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20154_ spi0.data_packed\[15\] net211 _12006_ VGND VGND VPWR VPWR _12007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24962_ _04306_ _04312_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__xnor2_1
X_20085_ top0.cordic0.slte0.opA\[11\] _11785_ VGND VGND VPWR VPWR _11946_ sky130_fd_sc_hd__nor2_1
X_26701_ clknet_leaf_83_clk_sys net877 net649 VGND VGND VPWR VPWR top0.pid_d.prev_error\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_23913_ _03231_ _03266_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24893_ _04244_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26632_ clknet_leaf_74_clk_sys _00249_ net655 VGND VGND VPWR VPWR top0.pid_d.out\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_23844_ _03063_ _03064_ _03103_ _03104_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__o22a_1
XFILLER_0_170_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26563_ clknet_leaf_50_clk_sys _00186_ net671 VGND VGND VPWR VPWR top0.pid_q.curr_error\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_23775_ _03110_ _03130_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__and2_1
XFILLER_0_200_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20987_ net213 _12832_ _12833_ _12817_ _12773_ VGND VGND VPWR VPWR _12834_ sky130_fd_sc_hd__a311oi_1
X_25514_ top0.matmul0.matmul_stage_inst.mult1\[13\] _04710_ _03148_ VGND VGND VPWR
+ VPWR _04843_ sky130_fd_sc_hd__mux2_1
X_22726_ _02254_ _02275_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__xnor2_1
X_26494_ clknet_leaf_71_clk_sys _00117_ net657 VGND VGND VPWR VPWR top0.pid_d.prev_int\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_83_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25445_ _03722_ _04174_ _04518_ _04272_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__a211o_1
XFILLER_0_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22657_ _02208_ _02209_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21608_ _01162_ _01169_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13390_ top0.c_out_calc\[10\] _05464_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__nand2_4
X_25376_ _04691_ _04690_ _04718_ _04719_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__o22a_1
X_22588_ _02111_ _02114_ _02141_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27115_ clknet_leaf_89_clk_sys _00729_ net603 VGND VGND VPWR VPWR top0.clarke_done
+ sky130_fd_sc_hd__dfrtp_1
X_24327_ _03680_ _03683_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__xnor2_4
X_21539_ net118 _01100_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_50_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15060_ _07155_ _07158_ VGND VGND VPWR VPWR _07159_ sky130_fd_sc_hd__xnor2_2
X_24258_ _03536_ _03537_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__nand2_1
X_27046_ clknet_leaf_16_clk_sys _00663_ net612 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14011_ _06094_ _05543_ _05545_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__or3_1
X_23209_ _11526_ _02660_ net174 VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__o21a_1
X_24189_ _03540_ _03546_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18750_ _10725_ _10726_ VGND VGND VPWR VPWR _10727_ sky130_fd_sc_hd__or2_1
XFILLER_0_179_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15962_ _07913_ _07917_ _08056_ VGND VGND VPWR VPWR _08057_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17701_ net387 VGND VGND VPWR VPWR _09688_ sky130_fd_sc_hd__inv_2
X_14913_ _07077_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__clkbuf_1
X_18681_ net390 net387 _10495_ VGND VGND VPWR VPWR _10659_ sky130_fd_sc_hd__and3_1
X_15893_ _07888_ _07889_ _07988_ VGND VGND VPWR VPWR _07989_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_175_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17632_ _09608_ _09618_ VGND VGND VPWR VPWR _09619_ sky130_fd_sc_hd__xor2_2
X_14844_ net7 _07039_ _07040_ net744 VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__o22a_1
XFILLER_0_188_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17563_ net418 net340 VGND VGND VPWR VPWR _09550_ sky130_fd_sc_hd__nor2_1
X_14775_ net21 _05666_ VGND VGND VPWR VPWR _06976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19302_ net437 _11240_ _11243_ _11125_ VGND VGND VPWR VPWR _11244_ sky130_fd_sc_hd__a211o_1
XFILLER_0_105_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16514_ _08600_ _08601_ VGND VGND VPWR VPWR _08602_ sky130_fd_sc_hd__or2_1
X_13726_ net47 _05683_ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__nand2_1
X_17494_ _09411_ _09412_ VGND VGND VPWR VPWR _09481_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19233_ top0.matmul0.alpha_pass\[4\] net76 _11150_ top0.matmul0.alpha_pass\[6\] VGND
+ VGND VPWR VPWR _11181_ sky130_fd_sc_hd__o31ai_2
X_16445_ net468 net473 net476 _08286_ VGND VGND VPWR VPWR _08534_ sky130_fd_sc_hd__nand4_2
X_13657_ net1027 _05478_ _05479_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19164_ top0.pid_d.prev_error\[0\] top0.pid_d.curr_error\[0\] VGND VGND VPWR VPWR
+ _11118_ sky130_fd_sc_hd__xor2_1
XFILLER_0_147_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16376_ _08463_ _08465_ VGND VGND VPWR VPWR _08466_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13588_ _05649_ _05800_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_182_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18115_ net332 net389 VGND VGND VPWR VPWR _10099_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15327_ _07418_ _07423_ _07425_ VGND VGND VPWR VPWR _07426_ sky130_fd_sc_hd__o21ba_1
X_19095_ _11065_ _11066_ VGND VGND VPWR VPWR _11067_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18046_ _09919_ _09920_ _10030_ VGND VGND VPWR VPWR _10031_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_197_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15258_ net524 net495 VGND VGND VPWR VPWR _07357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14209_ _06317_ _06318_ _06338_ _06328_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15189_ _07188_ _07189_ _07287_ VGND VGND VPWR VPWR _07288_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_111_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout408 top0.pid_d.mult0.a\[5\] VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__clkbuf_4
Xfanout419 net420 VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__clkbuf_2
X_19997_ _11774_ _11861_ _11862_ _11863_ VGND VGND VPWR VPWR _11864_ sky130_fd_sc_hd__a31o_1
X_18948_ _10922_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18879_ net383 _10852_ _10853_ VGND VGND VPWR VPWR _10854_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_154_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20910_ net265 _12095_ _12715_ VGND VGND VPWR VPWR _12758_ sky130_fd_sc_hd__nor3_1
X_21890_ _01366_ _01407_ _01451_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__a21oi_1
X_20841_ _12215_ _12688_ _12689_ VGND VGND VPWR VPWR _12690_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_194_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23560_ _02946_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__clkbuf_1
X_20772_ _11527_ _12109_ VGND VGND VPWR VPWR _12621_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout15 net530 VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__clkbuf_4
Xfanout26 net27 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_175_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22511_ _01821_ _02065_ _02066_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__o21ai_4
Xfanout37 net38 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_4
Xfanout48 net49 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
X_23491_ _02910_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__clkbuf_1
Xfanout59 top0.periodTop_r\[2\] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_4
XFILLER_0_18_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25230_ _04512_ _04572_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__xnor2_1
X_22442_ _01809_ _01891_ _01998_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__and3_1
XFILLER_0_190_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25161_ _03355_ _04252_ _03502_ _04339_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__a31o_2
XFILLER_0_33_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22373_ _01909_ _01930_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__nand2_1
X_24112_ _03396_ _03469_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21324_ net242 _13124_ VGND VGND VPWR VPWR _13166_ sky130_fd_sc_hd__and2_1
X_25092_ _04437_ _04440_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24043_ _03398_ _03400_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__nor2_1
X_21255_ _12965_ _13007_ VGND VGND VPWR VPWR _13099_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20206_ _12052_ _12053_ _12041_ VGND VGND VPWR VPWR _12055_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21186_ _12207_ _13029_ net262 VGND VGND VPWR VPWR _13030_ sky130_fd_sc_hd__mux2_1
X_20137_ net212 _11413_ _11519_ VGND VGND VPWR VPWR _11993_ sky130_fd_sc_hd__and3_1
X_25994_ _05164_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__buf_4
XFILLER_0_99_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24945_ _04199_ _04200_ _04201_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__a21o_1
X_20068_ _11903_ _11929_ net181 VGND VGND VPWR VPWR _11930_ sky130_fd_sc_hd__a21oi_1
X_24876_ _04021_ _04022_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__nor2_1
X_26615_ clknet_leaf_27_clk_sys _00232_ net621 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_23827_ _03027_ _03028_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__nor2_4
XFILLER_0_185_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14560_ _06707_ _06709_ _06765_ VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__a21o_1
X_26546_ clknet_leaf_49_clk_sys _00169_ net675 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23758_ _03036_ _03037_ _03069_ _03071_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__o22a_1
XFILLER_0_184_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13511_ _05617_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_165_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22709_ _02258_ _02259_ _02171_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__a21o_1
X_14491_ _06636_ _06650_ _06638_ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26477_ clknet_leaf_89_clk_sys _00108_ net603 VGND VGND VPWR VPWR top0.periodTop\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_23689_ _03045_ _03046_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__nor2_2
XFILLER_0_55_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16230_ top0.pid_q.out\[7\] _08321_ _07700_ VGND VGND VPWR VPWR _08322_ sky130_fd_sc_hd__mux2_1
X_25428_ _04743_ _04744_ _04518_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__a21o_1
X_13442_ _05548_ _05555_ _05654_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_181_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13373_ _05585_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__buf_4
X_16161_ _08219_ _08223_ _08217_ VGND VGND VPWR VPWR _08253_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25359_ _04521_ _04645_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15112_ _07149_ _07159_ _07154_ VGND VGND VPWR VPWR _07211_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16092_ net529 net443 VGND VGND VPWR VPWR _08185_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_121_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27029_ clknet_3_3__leaf_clk_sys _00646_ net615 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_15043_ net917 _07139_ _07143_ top0.pid_d.curr_int\[13\] VGND VGND VPWR VPWR _00130_
+ sky130_fd_sc_hd__a22o_1
X_19920_ _11791_ _11792_ VGND VGND VPWR VPWR _11793_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19851_ _11717_ _11719_ VGND VGND VPWR VPWR _11728_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_66_clk_sys clknet_3_5__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_66_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_107_clk_sys clknet_3_0__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_107_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_177_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18802_ net371 net318 VGND VGND VPWR VPWR _10778_ sky130_fd_sc_hd__nand2_1
X_19782_ _11661_ _11663_ VGND VGND VPWR VPWR _11664_ sky130_fd_sc_hd__xnor2_2
X_16994_ _09027_ _09047_ _09048_ VGND VGND VPWR VPWR _09049_ sky130_fd_sc_hd__o21a_1
X_18733_ net327 net362 VGND VGND VPWR VPWR _10710_ sky130_fd_sc_hd__nand2_1
X_15945_ _07944_ _07959_ _07960_ VGND VGND VPWR VPWR _08040_ sky130_fd_sc_hd__o21a_1
X_18664_ _10633_ _10641_ VGND VGND VPWR VPWR _10642_ sky130_fd_sc_hd__xnor2_1
X_15876_ _07821_ _07822_ _07971_ VGND VGND VPWR VPWR _07972_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_116_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17615_ _09547_ _09548_ _09601_ VGND VGND VPWR VPWR _09602_ sky130_fd_sc_hd__a21o_1
X_14827_ _07025_ _07026_ VGND VGND VPWR VPWR _07027_ sky130_fd_sc_hd__or2b_1
XFILLER_0_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18595_ _10490_ _10502_ _10492_ VGND VGND VPWR VPWR _10574_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_25_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17546_ net407 _09530_ _09532_ net412 VGND VGND VPWR VPWR _09533_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14758_ _06957_ _06959_ VGND VGND VPWR VPWR _06960_ sky130_fd_sc_hd__xor2_2
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13709_ _05909_ _05921_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__nand2_1
X_17477_ net398 _09462_ _09463_ net400 VGND VGND VPWR VPWR _09464_ sky130_fd_sc_hd__a22o_1
X_14689_ _06887_ _06892_ VGND VGND VPWR VPWR _06893_ sky130_fd_sc_hd__xor2_1
XFILLER_0_157_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19216_ _11164_ _11156_ top0.pid_d.prev_error\[4\] VGND VGND VPWR VPWR _11165_ sky130_fd_sc_hd__o21ba_1
X_16428_ _08430_ _08432_ _08516_ VGND VGND VPWR VPWR _08517_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19147_ top0.kid\[8\] _11098_ _11100_ top0.kpd\[8\] VGND VGND VPWR VPWR _11109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16359_ _07493_ _08448_ VGND VGND VPWR VPWR _08449_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19078_ _10845_ _11047_ _11048_ _11049_ VGND VGND VPWR VPWR _11050_ sky130_fd_sc_hd__o31a_1
XFILLER_0_30_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18029_ _09910_ _09911_ _09912_ VGND VGND VPWR VPWR _10014_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21040_ _12879_ _12880_ _12882_ _12883_ _12886_ VGND VGND VPWR VPWR _12887_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout205 top0.state\[2\] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_2
Xfanout216 net217 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_2
Xfanout227 net228 VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_4
Xfanout238 net239 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__buf_4
XFILLER_0_10_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout249 top0.cordic0.vec\[0\]\[10\] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__buf_4
XFILLER_0_66_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22991_ _02497_ _02493_ _02360_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__o21a_1
X_24730_ _03883_ _03884_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__nor2_1
X_21942_ net151 net136 net165 VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24661_ _03057_ _03058_ _03717_ _03718_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__o22a_1
X_21873_ _01379_ _01434_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_173_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26400_ clknet_leaf_98_clk_sys _00041_ net588 VGND VGND VPWR VPWR top0.kpd\[5\] sky130_fd_sc_hd__dfrtp_1
X_23612_ top0.matmul0.alpha_pass\[13\] _09325_ net560 VGND VGND VPWR VPWR _02973_
+ sky130_fd_sc_hd__mux2_1
X_20824_ _12669_ _12672_ VGND VGND VPWR VPWR _12673_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24592_ _03931_ _03946_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26331_ _05397_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23543_ top0.a_in_matmul\[11\] top0.matmul0.a\[11\] _02937_ VGND VGND VPWR VPWR _02938_
+ sky130_fd_sc_hd__mux2_1
X_20755_ _12598_ _12601_ _12603_ net287 VGND VGND VPWR VPWR _12604_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_9_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26262_ spi0.data_packed\[29\] spi0.data_packed\[30\] net696 VGND VGND VPWR VPWR
+ _05363_ sky130_fd_sc_hd__mux2_1
X_23474_ _02901_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20686_ _12324_ _12534_ VGND VGND VPWR VPWR _12535_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_119_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25213_ _03363_ _04131_ _04559_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__a21o_1
X_22425_ _01979_ _01982_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__xor2_1
XFILLER_0_169_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26193_ _05326_ top0.cordic0.slte0.opB\[14\] _12003_ VGND VGND VPWR VPWR _05327_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25144_ _04427_ _04432_ _04491_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22356_ net138 net123 _01910_ _01914_ top0.cordic0.vec\[1\]\[9\] VGND VGND VPWR VPWR
+ _01915_ sky130_fd_sc_hd__a311o_1
XFILLER_0_20_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21307_ _13142_ _13149_ VGND VGND VPWR VPWR _13150_ sky130_fd_sc_hd__xnor2_2
X_25075_ _04420_ _04423_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__xnor2_1
X_22287_ net101 net86 net96 VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__o21ai_1
X_24026_ _03379_ _03383_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__and2_2
Xhold270 top0.pid_q.prev_int\[9\] VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__dlygate4sd3_1
X_21238_ _12628_ VGND VGND VPWR VPWR _13082_ sky130_fd_sc_hd__inv_2
Xhold281 top0.cordic0.slte0.opA\[4\] VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 top0.cordic0.slte0.opA\[2\] VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__dlygate4sd3_1
X_21169_ net731 _12813_ _13013_ _12963_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13991_ _06181_ _06203_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__xnor2_2
X_25977_ top0.matmul0.beta_pass\[4\] _05169_ _05182_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15730_ _07745_ _07747_ _07743_ VGND VGND VPWR VPWR _07827_ sky130_fd_sc_hd__a21bo_1
X_24928_ _02982_ _04097_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15661_ _07753_ _07758_ VGND VGND VPWR VPWR _07759_ sky130_fd_sc_hd__xor2_1
X_24859_ _04198_ _04210_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17400_ net334 top0.pid_d.mult0.a\[0\] VGND VGND VPWR VPWR _09387_ sky130_fd_sc_hd__nand2_1
X_14612_ _06551_ _06807_ _06816_ VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__a21o_1
XFILLER_0_197_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18380_ _10358_ _10360_ VGND VGND VPWR VPWR _10361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15592_ _07220_ _07298_ VGND VGND VPWR VPWR _07691_ sky130_fd_sc_hd__or2_1
X_17331_ _09321_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14543_ _06699_ _06736_ _06738_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__a21o_2
X_26529_ clknet_leaf_61_clk_sys _00152_ net651 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17262_ _09262_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__clkbuf_1
X_14474_ _06672_ _06681_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_71_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19001_ _10972_ _10974_ VGND VGND VPWR VPWR _10975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16213_ _08182_ _08215_ _08214_ VGND VGND VPWR VPWR _08305_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13425_ top0.matmul0.beta_pass\[9\] _05466_ _05470_ _05463_ top0.c_out_calc\[9\]
+ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__a32o_1
X_17193_ _09201_ _09195_ _09202_ VGND VGND VPWR VPWR _09203_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16144_ top0.pid_q.out\[6\] _07704_ VGND VGND VPWR VPWR _08237_ sky130_fd_sc_hd__nor2_1
X_13356_ _05513_ _05514_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16075_ net476 net499 VGND VGND VPWR VPWR _08168_ sky130_fd_sc_hd__nand2_2
X_13287_ net33 VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__clkinv_4
X_19903_ _11575_ net82 _11776_ VGND VGND VPWR VPWR _11777_ sky130_fd_sc_hd__mux2_1
X_15026_ top0.pid_d.state\[0\] top0.pid_d.state\[3\] _07136_ VGND VGND VPWR VPWR _07141_
+ sky130_fd_sc_hd__nor3_2
X_19834_ net244 _11705_ VGND VGND VPWR VPWR _11712_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16977_ top0.currT_r\[9\] top0.currT_r\[10\] _08997_ _09032_ _05601_ VGND VGND VPWR
+ VPWR _09033_ sky130_fd_sc_hd__o32a_2
X_19765_ net180 _11413_ VGND VGND VPWR VPWR _11648_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15928_ _08021_ _08022_ VGND VGND VPWR VPWR _08023_ sky130_fd_sc_hd__xor2_2
X_18716_ net376 net316 VGND VGND VPWR VPWR _10693_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19696_ _11424_ _11528_ _11540_ _11565_ VGND VGND VPWR VPWR _11582_ sky130_fd_sc_hd__or4b_2
X_18647_ _10621_ _10624_ VGND VGND VPWR VPWR _10625_ sky130_fd_sc_hd__nand2_1
X_15859_ _07849_ _07851_ _07850_ VGND VGND VPWR VPWR _07955_ sky130_fd_sc_hd__o21a_1
XFILLER_0_188_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18578_ _10481_ _10485_ _10556_ VGND VGND VPWR VPWR _10557_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17529_ _09448_ _09449_ _09515_ VGND VGND VPWR VPWR _09516_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20540_ _12372_ _12276_ VGND VGND VPWR VPWR _12389_ sky130_fd_sc_hd__or2_1
XFILLER_0_188_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20471_ _11726_ _12246_ _12318_ VGND VGND VPWR VPWR _12320_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_144_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22210_ _01113_ _01770_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__xor2_2
XFILLER_0_70_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23190_ _02646_ _06860_ _02649_ net814 VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22141_ _01311_ _01076_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22072_ _01568_ _01588_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__and2b_1
XFILLER_0_199_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25900_ net429 _05116_ _05114_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__a21o_1
X_21023_ _12869_ _12783_ _12708_ VGND VGND VPWR VPWR _12870_ sky130_fd_sc_hd__o21a_1
X_26880_ clknet_leaf_41_clk_sys _00497_ net685 VGND VGND VPWR VPWR top0.svm0.tB\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_25831_ _05053_ _05054_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25762_ top0.matmul0.matmul_stage_inst.a\[9\] _04898_ _05457_ VGND VGND VPWR VPWR
+ _05002_ sky130_fd_sc_hd__mux2_1
X_22974_ net170 _02483_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_198_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24713_ _04049_ _04056_ _04065_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__o21a_1
X_21925_ net156 net137 VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__nand2_1
X_25693_ _05457_ _04958_ _04959_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__and3_1
XFILLER_0_179_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24644_ _03024_ _03025_ _03069_ _03071_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_6_clk_sys clknet_3_2__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_6_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_14_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_14_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_21856_ _01268_ _01413_ _01417_ net152 VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__a22o_2
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20807_ net273 _11673_ _12559_ _12650_ _12655_ VGND VGND VPWR VPWR _12656_ sky130_fd_sc_hd__a32o_1
XFILLER_0_72_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24575_ _03783_ _03814_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21787_ net132 net118 _01065_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__a21o_1
XFILLER_0_182_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26314_ spi0.data_packed\[55\] spi0.data_packed\[56\] net698 VGND VGND VPWR VPWR
+ _05389_ sky130_fd_sc_hd__mux2_1
X_23526_ top0.a_in_matmul\[3\] top0.matmul0.a\[3\] _02926_ VGND VGND VPWR VPWR _02929_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20738_ _12284_ _12585_ _12586_ _12285_ VGND VGND VPWR VPWR _12587_ sky130_fd_sc_hd__a22o_1
X_27294_ clknet_3_0__leaf_clk_mosi _00908_ VGND VGND VPWR VPWR spi0.opcode\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26245_ _05354_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20669_ _12471_ _12482_ _12477_ VGND VGND VPWR VPWR _12518_ sky130_fd_sc_hd__o21bai_1
X_23457_ _11789_ _02891_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13210_ _05435_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__buf_4
X_22408_ _01771_ _01965_ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__xnor2_2
X_14190_ _06289_ _06399_ _06400_ VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__o21a_1
X_26176_ _05313_ VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__clkbuf_1
X_23388_ _02809_ _02818_ _02828_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25127_ _04419_ _04452_ _04453_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__o21a_2
X_22339_ _01863_ _01865_ _01897_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25058_ _04406_ _04396_ _04394_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__o21a_1
X_16900_ top0.currT_r\[6\] _08960_ VGND VGND VPWR VPWR _08961_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_76_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24009_ _03195_ _03250_ _03217_ VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__or3_1
X_17880_ net378 net355 net375 net359 VGND VGND VPWR VPWR _09867_ sky130_fd_sc_hd__nand4_1
XFILLER_0_40_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16831_ _08895_ _08896_ VGND VGND VPWR VPWR _08897_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_189_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout580 net581 VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__clkbuf_4
X_19550_ _11430_ VGND VGND VPWR VPWR _11439_ sky130_fd_sc_hd__clkbuf_2
Xfanout591 net598 VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__clkbuf_4
X_16762_ _08794_ _08844_ _08845_ VGND VGND VPWR VPWR _08846_ sky130_fd_sc_hd__a21o_1
X_13974_ net51 _05605_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__nand2_1
X_18501_ _10369_ _10378_ _10377_ VGND VGND VPWR VPWR _10481_ sky130_fd_sc_hd__a21oi_2
X_15713_ _07793_ _07807_ _07809_ _07792_ VGND VGND VPWR VPWR _07810_ sky130_fd_sc_hd__a31o_2
XFILLER_0_87_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19481_ _10905_ _11374_ VGND VGND VPWR VPWR _11375_ sky130_fd_sc_hd__xnor2_1
X_16693_ _08757_ _08776_ VGND VGND VPWR VPWR _08778_ sky130_fd_sc_hd__and2_1
X_18432_ _10308_ _10412_ _10229_ VGND VGND VPWR VPWR _10413_ sky130_fd_sc_hd__o21a_1
X_15644_ _07740_ _07741_ VGND VGND VPWR VPWR _07742_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_85_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18363_ _10331_ _10343_ VGND VGND VPWR VPWR _10344_ sky130_fd_sc_hd__nor2_1
X_15575_ _07564_ _07583_ VGND VGND VPWR VPWR _07674_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17314_ top0.matmul0.matmul_stage_inst.mult1\[10\] top0.matmul0.matmul_stage_inst.mult2\[10\]
+ VGND VGND VPWR VPWR _09307_ sky130_fd_sc_hd__xor2_1
XFILLER_0_200_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14526_ net45 _06268_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18294_ _10175_ _10177_ _10176_ VGND VGND VPWR VPWR _10276_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17245_ top0.pid_q.curr_int\[15\] _09140_ _09192_ _08849_ VGND VGND VPWR VPWR _09249_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14457_ _06596_ _06594_ VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13408_ _05620_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__buf_2
XFILLER_0_52_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17176_ top0.pid_q.curr_int\[7\] top0.pid_q.prev_int\[7\] VGND VGND VPWR VPWR _09188_
+ sky130_fd_sc_hd__xor2_1
X_14388_ net51 _06268_ VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16127_ net483 _08003_ net499 VGND VGND VPWR VPWR _08220_ sky130_fd_sc_hd__o21a_2
XFILLER_0_49_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13339_ net57 _05551_ _05549_ _05550_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_122_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_94_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16058_ _08149_ _08151_ VGND VGND VPWR VPWR _08152_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15009_ spi0.data_packed\[10\] top0.periodTop\[10\] _07125_ VGND VGND VPWR VPWR _07130_
+ sky130_fd_sc_hd__mux2_1
X_19817_ _11695_ _11696_ VGND VGND VPWR VPWR _11697_ sky130_fd_sc_hd__and2b_1
XFILLER_0_155_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19748_ net180 _11630_ VGND VGND VPWR VPWR _11631_ sky130_fd_sc_hd__or2_1
X_19679_ _11424_ _11528_ _11540_ _11512_ VGND VGND VPWR VPWR _11566_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_155_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21710_ net162 net141 _01268_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__or3_1
XFILLER_0_63_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22690_ _02237_ _02240_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21641_ net144 _01101_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24360_ net571 net575 top0.matmul0.matmul_stage_inst.f\[14\] VGND VGND VPWR VPWR
+ _03717_ sky130_fd_sc_hd__o21a_2
XFILLER_0_117_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21572_ net114 _01074_ _01132_ _01122_ _01133_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__a221o_2
XFILLER_0_75_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_10 net1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_21 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_32 _03110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_191_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_43 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20523_ _12370_ _12371_ VGND VGND VPWR VPWR _12372_ sky130_fd_sc_hd__xor2_4
X_23311_ _11512_ _02741_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__xnor2_1
X_24291_ _03624_ _03625_ _03635_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26030_ top0.a_in_matmul\[0\] _05223_ _05196_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20454_ _12301_ _12302_ VGND VGND VPWR VPWR _12303_ sky130_fd_sc_hd__nand2_1
X_23242_ _11425_ _02691_ _02668_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_63_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23173_ _05717_ _06971_ _02644_ net806 VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__a22o_1
XFILLER_0_160_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20385_ _12139_ _12141_ VGND VGND VPWR VPWR _12234_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22124_ _01215_ _01219_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22055_ net102 _01616_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__nand2_2
X_26932_ clknet_leaf_7_clk_sys _00549_ net593 VGND VGND VPWR VPWR top0.matmul0.cos\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_21006_ net225 net222 VGND VGND VPWR VPWR _12853_ sky130_fd_sc_hd__nor2b_2
X_26863_ clknet_leaf_41_clk_sys _00480_ net683 VGND VGND VPWR VPWR top0.svm0.tA\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25814_ _05034_ _05033_ _05035_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__mux2_1
X_26794_ clknet_leaf_92_clk_sys _00411_ net599 VGND VGND VPWR VPWR top0.cordic0.out_valid
+ sky130_fd_sc_hd__dfrtp_2
Xmax_cap12 _05066_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_173_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25745_ _04993_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22957_ _02466_ _02468_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_195_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21908_ _01393_ _01436_ _01438_ _01392_ _01469_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__o221a_1
XFILLER_0_179_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13690_ _05886_ _05899_ _05902_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__o21a_1
X_25676_ _04884_ _04942_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__and2_1
X_22888_ _02313_ top0.svm0.tB\[15\] top0.svm0.tB\[14\] _02404_ _02406_ VGND VGND VPWR
+ VPWR _02407_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24627_ _03150_ _03151_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__or2_2
XFILLER_0_38_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21839_ _01384_ _01391_ _01400_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_77_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15360_ net486 _07456_ _07458_ net537 VGND VGND VPWR VPWR _07459_ sky130_fd_sc_hd__o211a_1
X_24558_ _03909_ _03912_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14311_ _06517_ _06520_ VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23509_ top0.cordic0.cos\[9\] top0.matmul0.cos\[9\] _02915_ VGND VGND VPWR VPWR _02920_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27277_ clknet_3_5__leaf_clk_mosi _00891_ VGND VGND VPWR VPWR spi0.data_packed\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_15291_ _07365_ _07389_ VGND VGND VPWR VPWR _07390_ sky130_fd_sc_hd__xor2_2
XFILLER_0_108_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24489_ _03842_ _03844_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17030_ _09081_ top0.currT_r\[13\] _08899_ VGND VGND VPWR VPWR _09082_ sky130_fd_sc_hd__or3_1
X_14242_ _06295_ _06452_ _06301_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__a21o_1
X_26228_ spi0.data_packed\[12\] spi0.data_packed\[13\] net695 VGND VGND VPWR VPWR
+ _05346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14173_ _06273_ _06382_ _06383_ _06257_ VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__o22a_1
XFILLER_0_180_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26159_ net18 _05299_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18981_ _10632_ _10878_ net363 VGND VGND VPWR VPWR _10955_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_21_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17932_ _09833_ _09838_ _09917_ VGND VGND VPWR VPWR _09918_ sky130_fd_sc_hd__a21o_1
XFILLER_0_175_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17863_ net389 net346 net384 net351 VGND VGND VPWR VPWR _09850_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19602_ _11486_ _11490_ top0.cordic0.slte0.opA\[9\] VGND VGND VPWR VPWR _11491_ sky130_fd_sc_hd__a21oi_1
X_16814_ _08880_ VGND VGND VPWR VPWR _08881_ sky130_fd_sc_hd__buf_2
X_17794_ _09649_ _09650_ _09648_ VGND VGND VPWR VPWR _09781_ sky130_fd_sc_hd__o21ai_1
X_16745_ _08648_ _08828_ VGND VGND VPWR VPWR _08829_ sky130_fd_sc_hd__xor2_1
X_19533_ _11414_ _11421_ _11422_ VGND VGND VPWR VPWR _11423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13957_ _06085_ _06169_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__xor2_2
XFILLER_0_88_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19464_ top0.pid_d.curr_int\[10\] top0.pid_d.prev_int\[10\] VGND VGND VPWR VPWR _11360_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16676_ _08759_ _08760_ VGND VGND VPWR VPWR _08761_ sky130_fd_sc_hd__xor2_1
X_13888_ _06099_ _06092_ _06093_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__and3_1
XFILLER_0_159_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18415_ _10395_ _10297_ _10286_ VGND VGND VPWR VPWR _10396_ sky130_fd_sc_hd__a21o_1
X_15627_ _07624_ _07625_ _07724_ VGND VGND VPWR VPWR _07725_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_201_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19395_ net431 _09977_ _11299_ net442 _11129_ VGND VGND VPWR VPWR _11300_ sky130_fd_sc_hd__a221o_1
XFILLER_0_174_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18346_ _10238_ _10239_ _10327_ VGND VGND VPWR VPWR _10328_ sky130_fd_sc_hd__a21o_1
X_15558_ _07648_ _07655_ VGND VGND VPWR VPWR _07657_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14509_ _06212_ _06715_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__nor2_1
XFILLER_0_173_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18277_ net396 net317 VGND VGND VPWR VPWR _10259_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15489_ _07194_ _07295_ VGND VGND VPWR VPWR _07588_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17228_ net551 _09055_ _09233_ net554 VGND VGND VPWR VPWR _09234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17159_ top0.pid_q.curr_int\[5\] top0.pid_q.prev_int\[5\] VGND VGND VPWR VPWR _09173_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20170_ top0.cordic0.out_valid top0.cordic_done VGND VGND VPWR VPWR _12022_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23860_ _03102_ _03105_ _03124_ _03217_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_79_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22811_ top0.svm0.counter\[5\] VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__inv_2
X_23791_ top0.matmul0.matmul_stage_inst.f\[0\] _03146_ _03148_ top0.matmul0.matmul_stage_inst.e\[0\]
+ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_149_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25530_ _04851_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__clkbuf_1
X_22742_ net191 _02286_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_181_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25461_ _04742_ _04739_ _04572_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__and3b_1
XFILLER_0_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22673_ _02207_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27200_ clknet_leaf_91_clk_sys _00814_ net600 VGND VGND VPWR VPWR top0.cordic0.slte0.opB\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24412_ _03185_ _03743_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__nor2_2
X_21624_ _01147_ _01185_ _01148_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_63_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25392_ _04734_ _04735_ _04518_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_191_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27131_ clknet_leaf_33_clk_sys _00745_ net664 VGND VGND VPWR VPWR top0.c_out_calc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24343_ _03698_ _03699_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__nor2_1
X_21555_ net109 _01115_ _01116_ VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27062_ clknet_leaf_110_clk_sys _00679_ net578 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.c\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_20506_ _12299_ _12354_ VGND VGND VPWR VPWR _12355_ sky130_fd_sc_hd__xnor2_1
X_24274_ _03626_ _03631_ _03623_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_50_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21486_ _01022_ _01036_ _01033_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26013_ top0.matmul0.beta_pass\[12\] _05203_ _05210_ VGND VGND VPWR VPWR _05211_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20437_ _12284_ _12285_ net274 VGND VGND VPWR VPWR _12286_ sky130_fd_sc_hd__mux2_1
X_23225_ net161 _02674_ _02675_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_114_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23156_ net902 _06381_ _02639_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__o21a_1
X_20368_ _12040_ _12216_ VGND VGND VPWR VPWR _12217_ sky130_fd_sc_hd__xnor2_2
X_22107_ _01406_ _01608_ _01363_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__o21ba_1
X_23087_ net36 top0.svm0.counter\[11\] VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__xor2_1
X_20299_ _12137_ _12146_ _12147_ VGND VGND VPWR VPWR _12148_ sky130_fd_sc_hd__nand3_2
X_22038_ net122 net113 net106 _01596_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__a31o_1
X_26915_ clknet_leaf_7_clk_sys _00532_ net583 VGND VGND VPWR VPWR top0.matmul0.sin\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_26846_ clknet_leaf_44_clk_sys _00463_ net681 VGND VGND VPWR VPWR top0.svm0.delta\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14860_ _07049_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13811_ net62 _06023_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__nand2_1
X_14791_ _06942_ VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__clkinvlp_2
X_26777_ clknet_leaf_7_clk_sys _00394_ net593 VGND VGND VPWR VPWR top0.cordic0.cos\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_23989_ _03317_ _03318_ _03313_ _03315_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16530_ _08610_ _08617_ _07710_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__o21a_1
X_13742_ _05949_ _05954_ _05860_ _05908_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25728_ net74 _04942_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__nand2_1
X_16461_ _08491_ _08549_ VGND VGND VPWR VPWR _08550_ sky130_fd_sc_hd__xnor2_2
X_13673_ _05884_ _05885_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__xnor2_2
X_25659_ net71 top0.matmul0.sin\[6\] VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18200_ _10172_ _10182_ VGND VGND VPWR VPWR _10183_ sky130_fd_sc_hd__xor2_2
XFILLER_0_35_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15412_ _07489_ _07479_ _07490_ VGND VGND VPWR VPWR _07511_ sky130_fd_sc_hd__or3_1
XFILLER_0_66_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19180_ _11125_ _11129_ _11131_ _11132_ _07800_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__o311a_1
XFILLER_0_26_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16392_ net1018 _08481_ VGND VGND VPWR VPWR _08482_ sky130_fd_sc_hd__and2_1
XFILLER_0_182_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_159_Left_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18131_ net350 top0.pid_d.mult0.a\[14\] VGND VGND VPWR VPWR _10115_ sky130_fd_sc_hd__nand2_2
XFILLER_0_136_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15343_ _07434_ _07435_ _07440_ _07441_ VGND VGND VPWR VPWR _07442_ sky130_fd_sc_hd__or4_2
XFILLER_0_109_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18062_ _10045_ _10046_ VGND VGND VPWR VPWR _10047_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15274_ net524 net495 net491 net527 VGND VGND VPWR VPWR _07373_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17013_ _05662_ top0.currT_r\[13\] _05437_ _09059_ net428 VGND VGND VPWR VPWR _09066_
+ sky130_fd_sc_hd__o2111a_1
X_14225_ net28 _05520_ _05521_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__and3_1
XFILLER_0_184_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14156_ _06239_ _06251_ _06252_ _06366_ VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14087_ _06189_ _06196_ VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__nor2_1
X_18964_ _10880_ _10885_ _10723_ VGND VGND VPWR VPWR _10938_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_168_Left_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17915_ top0.pid_d.out\[0\] top0.pid_d.curr_int\[0\] _09899_ VGND VGND VPWR VPWR
+ _09901_ sky130_fd_sc_hd__nand3_1
X_18895_ net318 net370 VGND VGND VPWR VPWR _10870_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17846_ _09783_ _09784_ _09832_ VGND VGND VPWR VPWR _09833_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_135_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14989_ _07119_ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__clkbuf_1
X_17777_ _09636_ _09762_ _09763_ VGND VGND VPWR VPWR _09764_ sky130_fd_sc_hd__a21o_1
X_19516_ _11341_ _11398_ _11404_ _11292_ _11406_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__a221o_1
XFILLER_0_152_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16728_ net447 _08811_ VGND VGND VPWR VPWR _08812_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19447_ top0.pid_d.curr_int\[7\] _11343_ _11344_ VGND VGND VPWR VPWR _11345_ sky130_fd_sc_hd__o21ai_2
X_16659_ net16 _08744_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__nor2_1
XFILLER_0_202_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_177_Left_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19378_ top0.pid_d.prev_error\[11\] _11284_ _11287_ net760 VGND VGND VPWR VPWR _00321_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18329_ net310 VGND VGND VPWR VPWR _10311_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21340_ _13169_ _13181_ VGND VGND VPWR VPWR _13182_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21271_ net246 _13028_ VGND VGND VPWR VPWR _13114_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23010_ top0.svm0.delta\[12\] VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20222_ _12054_ _12055_ _12060_ VGND VGND VPWR VPWR _12071_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20153_ _12003_ VGND VGND VPWR VPWR _12006_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24961_ _04307_ _04231_ _04309_ _04069_ _04311_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__a221o_1
X_20084_ net1014 _11944_ net177 VGND VGND VPWR VPWR _11945_ sky130_fd_sc_hd__o21ai_1
X_26700_ clknet_leaf_62_clk_sys net881 net648 VGND VGND VPWR VPWR top0.pid_d.prev_error\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_23912_ _03231_ _03266_ _03269_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__a21oi_1
X_24892_ top0.matmul0.matmul_stage_inst.mult2\[6\] _04243_ _03642_ VGND VGND VPWR
+ VPWR _04244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26631_ clknet_leaf_82_clk_sys _00248_ net637 VGND VGND VPWR VPWR top0.pid_d.out\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_23843_ _03114_ _03200_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26562_ clknet_leaf_51_clk_sys _00185_ net671 VGND VGND VPWR VPWR top0.pid_q.curr_error\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23774_ _03087_ _03100_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__nor2_1
X_20986_ net227 _12180_ VGND VGND VPWR VPWR _12833_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25513_ _04842_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22725_ _02273_ _02274_ _01230_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26493_ clknet_leaf_86_clk_sys _00013_ net640 VGND VGND VPWR VPWR state\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_193_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25444_ _03720_ _03829_ _04131_ _04182_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22656_ _02186_ _02207_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21607_ _01165_ _01168_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__or2_1
X_25375_ _04572_ _04694_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__nor2_1
X_22587_ _02111_ _02114_ _02108_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_8_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27114_ clknet_leaf_86_clk_sys _00728_ net600 VGND VGND VPWR VPWR top0.cordic0.in_valid
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_105_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24326_ _03681_ _03682_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21538_ net126 net123 VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_35_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27045_ clknet_leaf_8_clk_sys _00662_ net592 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24257_ _03604_ _03609_ _03612_ _03614_ _03524_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__a32o_1
X_21469_ _00977_ _01008_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14010_ _05565_ _05538_ _05539_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23208_ _02659_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__buf_2
X_24188_ _03464_ _03545_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__nand2_2
XFILLER_0_120_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23139_ top0.svm0.delta\[12\] _02625_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__or2_1
X_15961_ _07913_ _07917_ _07910_ VGND VGND VPWR VPWR _08056_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_65_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17700_ net381 net358 VGND VGND VPWR VPWR _09687_ sky130_fd_sc_hd__nand2_1
X_14912_ spi0.data_packed\[63\] top0.kpq\[15\] _07075_ VGND VGND VPWR VPWR _07077_
+ sky130_fd_sc_hd__mux2_1
X_18680_ _10519_ _10534_ _10533_ VGND VGND VPWR VPWR _10658_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15892_ _07888_ _07889_ _07882_ VGND VGND VPWR VPWR _07988_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17631_ _09609_ _09611_ _09615_ _09616_ _09617_ VGND VGND VPWR VPWR _09618_ sky130_fd_sc_hd__o221a_1
X_14843_ state\[0\] _05426_ net7 VGND VGND VPWR VPWR _07040_ sky130_fd_sc_hd__a21boi_1
X_26829_ clknet_leaf_46_clk_sys _00446_ net680 VGND VGND VPWR VPWR top0.svm0.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_37_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17562_ net418 net340 VGND VGND VPWR VPWR _09549_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14774_ net26 _06824_ VGND VGND VPWR VPWR _06975_ sky130_fd_sc_hd__nand2_1
X_16513_ _08596_ _08598_ VGND VGND VPWR VPWR _08601_ sky130_fd_sc_hd__nor2_1
X_19301_ _11120_ _11241_ _11242_ VGND VGND VPWR VPWR _11243_ sky130_fd_sc_hd__and3_1
X_13725_ net50 _05894_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__nand2_1
X_17493_ _09472_ _09479_ VGND VGND VPWR VPWR _09480_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_103_clk_sys clknet_3_0__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_103_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_62_clk_sys clknet_3_4__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_62_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_16444_ _08442_ _08457_ _08456_ VGND VGND VPWR VPWR _08533_ sky130_fd_sc_hd__a21o_1
X_19232_ top0.matmul0.alpha_pass\[4\] net76 top0.matmul0.alpha_pass\[6\] _11150_ VGND
+ VGND VPWR VPWR _11180_ sky130_fd_sc_hd__or4_2
X_13656_ net54 _05520_ _05521_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19163_ _11094_ VGND VGND VPWR VPWR _11117_ sky130_fd_sc_hd__clkbuf_4
X_16375_ _08464_ VGND VGND VPWR VPWR _08465_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13587_ _05651_ _05714_ VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18114_ net338 net378 VGND VGND VPWR VPWR _10098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15326_ _07393_ _07394_ VGND VGND VPWR VPWR _07425_ sky130_fd_sc_hd__xor2_1
XFILLER_0_170_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19094_ _11047_ _10955_ _10845_ VGND VGND VPWR VPWR _11066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18045_ _09919_ _09920_ _09921_ VGND VGND VPWR VPWR _10030_ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15257_ net527 net491 VGND VGND VPWR VPWR _07356_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14208_ _06328_ _06338_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15188_ _07188_ _07189_ _07187_ VGND VGND VPWR VPWR _07287_ sky130_fd_sc_hd__o21ba_1
X_14139_ _06131_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__buf_4
XFILLER_0_123_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout409 top0.pid_d.mult0.a\[5\] VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19996_ net202 _11573_ _11510_ _11612_ _11632_ VGND VGND VPWR VPWR _11863_ sky130_fd_sc_hd__o311a_1
XFILLER_0_123_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18947_ _05449_ _10921_ VGND VGND VPWR VPWR _10922_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18878_ net308 _10775_ _10851_ _09706_ VGND VGND VPWR VPWR _10853_ sky130_fd_sc_hd__a211o_1
X_17829_ _09812_ _09815_ VGND VGND VPWR VPWR _09816_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20840_ _12066_ _12215_ _12212_ _12040_ VGND VGND VPWR VPWR _12689_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_7_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20771_ _12610_ _12619_ VGND VGND VPWR VPWR _12620_ sky130_fd_sc_hd__xnor2_2
Xfanout16 net53 VGND VGND VPWR VPWR net1027 sky130_fd_sc_hd__buf_4
XFILLER_0_58_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout27 net28 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_2
XFILLER_0_146_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22510_ net111 net107 net98 _01230_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout38 top0.periodTop_r\[11\] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
Xfanout49 top0.periodTop_r\[6\] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_4
XFILLER_0_9_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23490_ net732 top0.matmul0.cos\[0\] _02904_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22441_ _01944_ _01987_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25160_ _04436_ _04447_ _04507_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__o21a_1
X_22372_ _01909_ _01930_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24111_ _03387_ _03392_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__xor2_2
X_21323_ _12699_ _13125_ _13162_ net242 _13164_ VGND VGND VPWR VPWR _13165_ sky130_fd_sc_hd__a221o_1
X_25091_ _04438_ _04439_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24042_ _03361_ _03399_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__xnor2_4
X_21254_ _13096_ _13097_ _12940_ _12941_ _13008_ VGND VGND VPWR VPWR _13098_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_41_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20205_ _12041_ _12052_ _12053_ VGND VGND VPWR VPWR _12054_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21185_ net238 net246 VGND VGND VPWR VPWR _13029_ sky130_fd_sc_hd__and2b_1
X_20136_ net212 _11434_ _11947_ _11978_ top0.cordic0.slte0.opA\[16\] VGND VGND VPWR
+ VPWR _11992_ sky130_fd_sc_hd__a41o_1
X_25993_ top0.matmul0.beta_pass\[8\] _05169_ _05194_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__a21o_1
X_24944_ _04188_ _04191_ _04294_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__o21a_1
X_20067_ net195 _11926_ _11928_ _11810_ VGND VGND VPWR VPWR _11929_ sky130_fd_sc_hd__a22oi_1
X_24875_ _04021_ _04022_ _04023_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26614_ clknet_leaf_30_clk_sys _00231_ net623 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_23826_ _02983_ _03182_ _03183_ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_197_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26545_ clknet_leaf_49_clk_sys _00168_ net675 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23757_ _03112_ _03114_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__nor2_2
XFILLER_0_71_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20969_ _12698_ _12815_ net241 VGND VGND VPWR VPWR _12816_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_68_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13510_ _05616_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_166_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22708_ _02186_ _02207_ _02224_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__or3_1
X_14490_ _06693_ _06694_ _06696_ VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__o21ai_4
X_26476_ clknet_leaf_11_clk_sys _00107_ net603 VGND VGND VPWR VPWR top0.periodTop\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_23688_ _03023_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25427_ _04745_ _04769_ _04694_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__mux2_1
X_13441_ _05548_ _05555_ _05553_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_48_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22639_ _11674_ net93 _01115_ _02188_ _02191_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__o311a_2
XFILLER_0_180_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16160_ _08227_ _08225_ VGND VGND VPWR VPWR _08252_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25358_ _04382_ _04647_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__or2_1
XFILLER_0_180_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13372_ _05531_ _05532_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__nor2_2
XFILLER_0_23_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15111_ _07201_ _07209_ VGND VGND VPWR VPWR _07210_ sky130_fd_sc_hd__xnor2_2
X_24309_ _03225_ _03226_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16091_ _08108_ _08119_ _08183_ VGND VGND VPWR VPWR _08184_ sky130_fd_sc_hd__o21a_1
X_25289_ _04628_ _04634_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__and2b_1
X_27028_ clknet_leaf_18_clk_sys _00645_ net614 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_15042_ top0.pid_d.prev_int\[12\] _07139_ _07143_ net978 VGND VGND VPWR VPWR _00129_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19850_ _11726_ VGND VGND VPWR VPWR _11727_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18801_ _10775_ _10776_ VGND VGND VPWR VPWR _10777_ sky130_fd_sc_hd__xor2_2
X_19781_ _11513_ _11662_ VGND VGND VPWR VPWR _11663_ sky130_fd_sc_hd__nand2_1
X_16993_ top0.pid_q.prev_error\[11\] top0.pid_q.curr_error\[11\] VGND VGND VPWR VPWR
+ _09048_ sky130_fd_sc_hd__nand2_1
X_18732_ _10636_ _10638_ _10708_ VGND VGND VPWR VPWR _10709_ sky130_fd_sc_hd__a21bo_1
X_15944_ _08012_ _08038_ VGND VGND VPWR VPWR _08039_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_183_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18663_ _10635_ _10640_ VGND VGND VPWR VPWR _10641_ sky130_fd_sc_hd__xnor2_1
X_15875_ _07821_ _07822_ _07820_ VGND VGND VPWR VPWR _07971_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_153_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14826_ _07021_ _07024_ VGND VGND VPWR VPWR _07026_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17614_ _09563_ _09566_ _09600_ VGND VGND VPWR VPWR _09601_ sky130_fd_sc_hd__a21o_1
XFILLER_0_192_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18594_ _10559_ _10572_ VGND VGND VPWR VPWR _10573_ sky130_fd_sc_hd__xor2_4
XFILLER_0_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14757_ _06958_ _05629_ net20 VGND VGND VPWR VPWR _06959_ sky130_fd_sc_hd__or3b_1
X_17545_ net407 _09531_ _09460_ VGND VGND VPWR VPWR _09532_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13708_ _05913_ _05918_ _05920_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__a21o_1
X_17476_ net395 _09431_ _09433_ VGND VGND VPWR VPWR _09463_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14688_ _06888_ _06891_ VGND VGND VPWR VPWR _06892_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19215_ top0.pid_d.curr_error\[4\] VGND VGND VPWR VPWR _11164_ sky130_fd_sc_hd__inv_2
X_13639_ _05828_ _05851_ _05849_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__o21a_1
X_16427_ _08430_ _08432_ _08431_ VGND VGND VPWR VPWR _08516_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16358_ net476 net473 VGND VGND VPWR VPWR _08448_ sky130_fd_sc_hd__or2b_1
X_19146_ net397 _11096_ _11108_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15309_ net542 net471 _07407_ VGND VGND VPWR VPWR _07408_ sky130_fd_sc_hd__and3_1
XFILLER_0_140_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16289_ _08377_ _08379_ VGND VGND VPWR VPWR _08380_ sky130_fd_sc_hd__xnor2_1
X_19077_ _10955_ _11012_ _10845_ VGND VGND VPWR VPWR _11049_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18028_ net307 _10012_ VGND VGND VPWR VPWR _10013_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_160_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout206 top0.state\[2\] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
Xfanout217 net220 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout228 top0.cordic0.vec\[0\]\[15\] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__buf_2
Xfanout239 net240 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19979_ net183 _11573_ _11509_ _11810_ VGND VGND VPWR VPWR _11847_ sky130_fd_sc_hd__or4b_1
XFILLER_0_201_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22990_ top0.svm0.delta\[9\] VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__inv_2
XFILLER_0_198_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21941_ net159 net136 _01136_ _01301_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__o31a_1
XFILLER_0_55_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24660_ _03207_ _03208_ _03196_ _03197_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__o22a_1
X_21872_ _01424_ _01433_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23611_ _02972_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__clkbuf_1
X_20823_ _12670_ _12400_ _12671_ _12399_ _12408_ VGND VGND VPWR VPWR _12672_ sky130_fd_sc_hd__a221o_1
X_24591_ _03934_ _03945_ VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_148_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26330_ spi0.data_packed\[63\] spi0.data_packed\[64\] net695 VGND VGND VPWR VPWR
+ _05397_ sky130_fd_sc_hd__mux2_1
X_23542_ _05460_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20754_ _12602_ _12598_ _11593_ net258 VGND VGND VPWR VPWR _12603_ sky130_fd_sc_hd__a211o_1
XFILLER_0_148_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26261_ _05362_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23473_ net1005 top0.matmul0.sin\[6\] _05461_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__mux2_1
X_20685_ _12261_ _12357_ VGND VGND VPWR VPWR _12534_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25212_ _03254_ _04174_ _03325_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22424_ _01980_ _01981_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__or2_2
X_26192_ spi0.data_packed\[12\] _05325_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25143_ _04427_ _04432_ _04424_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_165_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22355_ _01225_ _01327_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21306_ _13014_ _13144_ _13148_ VGND VGND VPWR VPWR _13149_ sky130_fd_sc_hd__a21oi_1
X_25074_ _04421_ _04422_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22286_ net101 net96 VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__and2_1
XFILLER_0_198_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_2_clk_sys clknet_3_2__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_2_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_10_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_10_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_24025_ _03380_ _03381_ _03382_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__a21o_2
Xhold260 top0.currT_r\[6\] VGND VGND VPWR VPWR net960 sky130_fd_sc_hd__dlygate4sd3_1
X_21237_ _12610_ _12628_ VGND VGND VPWR VPWR _13081_ sky130_fd_sc_hd__or2b_1
Xhold271 top0.pid_d.prev_int\[2\] VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 top0.pid_q.prev_int\[4\] VGND VGND VPWR VPWR net982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 top0.matmul0.matmul_stage_inst.a\[0\] VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__dlygate4sd3_1
X_21168_ _13010_ _13012_ VGND VGND VPWR VPWR _13013_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20119_ net177 top0.cordic0.slte0.opA\[15\] VGND VGND VPWR VPWR _11976_ sky130_fd_sc_hd__nand2_1
X_13990_ _06198_ _06202_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__xnor2_2
X_21099_ _12746_ _12943_ VGND VGND VPWR VPWR _12945_ sky130_fd_sc_hd__nor2_1
X_25976_ top0.pid_q.out\[4\] _12032_ _05014_ spi0.data_packed\[52\] VGND VGND VPWR
+ VPWR _05182_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24927_ _04180_ _04181_ _04277_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_172_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15660_ _07754_ _07757_ VGND VGND VPWR VPWR _07758_ sky130_fd_sc_hd__xnor2_1
X_24858_ _04203_ _04209_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_197_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14611_ _06792_ _06808_ _06812_ _06815_ VGND VGND VPWR VPWR _06816_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_158_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23809_ _03154_ _03166_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__xor2_1
X_15591_ _07610_ _07689_ _07220_ _07298_ VGND VGND VPWR VPWR _07690_ sky130_fd_sc_hd__a2bb2o_1
X_24789_ _04038_ _04045_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__nand2_2
XFILLER_0_96_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17330_ top0.matmul0.beta_pass\[12\] _09320_ net562 VGND VGND VPWR VPWR _09321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14542_ net861 _06280_ _06748_ _06381_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__a22o_1
X_26528_ clknet_leaf_61_clk_sys _00151_ net651 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_166_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17261_ top0.matmul0.beta_pass\[2\] _09261_ net563 VGND VGND VPWR VPWR _09262_ sky130_fd_sc_hd__mux2_1
X_14473_ _06608_ _06673_ _06675_ _06609_ _06680_ VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__a221o_2
X_26459_ clknet_leaf_91_clk_sys net692 net600 VGND VGND VPWR VPWR spi0.cs_sync\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_166_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16212_ _08283_ _08303_ VGND VGND VPWR VPWR _08304_ sky130_fd_sc_hd__xnor2_2
X_19000_ _10973_ VGND VGND VPWR VPWR _10974_ sky130_fd_sc_hd__inv_2
XFILLER_0_180_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13424_ top0.matmul0.alpha_pass\[9\] _05466_ _05467_ VGND VGND VPWR VPWR _05637_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_153_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17192_ _09201_ _09195_ _08404_ VGND VGND VPWR VPWR _09202_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16143_ _07701_ _08235_ VGND VGND VPWR VPWR _08236_ sky130_fd_sc_hd__nor2_1
X_13355_ _05565_ _05567_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16074_ _08124_ _08125_ _08166_ VGND VGND VPWR VPWR _08167_ sky130_fd_sc_hd__a21bo_1
X_13286_ _05487_ _05492_ _05498_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19902_ net181 _11775_ VGND VGND VPWR VPWR _11776_ sky130_fd_sc_hd__or2_1
X_15025_ _07139_ VGND VGND VPWR VPWR _07140_ sky130_fd_sc_hd__clkbuf_4
X_19833_ net244 _11705_ VGND VGND VPWR VPWR _11711_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19764_ net266 _11435_ VGND VGND VPWR VPWR _11647_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16976_ net429 _09030_ _09031_ _09011_ VGND VGND VPWR VPWR _09032_ sky130_fd_sc_hd__o2bb2a_1
X_18715_ net374 net365 _10689_ _10691_ VGND VGND VPWR VPWR _10692_ sky130_fd_sc_hd__a31o_1
X_15927_ net532 net446 VGND VGND VPWR VPWR _08022_ sky130_fd_sc_hd__nand2_1
X_19695_ _11425_ _11577_ _11579_ _11580_ net82 VGND VGND VPWR VPWR _11581_ sky130_fd_sc_hd__a32o_2
XFILLER_0_189_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18646_ _10622_ _10623_ net364 VGND VGND VPWR VPWR _10624_ sky130_fd_sc_hd__o21ai_1
X_15858_ _07833_ _07835_ _07953_ VGND VGND VPWR VPWR _07954_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_143_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14809_ _06972_ VGND VGND VPWR VPWR _07009_ sky130_fd_sc_hd__inv_2
X_18577_ _10481_ _10485_ _10480_ VGND VGND VPWR VPWR _10556_ sky130_fd_sc_hd__a21o_1
X_15789_ net508 _07767_ _07883_ _07885_ VGND VGND VPWR VPWR _07886_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17528_ _09456_ _09514_ VGND VGND VPWR VPWR _09515_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17459_ _09427_ _09445_ VGND VGND VPWR VPWR _09446_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20470_ _11726_ _12246_ _12318_ VGND VGND VPWR VPWR _12319_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_104_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19129_ top0.pid_d.state\[3\] _05442_ _11094_ VGND VGND VPWR VPWR _11099_ sky130_fd_sc_hd__and3_2
XFILLER_0_113_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22140_ _01311_ _01076_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22071_ _01588_ _01568_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_61_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21022_ _12785_ VGND VGND VPWR VPWR _12869_ sky130_fd_sc_hd__inv_2
XFILLER_0_195_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25830_ top0.matmul0.alpha_pass\[4\] top0.matmul0.beta_pass\[4\] VGND VGND VPWR VPWR
+ _05054_ sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_113_Left_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25761_ _05001_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22973_ _02440_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__clkbuf_4
X_24712_ _04049_ _04056_ _04053_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_93_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21924_ _01281_ _01484_ _01485_ _01442_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__a22o_1
X_25692_ _04886_ top0.matmul0.sin\[13\] net73 VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_195_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_182_Right_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24643_ _02979_ _02980_ _03061_ _03062_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__o22a_1
X_21855_ net158 _01178_ _01414_ _01416_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__a31o_1
XFILLER_0_171_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20806_ _12651_ _12652_ _12653_ _12654_ VGND VGND VPWR VPWR _12655_ sky130_fd_sc_hd__o22ai_1
X_24574_ _03783_ _03814_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21786_ _01347_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26313_ _05388_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23525_ _02928_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_122_Left_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20737_ _12348_ _12584_ _12551_ VGND VGND VPWR VPWR _12586_ sky130_fd_sc_hd__mux2_1
X_27293_ clknet_3_0__leaf_clk_mosi _00907_ VGND VGND VPWR VPWR spi0.data_packed\[79\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26244_ spi0.data_packed\[20\] spi0.data_packed\[21\] net698 VGND VGND VPWR VPWR
+ _05354_ sky130_fd_sc_hd__mux2_1
X_23456_ _02885_ _02886_ _02888_ _02890_ VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__a211o_1
X_20668_ _12471_ _12482_ _12477_ VGND VGND VPWR VPWR _12517_ sky130_fd_sc_hd__or3b_1
XFILLER_0_34_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22407_ _01408_ _01964_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__xnor2_1
X_26175_ _05312_ top0.cordic0.slte0.opB\[10\] _12006_ VGND VGND VPWR VPWR _05313_
+ sky130_fd_sc_hd__mux2_1
X_23387_ _02809_ _02818_ net116 VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__o21a_1
X_20599_ _11408_ _12059_ _12333_ VGND VGND VPWR VPWR _12448_ sky130_fd_sc_hd__a21oi_1
X_25126_ _04461_ _04472_ _04473_ _04386_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_104_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22338_ _01863_ _01865_ _01861_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25057_ _04306_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__buf_4
XFILLER_0_103_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22269_ _01824_ _01828_ _01819_ VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__a21oi_1
X_24008_ _03363_ _03324_ _03056_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_131_Left_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16830_ top0.pid_q.prev_error\[1\] top0.pid_q.curr_error\[1\] VGND VGND VPWR VPWR
+ _08896_ sky130_fd_sc_hd__xor2_1
Xfanout570 top0.matmul0.matmul_stage_inst.state\[2\] VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__buf_4
Xfanout581 net585 VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__clkbuf_2
Xfanout592 net597 VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__clkbuf_4
X_13973_ _06182_ _06185_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__xnor2_2
X_16761_ top0.pid_q.out\[14\] top0.pid_q.curr_int\[14\] VGND VGND VPWR VPWR _08845_
+ sky130_fd_sc_hd__nor2_1
X_25959_ _05168_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__buf_2
X_18500_ _10469_ _10479_ VGND VGND VPWR VPWR _10480_ sky130_fd_sc_hd__xnor2_1
X_15712_ _07695_ _07808_ _07694_ VGND VGND VPWR VPWR _07809_ sky130_fd_sc_hd__o21bai_1
X_16692_ _08757_ _08776_ VGND VGND VPWR VPWR _08777_ sky130_fd_sc_hd__or2_1
X_19480_ _10828_ _10923_ _10924_ VGND VGND VPWR VPWR _11374_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18431_ _10314_ VGND VGND VPWR VPWR _10412_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15643_ net460 net525 VGND VGND VPWR VPWR _07741_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18362_ _10165_ _10251_ _10326_ _10329_ _10250_ VGND VGND VPWR VPWR _10343_ sky130_fd_sc_hd__o221a_1
X_15574_ _07564_ _07672_ _07581_ VGND VGND VPWR VPWR _07673_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_140_Left_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14525_ net45 _06351_ _06730_ _06731_ VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__a31o_1
X_17313_ _09304_ _09300_ _09305_ VGND VGND VPWR VPWR _09306_ sky130_fd_sc_hd__a21o_1
XFILLER_0_166_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18293_ _10271_ _10274_ VGND VGND VPWR VPWR _10275_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14456_ _06597_ _06600_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__nor2_1
X_17244_ _09246_ _09247_ VGND VGND VPWR VPWR _09248_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13407_ net64 _05602_ _05603_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17175_ top0.pid_q.curr_int\[6\] _09184_ _09186_ VGND VGND VPWR VPWR _09187_ sky130_fd_sc_hd__o21ai_2
X_14387_ _06489_ _06490_ _06595_ VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16126_ _08092_ _08135_ _08218_ VGND VGND VPWR VPWR _08219_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13338_ _05538_ _05539_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__nor2_2
XFILLER_0_40_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16057_ _08001_ _08007_ _08150_ VGND VGND VPWR VPWR _08151_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13269_ _05473_ _05481_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15008_ _07129_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19816_ _11684_ _11690_ _11694_ VGND VGND VPWR VPWR _11696_ sky130_fd_sc_hd__or3_1
X_19747_ _11573_ _11629_ _11576_ VGND VGND VPWR VPWR _11630_ sky130_fd_sc_hd__a21oi_1
X_16959_ _09014_ _09015_ net547 VGND VGND VPWR VPWR _09016_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19678_ net182 _11559_ _11564_ VGND VGND VPWR VPWR _11565_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_154_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18629_ _10573_ _10577_ _10575_ VGND VGND VPWR VPWR _10607_ sky130_fd_sc_hd__o21a_1
XFILLER_0_52_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21640_ _01078_ _01199_ _01198_ net144 _01201_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21571_ net120 net114 VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__nor2_1
XANTENNA_11 net1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_23310_ net140 _02744_ _02707_ net144 _02719_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__o2111a_1
XANTENNA_33 _05500_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20522_ _11758_ _12075_ VGND VGND VPWR VPWR _12371_ sky130_fd_sc_hd__xnor2_4
XANTENNA_44 net1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24290_ _03624_ _03625_ _03635_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23241_ _02687_ _02688_ _02689_ _02690_ _11572_ _11420_ VGND VGND VPWR VPWR _02691_
+ sky130_fd_sc_hd__mux4_1
X_20453_ net294 net274 VGND VGND VPWR VPWR _12302_ sky130_fd_sc_hd__or2b_1
XFILLER_0_162_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23172_ _05717_ _06945_ _02644_ net781 VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__a22o_1
X_20384_ _12125_ _12231_ _12232_ VGND VGND VPWR VPWR _12233_ sky130_fd_sc_hd__o21a_1
XFILLER_0_179_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22123_ net78 net99 net86 VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22054_ net119 net105 VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__nand2_2
X_26931_ clknet_leaf_7_clk_sys _00548_ net592 VGND VGND VPWR VPWR top0.matmul0.cos\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21005_ net225 net221 _12696_ net234 VGND VGND VPWR VPWR _12852_ sky130_fd_sc_hd__a211o_1
X_26862_ clknet_leaf_40_clk_sys _00479_ net682 VGND VGND VPWR VPWR top0.svm0.tA\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_25813_ top0.matmul0.alpha_pass\[2\] top0.matmul0.beta_pass\[2\] VGND VGND VPWR VPWR
+ _05039_ sky130_fd_sc_hd__xnor2_2
X_26793_ clknet_leaf_109_clk_sys _00410_ net578 VGND VGND VPWR VPWR top0.cordic0.sin\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25744_ net993 _04882_ _05458_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__mux2_1
Xmax_cap13 _07699_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
X_22956_ _02458_ _02461_ _02467_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__a21o_1
X_21907_ _01358_ _01436_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__nand2_1
X_25675_ net805 _04904_ _04946_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_70_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22887_ top0.svm0.tB\[14\] _02404_ _02405_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__o21a_1
XFILLER_0_167_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24626_ _03975_ _03976_ _03978_ _03742_ _03979_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__o221ai_4
X_21838_ _01398_ _01399_ _01390_ _01391_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__o211a_1
XFILLER_0_183_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24557_ _03910_ _03911_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21769_ net135 _01327_ _01329_ _01330_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__a211o_2
XFILLER_0_194_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14310_ _06518_ _06519_ VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23508_ _02919_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27276_ clknet_3_7__leaf_clk_mosi _00890_ VGND VGND VPWR VPWR spi0.data_packed\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_15290_ _07321_ _07382_ _07384_ net525 _07388_ VGND VGND VPWR VPWR _07389_ sky130_fd_sc_hd__a221o_1
X_24488_ _03738_ _03745_ _03843_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14241_ _06296_ _06297_ _06298_ _06299_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26227_ _05345_ VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__clkbuf_1
X_23439_ _02875_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14172_ _06373_ _06377_ _06370_ VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__mux2_1
X_26158_ spi0.data_packed\[3\] spi0.data_packed\[4\] _05292_ VGND VGND VPWR VPWR _05299_
+ sky130_fd_sc_hd__and3_1
X_25109_ _04336_ _04344_ _04345_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_21_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26089_ top0.matmul0.alpha_pass\[14\] _05168_ _05268_ VGND VGND VPWR VPWR _05269_
+ sky130_fd_sc_hd__a21o_1
X_18980_ _10950_ _10953_ VGND VGND VPWR VPWR _10954_ sky130_fd_sc_hd__xnor2_2
X_17931_ _09833_ _09838_ _09831_ VGND VGND VPWR VPWR _09917_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_84_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17862_ net389 net346 net384 net351 VGND VGND VPWR VPWR _09849_ sky130_fd_sc_hd__nand4_1
XFILLER_0_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19601_ _11485_ top0.cordic0.slte0.opA\[8\] _11488_ _11489_ VGND VGND VPWR VPWR _11490_
+ sky130_fd_sc_hd__a22o_1
X_16813_ _07698_ _08853_ VGND VGND VPWR VPWR _08880_ sky130_fd_sc_hd__or2_1
X_17793_ _09776_ _09779_ VGND VGND VPWR VPWR _09780_ sky130_fd_sc_hd__xnor2_1
X_19532_ net179 VGND VGND VPWR VPWR _11422_ sky130_fd_sc_hd__inv_2
X_16744_ net500 _08825_ _08827_ net444 VGND VGND VPWR VPWR _08828_ sky130_fd_sc_hd__a22o_1
X_13956_ _06162_ _06166_ _06167_ _06168_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_199_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_191_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19463_ _11357_ _11353_ _11358_ VGND VGND VPWR VPWR _11359_ sky130_fd_sc_hd__o21a_1
X_13887_ _06092_ _06093_ _06099_ VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__a21oi_2
X_16675_ net504 net445 VGND VGND VPWR VPWR _08760_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18414_ _10287_ VGND VGND VPWR VPWR _10395_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15626_ _07624_ _07625_ _07626_ VGND VGND VPWR VPWR _07724_ sky130_fd_sc_hd__o21ai_1
X_19394_ _11297_ _11298_ VGND VGND VPWR VPWR _11299_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18345_ _10238_ _10239_ _10236_ VGND VGND VPWR VPWR _10327_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_167_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15557_ _07648_ _07655_ VGND VGND VPWR VPWR _07656_ sky130_fd_sc_hd__nor2_1
XFILLER_0_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14508_ _05579_ _06640_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__nand2_1
X_18276_ net397 net366 _10257_ _09399_ _09363_ VGND VGND VPWR VPWR _10258_ sky130_fd_sc_hd__a32o_1
X_15488_ _07585_ _07546_ _07547_ VGND VGND VPWR VPWR _07587_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17227_ _09231_ _09232_ VGND VGND VPWR VPWR _09233_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14439_ _06643_ _06646_ VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_181_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17158_ top0.pid_q.prev_int\[4\] _09165_ _09171_ VGND VGND VPWR VPWR _09172_ sky130_fd_sc_hd__o21a_2
X_16109_ net466 net507 VGND VGND VPWR VPWR _08202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17089_ top0.pid_q.curr_error\[3\] _00011_ _09117_ VGND VGND VPWR VPWR _09121_ sky130_fd_sc_hd__and3_1
XFILLER_0_161_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_57_clk_sys clknet_3_4__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_57_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22810_ top0.svm0.counter\[5\] _02323_ _02327_ _02328_ _02329_ VGND VGND VPWR VPWR
+ _02330_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23790_ _03147_ VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__buf_4
XFILLER_0_196_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22741_ net174 net197 VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25460_ _04742_ _04739_ _04745_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__nor3_1
XFILLER_0_149_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22672_ _02206_ _02223_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__xnor2_2
X_24411_ _03007_ _02982_ _03764_ _03766_ VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__o31a_1
X_21623_ net154 _01151_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__xor2_1
X_25391_ _03123_ _04676_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27130_ clknet_leaf_33_clk_sys _00744_ net665 VGND VGND VPWR VPWR top0.c_out_calc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24342_ _03697_ _03695_ _03696_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__and3b_1
XFILLER_0_173_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21554_ net114 net109 VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27061_ clknet_leaf_21_clk_sys _00678_ net610 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.a\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_20505_ net274 _12353_ VGND VGND VPWR VPWR _12354_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24273_ _03620_ _03622_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__or2_1
X_21485_ _12180_ _12824_ _01046_ _01048_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__o31a_1
XFILLER_0_172_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26012_ top0.pid_q.out\[12\] _05198_ _05199_ spi0.data_packed\[60\] VGND VGND VPWR
+ VPWR _05210_ sky130_fd_sc_hd__a22o_1
X_23224_ net160 _11784_ _02673_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__or3_1
XFILLER_0_200_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20436_ _11407_ net299 VGND VGND VPWR VPWR _12285_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23155_ _02639_ _02640_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20367_ _12214_ _12215_ VGND VGND VPWR VPWR _12216_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22106_ _01662_ _01665_ _01667_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__mux2_1
X_23086_ _02576_ _02579_ _02584_ _02585_ _02586_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__a221o_1
X_20298_ _12139_ _12141_ _12145_ VGND VGND VPWR VPWR _12147_ sky130_fd_sc_hd__nand3_1
XFILLER_0_101_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22037_ _01595_ _01597_ _01598_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26914_ clknet_leaf_1_clk_sys _00531_ net582 VGND VGND VPWR VPWR top0.matmul0.sin\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26845_ clknet_leaf_44_clk_sys _00462_ net681 VGND VGND VPWR VPWR top0.svm0.delta\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_13810_ _05523_ _05524_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__and2_1
X_14790_ _06949_ _06990_ VGND VGND VPWR VPWR _06991_ sky130_fd_sc_hd__or2_1
XFILLER_0_202_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23988_ net1017 _03161_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__nor2_1
X_26776_ clknet_leaf_5_clk_sys _00393_ net590 VGND VGND VPWR VPWR top0.cordic0.cos\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13741_ _05950_ _05951_ _05952_ _05953_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__o22a_1
X_22939_ _02447_ _02452_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__nand2_1
X_25727_ net906 _04964_ _04913_ _04982_ VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13672_ _05837_ _05842_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__xnor2_1
X_16460_ _08547_ _08548_ VGND VGND VPWR VPWR _08549_ sky130_fd_sc_hd__or2b_1
XFILLER_0_167_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25658_ _04931_ _04932_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15411_ _07479_ _07502_ _07509_ VGND VGND VPWR VPWR _07510_ sky130_fd_sc_hd__o21a_1
X_24609_ _03863_ _03957_ _03962_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16391_ top0.pid_q.out\[9\] _08480_ net13 VGND VGND VPWR VPWR _08481_ sky130_fd_sc_hd__mux2_1
X_25589_ net73 VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18130_ _10015_ _10020_ _10113_ VGND VGND VPWR VPWR _10114_ sky130_fd_sc_hd__a21o_1
X_15342_ net542 net475 VGND VGND VPWR VPWR _07441_ sky130_fd_sc_hd__nand2_1
XFILLER_0_171_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18061_ net424 net310 VGND VGND VPWR VPWR _10046_ sky130_fd_sc_hd__nand2_1
X_15273_ net527 net524 net495 net491 VGND VGND VPWR VPWR _07372_ sky130_fd_sc_hd__and4_1
XFILLER_0_81_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27259_ clknet_3_3__leaf_clk_mosi _00873_ VGND VGND VPWR VPWR spi0.data_packed\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14224_ net30 net1015 VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__nand2_2
XFILLER_0_151_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17012_ _05662_ net428 top0.currT_r\[13\] _05437_ VGND VGND VPWR VPWR _09065_ sky130_fd_sc_hd__and4_1
XFILLER_0_34_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14155_ _06239_ _06252_ _06366_ VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14086_ _06189_ _06196_ _06186_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__a21oi_1
X_18963_ _10633_ _10936_ VGND VGND VPWR VPWR _10937_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17914_ top0.pid_d.out\[0\] top0.pid_d.curr_int\[0\] _09899_ VGND VGND VPWR VPWR
+ _09900_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18894_ _10867_ _10868_ VGND VGND VPWR VPWR _10869_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17845_ _09783_ _09784_ _09666_ VGND VGND VPWR VPWR _09832_ sky130_fd_sc_hd__o21bai_1
X_17776_ _09636_ _09762_ _09637_ VGND VGND VPWR VPWR _09763_ sky130_fd_sc_hd__o21a_1
XFILLER_0_156_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14988_ spi0.data_packed\[0\] top0.periodTop\[0\] _07108_ VGND VGND VPWR VPWR _07119_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19515_ top0.pid_d.curr_int\[15\] _11289_ _11341_ _11405_ VGND VGND VPWR VPWR _11406_
+ sky130_fd_sc_hd__a22o_1
X_16727_ _08809_ _08810_ VGND VGND VPWR VPWR _08811_ sky130_fd_sc_hd__nor2_1
X_13939_ _06146_ _06151_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19446_ _11342_ _11336_ VGND VGND VPWR VPWR _11344_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16658_ net549 _07700_ _08738_ _08743_ VGND VGND VPWR VPWR _08744_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_186_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15609_ _07707_ _07706_ top0.pid_q.out\[0\] VGND VGND VPWR VPWR _07708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19377_ net874 _11284_ _11287_ top0.pid_d.curr_error\[10\] VGND VGND VPWR VPWR _00320_
+ sky130_fd_sc_hd__a22o_1
X_16589_ _08673_ _08674_ _08675_ VGND VGND VPWR VPWR _08676_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18328_ _10103_ _10309_ VGND VGND VPWR VPWR _10310_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18259_ _10167_ _10241_ VGND VGND VPWR VPWR _10242_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21270_ net239 _13028_ VGND VGND VPWR VPWR _13113_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20221_ _12054_ _12055_ _12060_ _12069_ VGND VGND VPWR VPWR _12070_ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20152_ _12005_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__clkbuf_1
X_24960_ _04307_ _04231_ _04258_ _04310_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__o211a_1
X_20083_ _11942_ _11943_ VGND VGND VPWR VPWR _11944_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23911_ _03267_ _03268_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__nand2_2
XFILLER_0_58_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24891_ _04158_ _04242_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__xnor2_1
X_23842_ _03107_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__buf_4
X_26630_ clknet_leaf_74_clk_sys _00247_ net655 VGND VGND VPWR VPWR top0.pid_d.out\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_23773_ _03101_ _03111_ _03130_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__a21oi_2
X_26561_ clknet_leaf_51_clk_sys _00184_ net671 VGND VGND VPWR VPWR top0.pid_q.curr_error\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_68_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20985_ _11757_ net221 VGND VGND VPWR VPWR _12832_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25512_ top0.matmul0.matmul_stage_inst.mult1\[12\] _04659_ _03148_ VGND VGND VPWR
+ VPWR _04842_ sky130_fd_sc_hd__mux2_1
X_22724_ _01248_ _02112_ _02023_ _01948_ VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__o22a_1
X_26492_ clknet_leaf_85_clk_sys _00012_ net640 VGND VGND VPWR VPWR state\[0\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_48_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25443_ _04406_ _04785_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22655_ _02186_ _02207_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__or2_1
XFILLER_0_192_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21606_ net110 _01163_ _01167_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__and3_1
X_25374_ _04572_ _04694_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__and2_1
X_22586_ _02101_ _02116_ _02139_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__o21a_2
XFILLER_0_36_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24325_ _02994_ _02996_ _02979_ _02980_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27113_ clknet_leaf_89_clk_sys _00727_ net603 VGND VGND VPWR VPWR top0.matmul0.start
+ sky130_fd_sc_hd__dfrtp_2
X_21537_ net164 _01095_ _01097_ _01098_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27044_ clknet_leaf_16_clk_sys _00661_ net613 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_24256_ _03533_ _03613_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__xnor2_1
X_21468_ _01028_ _01029_ _01032_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_160_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23207_ _02656_ _02658_ net179 VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20419_ _11653_ _12267_ _12144_ VGND VGND VPWR VPWR _12268_ sky130_fd_sc_hd__o21bai_1
X_24187_ _03541_ _03544_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__xnor2_2
X_21399_ _00932_ _00951_ _00965_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__o21ai_4
X_23138_ net972 _02626_ _02627_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23069_ net170 _02564_ _02540_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__or3b_1
X_15960_ _07954_ _07956_ _08054_ VGND VGND VPWR VPWR _08055_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14911_ _07076_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__clkbuf_1
X_15891_ _07979_ _07986_ VGND VGND VPWR VPWR _07987_ sky130_fd_sc_hd__xnor2_1
X_17630_ net426 _09612_ _09609_ VGND VGND VPWR VPWR _09617_ sky130_fd_sc_hd__or3b_1
X_26828_ clknet_leaf_46_clk_sys _00445_ net680 VGND VGND VPWR VPWR top0.svm0.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14842_ state\[0\] _05425_ _05422_ VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_188_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17561_ _09544_ _09546_ _09535_ VGND VGND VPWR VPWR _09548_ sky130_fd_sc_hd__a21o_1
X_14773_ _06954_ _06955_ _06973_ VGND VGND VPWR VPWR _06974_ sky130_fd_sc_hd__o21a_1
X_26759_ clknet_leaf_94_clk_sys _00376_ net590 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_19300_ top0.matmul0.alpha_pass\[11\] _11221_ top0.matmul0.alpha_pass\[12\] VGND
+ VGND VPWR VPWR _11242_ sky130_fd_sc_hd__o21ai_1
X_16512_ _08599_ VGND VGND VPWR VPWR _08600_ sky130_fd_sc_hd__inv_2
X_13724_ net1027 _05496_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__nand2_1
X_17492_ _09475_ _09478_ VGND VGND VPWR VPWR _09479_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19231_ net440 _11177_ _11178_ VGND VGND VPWR VPWR _11179_ sky130_fd_sc_hd__and3_1
X_16443_ _08521_ _08531_ VGND VGND VPWR VPWR _08532_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_195_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13655_ net67 _05551_ _05866_ _05867_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__a31o_1
XFILLER_0_186_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19162_ net365 _11095_ _11116_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__a21o_1
X_13586_ _05716_ _05798_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__or2_1
X_16374_ _08459_ _08462_ VGND VGND VPWR VPWR _08464_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18113_ _10024_ _10035_ _10096_ VGND VGND VPWR VPWR _10097_ sky130_fd_sc_hd__o21a_1
X_15325_ _07418_ _07423_ VGND VGND VPWR VPWR _07424_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19093_ net363 _11064_ VGND VGND VPWR VPWR _11065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18044_ _10025_ _10028_ VGND VGND VPWR VPWR _10029_ sky130_fd_sc_hd__xnor2_2
X_15256_ net542 net539 net471 net475 VGND VGND VPWR VPWR _07355_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14207_ _06415_ _06416_ _06408_ VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15187_ _07282_ _07285_ VGND VGND VPWR VPWR _07286_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_105_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14138_ _06191_ _06193_ _06131_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__o21a_1
X_19995_ net202 net190 _11510_ VGND VGND VPWR VPWR _11862_ sky130_fd_sc_hd__or3_1
XFILLER_0_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14069_ net56 _05721_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__nand2_2
X_18946_ top0.pid_d.out\[12\] _10920_ _07141_ VGND VGND VPWR VPWR _10921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18877_ _10494_ _10851_ VGND VGND VPWR VPWR _10852_ sky130_fd_sc_hd__xnor2_1
X_17828_ _09644_ _09813_ _09814_ VGND VGND VPWR VPWR _09815_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17759_ _09516_ _09517_ _09603_ _09745_ VGND VGND VPWR VPWR _09746_ sky130_fd_sc_hd__a211o_1
XFILLER_0_178_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20770_ _12609_ _12616_ VGND VGND VPWR VPWR _12619_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_187_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout17 net519 VGND VGND VPWR VPWR net1028 sky130_fd_sc_hd__buf_4
X_19429_ top0.pid_d.prev_int\[5\] _11325_ top0.pid_d.curr_int\[5\] VGND VGND VPWR
+ VPWR _11329_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout28 net1030 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_4
Xfanout39 net40 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22440_ net727 _12004_ _12740_ _01997_ VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__a31o_1
XFILLER_0_73_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22371_ _01916_ _01929_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24110_ _03461_ _03462_ _03465_ _03466_ _03467_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__a32o_2
X_21322_ _13122_ _13163_ _13125_ VGND VGND VPWR VPWR _13164_ sky130_fd_sc_hd__o21ba_1
X_25090_ _03254_ _03743_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24041_ _03353_ _03358_ VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__xnor2_2
X_21253_ _12244_ _12673_ _12807_ _12736_ VGND VGND VPWR VPWR _13097_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_64_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20204_ _12044_ _12046_ _12051_ VGND VGND VPWR VPWR _12053_ sky130_fd_sc_hd__a21oi_1
X_21184_ net221 _12761_ VGND VGND VPWR VPWR _13028_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_187_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20135_ _11984_ _11985_ _11988_ net212 _11990_ VGND VGND VPWR VPWR _11991_ sky130_fd_sc_hd__o221a_1
X_25992_ top0.pid_q.out\[8\] _12032_ _05014_ spi0.data_packed\[56\] VGND VGND VPWR
+ VPWR _05194_ sky130_fd_sc_hd__a22o_1
X_24943_ _04188_ _04191_ _04189_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__a21o_1
X_20066_ _11654_ _11513_ _11927_ VGND VGND VPWR VPWR _11928_ sky130_fd_sc_hd__a21o_1
X_24874_ _04222_ _04225_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_197_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26613_ clknet_leaf_30_clk_sys _00230_ net623 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_197_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23825_ _02992_ _03001_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__nor2_1
XFILLER_0_200_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23756_ _03113_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__buf_4
X_26544_ clknet_leaf_51_clk_sys _00167_ net661 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20968_ _11726_ _11739_ VGND VGND VPWR VPWR _12815_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22707_ _02231_ _02224_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__nand2_1
X_23687_ _03022_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__clkbuf_4
X_26475_ clknet_leaf_11_clk_sys _00106_ net604 VGND VGND VPWR VPWR top0.periodTop\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20899_ net229 net221 net214 _12681_ VGND VGND VPWR VPWR _12747_ sky130_fd_sc_hd__a31o_1
XFILLER_0_192_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13440_ net65 _05615_ _05652_ _05633_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__o211ai_4
X_25426_ _04406_ _04745_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22638_ net110 _02190_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25357_ _04664_ _04701_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__xnor2_1
X_13371_ _05561_ _05562_ _05583_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22569_ _02122_ _02123_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_196_Left_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15110_ _07203_ _07208_ VGND VGND VPWR VPWR _07209_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24308_ _03130_ _03135_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__and2_1
X_16090_ _08108_ _08119_ _08106_ VGND VGND VPWR VPWR _08183_ sky130_fd_sc_hd__a21bo_1
X_25288_ _04630_ _04633_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__xor2_1
XFILLER_0_107_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15041_ top0.pid_d.prev_int\[11\] _07139_ _07143_ top0.pid_d.curr_int\[11\] VGND
+ VGND VPWR VPWR _00128_ sky130_fd_sc_hd__a22o_1
X_24239_ _03583_ _03585_ _03563_ _03565_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__a211o_1
X_27027_ clknet_leaf_15_clk_sys _00644_ net614 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18800_ net383 net309 VGND VGND VPWR VPWR _10776_ sky130_fd_sc_hd__nand2_1
X_19780_ _11640_ _11641_ VGND VGND VPWR VPWR _11662_ sky130_fd_sc_hd__nand2_1
X_16992_ top0.pid_q.prev_error\[11\] top0.pid_q.curr_error\[11\] VGND VGND VPWR VPWR
+ _09047_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_196_Right_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18731_ _10636_ _10638_ _10637_ VGND VGND VPWR VPWR _10708_ sky130_fd_sc_hd__o21ai_1
X_15943_ _08026_ _08037_ VGND VGND VPWR VPWR _08038_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18662_ _10636_ _10639_ VGND VGND VPWR VPWR _10640_ sky130_fd_sc_hd__xnor2_1
X_15874_ net505 net483 VGND VGND VPWR VPWR _07970_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17613_ _09565_ _09563_ _09592_ _09598_ _09599_ VGND VGND VPWR VPWR _09600_ sky130_fd_sc_hd__o221a_1
X_14825_ _07021_ _07024_ VGND VGND VPWR VPWR _07025_ sky130_fd_sc_hd__nor2_1
X_18593_ _10570_ _10571_ VGND VGND VPWR VPWR _10572_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_4__f_clk_sys clknet_0_clk_sys VGND VGND VPWR VPWR clknet_3_4__leaf_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_169_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17544_ net417 net358 VGND VGND VPWR VPWR _09531_ sky130_fd_sc_hd__nand2_1
X_14756_ _06924_ _06833_ VGND VGND VPWR VPWR _06958_ sky130_fd_sc_hd__and2b_1
XFILLER_0_153_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13707_ _05913_ _05918_ _05919_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17475_ net400 net394 net359 VGND VGND VPWR VPWR _09462_ sky130_fd_sc_hd__o21ai_1
X_14687_ _06889_ _06890_ VGND VGND VPWR VPWR _06891_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19214_ net342 _11117_ _11163_ _10067_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__o211a_1
X_16426_ _08422_ _08423_ _08514_ VGND VGND VPWR VPWR _08515_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_144_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13638_ _05830_ _05848_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19145_ top0.kid\[7\] _11098_ _11100_ top0.kpd\[7\] VGND VGND VPWR VPWR _11108_ sky130_fd_sc_hd__a22o_1
X_16357_ _08048_ _08340_ VGND VGND VPWR VPWR _08447_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13569_ _05779_ _05781_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15308_ net539 net478 VGND VGND VPWR VPWR _07407_ sky130_fd_sc_hd__nand2_1
X_19076_ _10957_ _11012_ VGND VGND VPWR VPWR _11048_ sky130_fd_sc_hd__nor2_1
X_16288_ _08270_ _08281_ _08378_ VGND VGND VPWR VPWR _08379_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18027_ _10010_ _10011_ VGND VGND VPWR VPWR _10012_ sky130_fd_sc_hd__xnor2_1
X_15239_ net520 net493 _07228_ VGND VGND VPWR VPWR _07338_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout207 top0.state\[1\] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_4
Xfanout218 net220 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_201_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout229 net230 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_8
X_19978_ _11509_ _11845_ _11413_ VGND VGND VPWR VPWR _11846_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_163_Right_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18929_ _10901_ _10902_ VGND VGND VPWR VPWR _10904_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21940_ net164 _01501_ _01295_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21871_ _01399_ _01390_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23610_ top0.matmul0.alpha_pass\[12\] _09320_ net559 VGND VGND VPWR VPWR _02972_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20822_ _12400_ _12417_ _12670_ VGND VGND VPWR VPWR _12671_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24590_ _03939_ _03944_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23541_ _02936_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__clkbuf_1
X_20753_ _12587_ _12588_ VGND VGND VPWR VPWR _12602_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26260_ spi0.data_packed\[28\] spi0.data_packed\[29\] net699 VGND VGND VPWR VPWR
+ _05362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23472_ _02900_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__clkbuf_1
X_20684_ _12516_ _12531_ _12532_ VGND VGND VPWR VPWR _12533_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_46_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25211_ _04484_ _04556_ _04557_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__a21o_1
X_22423_ net95 _01902_ _01845_ net91 VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_174_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26191_ spi0.data_packed\[11\] _05321_ net18 VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25142_ _04480_ _04489_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22354_ net123 _01910_ _01912_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21305_ _13146_ _13147_ _12883_ VGND VGND VPWR VPWR _13148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25073_ _02982_ _04182_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22285_ _01844_ _01550_ _01214_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__a21o_2
X_24024_ _03380_ _03381_ _03010_ _03157_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21236_ _12616_ VGND VGND VPWR VPWR _13080_ sky130_fd_sc_hd__inv_2
Xhold250 _05379_ VGND VGND VPWR VPWR net950 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold261 top0.pid_d.prev_error\[1\] VGND VGND VPWR VPWR net961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 top0.svm0.delta\[12\] VGND VGND VPWR VPWR net972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 top0.pid_q.curr_error\[1\] VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 top0.b_in_matmul\[14\] VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__dlygate4sd3_1
X_21167_ _12952_ _13011_ _12883_ VGND VGND VPWR VPWR _13012_ sky130_fd_sc_hd__o21a_1
XFILLER_0_102_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20118_ top0.cordic0.gm0.iter\[4\] _11974_ VGND VGND VPWR VPWR _11975_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25975_ _05181_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__clkbuf_1
X_21098_ _12746_ _12943_ VGND VGND VPWR VPWR _12944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24926_ _04180_ _04181_ _04183_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_137_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20049_ _11650_ _11912_ net1020 VGND VGND VPWR VPWR _11913_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24857_ _04206_ _04208_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__xnor2_1
X_14610_ _06685_ _06744_ _06813_ _06814_ VGND VGND VPWR VPWR _06815_ sky130_fd_sc_hd__o22a_1
XFILLER_0_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23808_ _03160_ _03165_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__xnor2_4
X_15590_ _07255_ _07604_ _07595_ _07594_ VGND VGND VPWR VPWR _07689_ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24788_ _04125_ _04140_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__xnor2_2
X_14541_ _06691_ _06747_ VGND VGND VPWR VPWR _06748_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26527_ clknet_leaf_61_clk_sys _00150_ net647 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_23739_ _03073_ _03074_ _03096_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__nand3_1
XFILLER_0_83_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17260_ _09259_ _09260_ VGND VGND VPWR VPWR _09261_ sky130_fd_sc_hd__xnor2_1
X_14472_ _06678_ _06679_ _06551_ VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__mux2_1
X_26458_ clknet_leaf_88_clk_sys _00099_ net642 VGND VGND VPWR VPWR top0.kiq\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16211_ _08285_ _08302_ VGND VGND VPWR VPWR _08303_ sky130_fd_sc_hd__xor2_1
X_25409_ _04721_ _04752_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__xnor2_1
X_13423_ _05615_ _05635_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__xnor2_2
X_17191_ top0.pid_q.prev_int\[8\] VGND VGND VPWR VPWR _09201_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26389_ clknet_leaf_39_clk_sys _00030_ net677 VGND VGND VPWR VPWR top0.svm0.tC\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13354_ _05566_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__buf_2
X_16142_ _08163_ _08234_ VGND VGND VPWR VPWR _08235_ sky130_fd_sc_hd__xnor2_1
X_13285_ _05487_ _05492_ _05497_ net42 VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__o211a_1
X_16073_ _08124_ _08125_ _08126_ VGND VGND VPWR VPWR _08166_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15024_ net435 _07138_ _05443_ VGND VGND VPWR VPWR _07139_ sky130_fd_sc_hd__o21a_2
X_19901_ net190 _11774_ VGND VGND VPWR VPWR _11775_ sky130_fd_sc_hd__or2_2
X_19832_ _11710_ VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19763_ _11643_ _11645_ VGND VGND VPWR VPWR _11646_ sky130_fd_sc_hd__xor2_1
X_16975_ net429 top0.currT_r\[10\] VGND VGND VPWR VPWR _09031_ sky130_fd_sc_hd__and2b_1
XFILLER_0_127_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18714_ net377 _10690_ _09364_ VGND VGND VPWR VPWR _10691_ sky130_fd_sc_hd__and3_1
X_15926_ net448 net529 VGND VGND VPWR VPWR _08021_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19694_ net193 net182 net187 net179 VGND VGND VPWR VPWR _11580_ sky130_fd_sc_hd__a31o_1
X_18645_ _10456_ _10552_ VGND VGND VPWR VPWR _10623_ sky130_fd_sc_hd__and2b_1
X_15857_ _07833_ _07835_ _07834_ VGND VGND VPWR VPWR _07953_ sky130_fd_sc_hd__o21a_1
XFILLER_0_189_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14808_ _06910_ _06992_ _07003_ _07007_ VGND VGND VPWR VPWR _07008_ sky130_fd_sc_hd__a31o_1
XFILLER_0_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18576_ _10549_ _10554_ VGND VGND VPWR VPWR _10555_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_148_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15788_ _07765_ _07884_ _07770_ VGND VGND VPWR VPWR _07885_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17527_ _09467_ _09513_ VGND VGND VPWR VPWR _09514_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14739_ _06939_ _06941_ VGND VGND VPWR VPWR _06942_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17458_ _09437_ _09444_ VGND VGND VPWR VPWR _09445_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16409_ net452 net506 VGND VGND VPWR VPWR _08498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17389_ _09373_ _09375_ VGND VGND VPWR VPWR _09376_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19128_ _11097_ VGND VGND VPWR VPWR _11098_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19059_ top0.pid_d.out\[13\] top0.pid_d.curr_int\[13\] _10911_ _10915_ _10910_ VGND
+ VGND VPWR VPWR _11032_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22070_ _01565_ _01630_ _01631_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_100_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21021_ _12752_ _12866_ _12867_ VGND VGND VPWR VPWR _12868_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_77_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22972_ _06277_ _02481_ net172 VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__o21ai_1
X_25760_ top0.matmul0.matmul_stage_inst.a\[8\] _04897_ _05457_ VGND VGND VPWR VPWR
+ _05001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24711_ _03963_ _04059_ _04060_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__o21ai_1
X_21923_ _01106_ _01107_ _01458_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25691_ net72 _04885_ top0.matmul0.sin\[13\] _04954_ VGND VGND VPWR VPWR _04958_
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_171_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24642_ _03018_ _03019_ _03054_ _03055_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__o22a_1
X_21854_ net158 _01178_ _01415_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20805_ _11608_ _12278_ VGND VGND VPWR VPWR _12654_ sky130_fd_sc_hd__or2_1
X_24573_ _03899_ _03927_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__xnor2_2
X_21785_ _01337_ _01340_ _01341_ _01343_ _01346_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__a311o_1
X_26312_ spi0.data_packed\[54\] spi0.data_packed\[55\] net698 VGND VGND VPWR VPWR
+ _05388_ sky130_fd_sc_hd__mux2_1
X_20736_ _12348_ _12584_ _12553_ VGND VGND VPWR VPWR _12585_ sky130_fd_sc_hd__mux2_1
X_23524_ net979 top0.matmul0.a\[2\] _02926_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27292_ clknet_3_0__leaf_clk_mosi _00906_ VGND VGND VPWR VPWR spi0.data_packed\[78\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23455_ _02877_ _02889_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__nor2_1
X_26243_ _05353_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__clkbuf_1
X_20667_ _12515_ VGND VGND VPWR VPWR _12516_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22406_ _01112_ _01963_ net127 VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__o21a_1
XFILLER_0_190_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23386_ _02824_ _02826_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__xnor2_2
X_26174_ spi0.data_packed\[8\] _05311_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__xnor2_1
X_20598_ _12272_ _12347_ VGND VGND VPWR VPWR _12447_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25125_ _04461_ _04463_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22337_ _01809_ _01891_ _01895_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_182_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25056_ _04395_ _04391_ _04392_ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__a21o_1
X_22268_ _01758_ _01763_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24007_ _03325_ _03363_ _03324_ _03364_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__a31o_1
X_21219_ _12544_ _12545_ _12578_ _12646_ VGND VGND VPWR VPWR _13063_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22199_ net77 net92 VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__xnor2_1
Xfanout560 net561 VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__buf_4
Xfanout571 top0.matmul0.matmul_stage_inst.state\[2\] VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__clkbuf_2
Xfanout582 net584 VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__clkbuf_4
X_16760_ top0.pid_q.out\[14\] top0.pid_q.curr_int\[14\] VGND VGND VPWR VPWR _08844_
+ sky130_fd_sc_hd__nand2_1
X_13972_ _06183_ _06184_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__xnor2_1
Xfanout593 net597 VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__clkbuf_4
X_25958_ _12030_ _05015_ net207 _08900_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__a211oi_4
X_15711_ _07531_ _07614_ VGND VGND VPWR VPWR _07808_ sky130_fd_sc_hd__nor2_1
X_24909_ _04219_ _04220_ _04259_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__o21a_2
X_16691_ _08769_ _08775_ VGND VGND VPWR VPWR _08776_ sky130_fd_sc_hd__xnor2_1
X_25889_ _05104_ _05105_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18430_ _10399_ _10410_ VGND VGND VPWR VPWR _10411_ sky130_fd_sc_hd__xnor2_1
X_15642_ net462 net522 VGND VGND VPWR VPWR _07740_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18361_ _10339_ _10340_ VGND VGND VPWR VPWR _10342_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15573_ _07288_ _07286_ _07291_ VGND VGND VPWR VPWR _07672_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17312_ _09304_ _09300_ top0.matmul0.matmul_stage_inst.mult1\[9\] VGND VGND VPWR
+ VPWR _09305_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_139_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14524_ _06616_ _06617_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__nor2_1
X_18292_ _10272_ _10273_ VGND VGND VPWR VPWR _10274_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17243_ top0.pid_q.curr_int\[15\] top0.pid_q.prev_int\[15\] VGND VGND VPWR VPWR _09247_
+ sky130_fd_sc_hd__xnor2_1
X_14455_ _06596_ _06594_ VGND VGND VPWR VPWR _06663_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13406_ _05618_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__buf_4
XFILLER_0_25_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17174_ top0.pid_q.prev_int\[5\] _09172_ _09185_ top0.pid_q.prev_int\[6\] VGND VGND
+ VPWR VPWR _09186_ sky130_fd_sc_hd__a211o_1
X_14386_ net51 _06351_ _06489_ _06490_ VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16125_ _08092_ _08135_ _08121_ VGND VGND VPWR VPWR _08218_ sky130_fd_sc_hd__a21bo_1
X_13337_ _05536_ _05543_ _05545_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16056_ _08001_ _08007_ _08008_ VGND VGND VPWR VPWR _08150_ sky130_fd_sc_hd__a21o_1
X_13268_ _05477_ _05480_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__xor2_1
X_15007_ spi0.data_packed\[9\] top0.periodTop\[9\] _07125_ VGND VGND VPWR VPWR _07129_
+ sky130_fd_sc_hd__mux2_1
X_13199_ spi0.opcode\[0\] spi0.opcode\[2\] spi0.opcode\[3\] spi0.opcode\[4\] VGND
+ VGND VPWR VPWR _05429_ sky130_fd_sc_hd__or4_2
X_19815_ _11684_ _11690_ _11694_ VGND VGND VPWR VPWR _11695_ sky130_fd_sc_hd__o21a_1
XFILLER_0_159_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16958_ top0.currT_r\[10\] _08900_ _09013_ VGND VGND VPWR VPWR _09015_ sky130_fd_sc_hd__or3_1
X_19746_ net194 net203 VGND VGND VPWR VPWR _11629_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15909_ net499 _08003_ VGND VGND VPWR VPWR _08004_ sky130_fd_sc_hd__nand2_1
X_19677_ net179 net84 _11560_ _11563_ VGND VGND VPWR VPWR _11564_ sky130_fd_sc_hd__a22o_1
X_16889_ top0.pid_q.curr_error\[4\] _08939_ _08950_ VGND VGND VPWR VPWR _08951_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18628_ _10579_ _10600_ _10601_ _10433_ _10605_ VGND VGND VPWR VPWR _10606_ sky130_fd_sc_hd__a221o_2
XFILLER_0_52_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18559_ net320 net379 VGND VGND VPWR VPWR _10538_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_53_clk_sys clknet_3_6__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_53_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_21570_ _01074_ _01131_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__or2b_1
XANTENNA_12 net1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20521_ _11739_ _12317_ VGND VGND VPWR VPWR _12370_ sky130_fd_sc_hd__nor2_2
XFILLER_0_7_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_23 net237 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 net1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_45 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23240_ net297 net291 net286 net279 net198 net192 VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__mux4_1
XFILLER_0_172_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20452_ net274 net294 VGND VGND VPWR VPWR _12301_ sky130_fd_sc_hd__or2b_1
XFILLER_0_104_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23171_ _02641_ _06907_ _02645_ net989 VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20383_ _12148_ _12149_ _12133_ VGND VGND VPWR VPWR _12232_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_70_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22122_ _01258_ _01683_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__nand2_2
XFILLER_0_141_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22053_ net115 net97 VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__nand2_2
X_26930_ clknet_leaf_3_clk_sys _00547_ net583 VGND VGND VPWR VPWR top0.matmul0.cos\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_21004_ net238 _12134_ _12269_ _12850_ _12197_ VGND VGND VPWR VPWR _12851_ sky130_fd_sc_hd__a221o_4
X_26861_ clknet_leaf_40_clk_sys _00478_ net682 VGND VGND VPWR VPWR top0.svm0.tA\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25812_ top0.c_out_calc\[1\] _05029_ _05031_ _05038_ VGND VGND VPWR VPWR _00732_
+ sky130_fd_sc_hd__a22o_1
X_26792_ clknet_leaf_0_clk_sys _00409_ net578 VGND VGND VPWR VPWR top0.cordic0.sin\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25743_ net711 _04925_ _04992_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__a21o_1
Xmax_cap14 _07141_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
XFILLER_0_202_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22955_ _02458_ _02461_ _02332_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__o21a_1
XFILLER_0_173_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21906_ _01465_ _01466_ _01467_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__and3_1
XFILLER_0_179_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25674_ net71 _04944_ _04945_ net74 _05456_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__a221o_1
X_22886_ net168 VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__inv_2
X_24625_ _03829_ _03974_ _03315_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__a21o_1
X_21837_ _01381_ _01382_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__nand2_2
XFILLER_0_195_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24556_ _03045_ _03046_ _03162_ _03163_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__o22a_1
X_21768_ net142 net135 VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20719_ _12156_ _12327_ _12506_ VGND VGND VPWR VPWR _12568_ sky130_fd_sc_hd__and3_1
X_23507_ net771 top0.matmul0.cos\[8\] _02915_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__mux2_1
X_27275_ clknet_3_7__leaf_clk_mosi _00889_ VGND VGND VPWR VPWR spi0.data_packed\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24487_ _03738_ _03745_ _03746_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__a21o_1
X_21699_ _01259_ _01260_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__or2b_1
XFILLER_0_124_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14240_ _06448_ _06449_ _06417_ _06418_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__o211ai_2
X_26226_ spi0.data_packed\[11\] spi0.data_packed\[12\] net695 VGND VGND VPWR VPWR
+ _05345_ sky130_fd_sc_hd__mux2_1
X_23438_ _02873_ _02874_ _01166_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14171_ _06255_ _06256_ _06370_ VGND VGND VPWR VPWR _06382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23369_ _11518_ _02796_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__nand2_1
X_26157_ _05298_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25108_ _04347_ _04379_ _04456_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__a21oi_1
X_26088_ top0.pid_d.out\[14\] _12031_ _05013_ spi0.data_packed\[78\] VGND VGND VPWR
+ VPWR _05268_ sky130_fd_sc_hd__a22o_1
X_17930_ _09907_ _09915_ VGND VGND VPWR VPWR _09916_ sky130_fd_sc_hd__xnor2_2
X_25039_ _04268_ _04301_ _04388_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__a21o_1
X_17861_ _09844_ _09847_ VGND VGND VPWR VPWR _09848_ sky130_fd_sc_hd__xnor2_2
X_19600_ top0.cordic0.slte0.opA\[7\] _11487_ VGND VGND VPWR VPWR _11489_ sky130_fd_sc_hd__or2_1
X_16812_ top0.pid_q.mult0.a\[15\] _08855_ _08858_ net937 _08879_ VGND VGND VPWR VPWR
+ _00164_ sky130_fd_sc_hd__a221o_1
X_17792_ _09777_ _09778_ VGND VGND VPWR VPWR _09779_ sky130_fd_sc_hd__xor2_1
XFILLER_0_108_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout390 net391 VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_4
X_19531_ _11415_ _11416_ _11417_ _11418_ _11419_ _11420_ VGND VGND VPWR VPWR _11421_
+ sky130_fd_sc_hd__mux4_1
X_16743_ _07781_ net445 _08141_ _08826_ _08287_ VGND VGND VPWR VPWR _08827_ sky130_fd_sc_hd__a32o_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13955_ _06164_ _06165_ _06138_ _06161_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19462_ _11357_ _11353_ _10756_ VGND VGND VPWR VPWR _11358_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16674_ net447 net500 VGND VGND VPWR VPWR _08759_ sky130_fd_sc_hd__nand2_1
X_13886_ _06095_ _06098_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_202_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18413_ _10380_ _10393_ VGND VGND VPWR VPWR _10394_ sky130_fd_sc_hd__xor2_2
XFILLER_0_97_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15625_ _07719_ _07722_ VGND VGND VPWR VPWR _07723_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19393_ top0.pid_d.curr_int\[1\] top0.pid_d.prev_int\[1\] VGND VGND VPWR VPWR _11298_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_189_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18344_ _10325_ VGND VGND VPWR VPWR _10326_ sky130_fd_sc_hd__inv_2
XFILLER_0_201_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15556_ _07649_ _07654_ VGND VGND VPWR VPWR _07655_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14507_ _06649_ _06713_ VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18275_ net401 _10203_ _09363_ VGND VGND VPWR VPWR _10257_ sky130_fd_sc_hd__o21ai_1
X_15487_ _07546_ _07547_ _07585_ VGND VGND VPWR VPWR _07586_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17226_ top0.pid_q.curr_int\[13\] top0.pid_q.prev_int\[13\] VGND VGND VPWR VPWR _09232_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14438_ _06644_ _06645_ VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17157_ top0.pid_q.prev_int\[4\] _09165_ top0.pid_q.curr_int\[4\] VGND VGND VPWR
+ VPWR _09171_ sky130_fd_sc_hd__a21o_1
X_14369_ _06523_ _06525_ VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16108_ net458 net1029 VGND VGND VPWR VPWR _08201_ sky130_fd_sc_hd__and2_1
X_17088_ net897 _09115_ _09120_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__a21o_1
X_16039_ _08045_ _08050_ _08051_ VGND VGND VPWR VPWR _08133_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19729_ net188 net179 VGND VGND VPWR VPWR _11613_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_9_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22740_ _02285_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22671_ _02215_ _02221_ _02222_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__a21boi_2
X_24410_ _03765_ net1017 _03681_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__or3b_1
XFILLER_0_137_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21622_ _01174_ _01182_ _01183_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_181_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25390_ _03123_ _04676_ _03124_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24341_ _03695_ _03696_ _03697_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_63_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21553_ net105 net86 VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_16_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20504_ net303 _12346_ _12350_ _12352_ VGND VGND VPWR VPWR _12353_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24272_ _03290_ _03629_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__xnor2_4
X_27060_ clknet_leaf_21_clk_sys _00677_ net610 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.d\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_21484_ net227 net219 _01047_ net231 net223 VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26011_ _05209_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__clkbuf_1
X_23223_ _11650_ _02673_ net1020 VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20435_ net302 _11437_ VGND VGND VPWR VPWR _12284_ sky130_fd_sc_hd__nor2_2
XFILLER_0_132_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23154_ net171 net9 top0.svm0.rising VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__a21bo_1
X_20366_ net291 net265 VGND VGND VPWR VPWR _12215_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22105_ _01172_ _01666_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23085_ net170 _02567_ _02568_ _02566_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__a22oi_1
X_20297_ _12139_ _12141_ _12145_ VGND VGND VPWR VPWR _12146_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22036_ _01595_ _01597_ _01316_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__a21bo_1
X_26913_ clknet_leaf_2_clk_sys _00530_ net582 VGND VGND VPWR VPWR top0.matmul0.sin\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26844_ clknet_leaf_44_clk_sys _00461_ net681 VGND VGND VPWR VPWR top0.svm0.delta\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26775_ clknet_leaf_7_clk_sys _00392_ net593 VGND VGND VPWR VPWR top0.cordic0.cos\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23987_ _03342_ _03344_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__and2_1
X_13740_ _05879_ _05880_ _05878_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25726_ top0.matmul0.sin\[9\] _04981_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__xnor2_1
X_22938_ _02443_ _02444_ _02445_ _02347_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13671_ _05834_ _05835_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25657_ _04883_ top0.matmul0.sin\[6\] _04926_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__nand3_1
X_22869_ top0.svm0.tB\[5\] _02387_ _02331_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15410_ _07501_ _07508_ _07490_ _07489_ VGND VGND VPWR VPWR _07509_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24608_ _03954_ _03956_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16390_ net545 _08408_ _08409_ net549 _08479_ VGND VGND VPWR VPWR _08480_ sky130_fd_sc_hd__a32o_1
X_25588_ net70 top0.matmul0.cos\[0\] VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__and2_1
X_15341_ _07436_ _07439_ VGND VGND VPWR VPWR _07440_ sky130_fd_sc_hd__xnor2_4
X_24539_ _03890_ _03891_ _03892_ _03893_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_26_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18060_ _09616_ net307 VGND VGND VPWR VPWR _10045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27258_ clknet_3_3__leaf_clk_mosi _00872_ VGND VGND VPWR VPWR spi0.data_packed\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_15272_ _07365_ _07370_ VGND VGND VPWR VPWR _07371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17011_ net448 _08890_ _09064_ _08930_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14223_ _06431_ _06432_ _06425_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__a21oi_2
X_26209_ _05336_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27189_ clknet_leaf_54_clk_sys _00803_ net668 VGND VGND VPWR VPWR top0.currT_r\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14154_ _06249_ _06359_ _06365_ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14085_ _06229_ _06231_ _06226_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__a21oi_1
X_18962_ _10880_ _10884_ _10845_ VGND VGND VPWR VPWR _10936_ sky130_fd_sc_hd__a21o_1
X_17913_ top0.pid_d.out\[1\] top0.pid_d.curr_int\[1\] VGND VGND VPWR VPWR _09899_
+ sky130_fd_sc_hd__xor2_1
X_18893_ net380 net308 VGND VGND VPWR VPWR _10868_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17844_ _09827_ _09830_ VGND VGND VPWR VPWR _09831_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17775_ net378 net359 VGND VGND VPWR VPWR _09762_ sky130_fd_sc_hd__nand2_1
X_14987_ _07118_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__clkbuf_1
X_16726_ net449 net452 net455 VGND VGND VPWR VPWR _08810_ sky130_fd_sc_hd__nor3_1
X_19514_ _11028_ _11029_ _11077_ VGND VGND VPWR VPWR _11405_ sky130_fd_sc_hd__mux2_1
X_13938_ _06147_ _06150_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19445_ _11342_ _11336_ VGND VGND VPWR VPWR _11343_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16657_ top0.pid_q.out\[13\] _07705_ _08742_ net544 VGND VGND VPWR VPWR _08743_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13869_ _05860_ _05908_ _05955_ _06081_ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15608_ _07706_ _07704_ VGND VGND VPWR VPWR _07707_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19376_ net889 _11285_ _11288_ top0.pid_d.curr_error\[9\] VGND VGND VPWR VPWR _00319_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16588_ _08593_ _08592_ VGND VGND VPWR VPWR _08675_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18327_ net411 net406 _09967_ VGND VGND VPWR VPWR _10309_ sky130_fd_sc_hd__and3_1
X_15539_ net465 net522 VGND VGND VPWR VPWR _07638_ sky130_fd_sc_hd__nand2_2
XFILLER_0_151_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18258_ _10236_ _10240_ VGND VGND VPWR VPWR _10241_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17209_ _09215_ _09209_ _09216_ VGND VGND VPWR VPWR _09217_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18189_ _10168_ _10171_ VGND VGND VPWR VPWR _10172_ sky130_fd_sc_hd__xnor2_2
X_20220_ _12064_ _12068_ VGND VGND VPWR VPWR _12069_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20151_ spi0.data_packed\[14\] top0.cordic0.domain\[0\] _12004_ VGND VGND VPWR VPWR
+ _12005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20082_ _11940_ _11941_ VGND VGND VPWR VPWR _11943_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23910_ _03195_ _03200_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__nor2_1
X_24890_ _04166_ _04241_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__xnor2_1
X_23841_ _03195_ _03198_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__nor2_2
XFILLER_0_19_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26560_ clknet_leaf_52_clk_sys _00183_ net670 VGND VGND VPWR VPWR top0.pid_q.curr_error\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_23772_ _03119_ _03129_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__xor2_4
X_20984_ _12773_ _12829_ _12830_ _12818_ VGND VGND VPWR VPWR _12831_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25511_ _04841_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__clkbuf_1
X_22723_ net104 net100 _01852_ _01167_ net78 VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__o32a_1
X_26491_ clknet_leaf_67_clk_sys _00011_ net659 VGND VGND VPWR VPWR top0.pid_q.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25442_ _04518_ _04784_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__nor2_1
X_22654_ _02205_ _02206_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__or2_2
XFILLER_0_47_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21605_ _01063_ _01166_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__nor2_1
X_25373_ _04712_ _04713_ _04715_ _04716_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__o31ai_4
X_22585_ _02101_ _02116_ _02117_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_35_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27112_ clknet_leaf_87_clk_sys _00726_ net644 VGND VGND VPWR VPWR top0.pid_d.iterate_enable
+ sky130_fd_sc_hd__dfrtp_1
X_24324_ _02985_ _02987_ _03024_ _03025_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__o22a_2
XFILLER_0_63_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21536_ net143 _01090_ _01088_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27043_ clknet_leaf_16_clk_sys _00660_ net612 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24255_ _03478_ _03489_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__xnor2_1
X_21467_ _01030_ _01031_ net241 VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_177_Right_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20418_ net256 net245 VGND VGND VPWR VPWR _12267_ sky130_fd_sc_hd__xor2_2
X_23206_ _02657_ net217 _11775_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__mux2_1
X_24186_ _03542_ _03543_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__xnor2_1
X_21398_ _00932_ _00951_ _00952_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__a21o_1
X_23137_ _02514_ _02598_ _02625_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__and3_1
X_20349_ net238 _12136_ _12197_ VGND VGND VPWR VPWR _12198_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23068_ _05573_ _02565_ _02566_ _02567_ _02568_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__o221a_1
XFILLER_0_179_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22019_ _01281_ _01442_ _01580_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__or3b_1
XFILLER_0_41_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14910_ spi0.data_packed\[62\] top0.kpq\[14\] _07075_ VGND VGND VPWR VPWR _07076_
+ sky130_fd_sc_hd__mux2_1
X_15890_ _07983_ _07985_ VGND VGND VPWR VPWR _07986_ sky130_fd_sc_hd__xor2_1
X_14841_ net858 _06279_ _07038_ _05465_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__a22o_1
X_26827_ clknet_leaf_46_clk_sys _00444_ net680 VGND VGND VPWR VPWR top0.svm0.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_17560_ _09544_ _09546_ VGND VGND VPWR VPWR _09547_ sky130_fd_sc_hd__or2_1
X_14772_ net31 _06824_ _06954_ _06955_ VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__a22o_1
X_26758_ clknet_leaf_5_clk_sys _00375_ net590 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16511_ _08596_ _08598_ VGND VGND VPWR VPWR _08599_ sky130_fd_sc_hd__nand2_1
X_13723_ _05931_ _05935_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__or2_1
X_25709_ net819 _04964_ _04936_ _04970_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__a22o_1
X_17491_ _09407_ _09476_ _09477_ VGND VGND VPWR VPWR _09478_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26689_ clknet_leaf_84_clk_sys _00306_ net641 VGND VGND VPWR VPWR top0.pid_d.curr_error\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19230_ _11175_ _11176_ VGND VGND VPWR VPWR _11178_ sky130_fd_sc_hd__or2_1
X_16442_ _08529_ _08530_ VGND VGND VPWR VPWR _08531_ sky130_fd_sc_hd__or2b_1
XFILLER_0_183_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13654_ net63 net61 _05585_ _05587_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__and4_1
XFILLER_0_156_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19161_ top0.kid\[15\] _11097_ _11099_ top0.kpd\[15\] VGND VGND VPWR VPWR _11116_
+ sky130_fd_sc_hd__a22o_1
X_16373_ _08459_ _08462_ VGND VGND VPWR VPWR _08463_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13585_ _05788_ _05797_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18112_ _10024_ _10035_ _10022_ VGND VGND VPWR VPWR _10096_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_186_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15324_ _07420_ _07422_ VGND VGND VPWR VPWR _07423_ sky130_fd_sc_hd__xnor2_1
X_19092_ _10947_ _11008_ _11063_ net356 VGND VGND VPWR VPWR _11064_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18043_ _10026_ _10027_ VGND VGND VPWR VPWR _10028_ sky130_fd_sc_hd__xnor2_1
X_15255_ _07312_ _07353_ VGND VGND VPWR VPWR _07354_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14206_ _06408_ _06415_ _06416_ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__nand3_2
XFILLER_0_151_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15186_ _07283_ _07284_ VGND VGND VPWR VPWR _07285_ sky130_fd_sc_hd__xor2_2
X_14137_ net60 _06135_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19994_ net189 _11511_ VGND VGND VPWR VPWR _11861_ sky130_fd_sc_hd__nand2_1
X_14068_ _05465_ _06275_ _06280_ net736 VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__a22o_1
X_18945_ net436 _10909_ _10916_ net432 _10919_ VGND VGND VPWR VPWR _10920_ sky130_fd_sc_hd__a221o_1
XFILLER_0_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18876_ net380 net374 _10495_ VGND VGND VPWR VPWR _10851_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17827_ _09641_ _09645_ VGND VGND VPWR VPWR _09814_ sky130_fd_sc_hd__and2b_1
XFILLER_0_179_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17758_ _09718_ _09740_ _09742_ _09744_ VGND VGND VPWR VPWR _09745_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16709_ top0.pid_q.curr_int\[13\] _08740_ _08793_ VGND VGND VPWR VPWR _08794_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17689_ net413 net408 net333 net339 VGND VGND VPWR VPWR _09676_ sky130_fd_sc_hd__and4_1
XFILLER_0_130_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19428_ top0.pid_d.curr_int\[5\] _11290_ _11293_ _11328_ VGND VGND VPWR VPWR _00331_
+ sky130_fd_sc_hd__a22o_1
Xfanout18 net19 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
Xfanout29 top0.periodTop_r\[14\] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_99_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19359_ net910 _11275_ _11278_ _11247_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22370_ _01921_ _01928_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21321_ net242 _13124_ VGND VGND VPWR VPWR _13163_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24040_ _03393_ _03397_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__and2_1
XFILLER_0_142_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21252_ _12543_ _13094_ _13095_ _12738_ _12420_ VGND VGND VPWR VPWR _13096_ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_4_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20203_ _12044_ _12046_ _12051_ VGND VGND VPWR VPWR _12052_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21183_ net267 _13022_ _13026_ VGND VGND VPWR VPWR _13027_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_99_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20134_ _11985_ _11989_ _11428_ VGND VGND VPWR VPWR _11990_ sky130_fd_sc_hd__a21o_1
X_25991_ _05193_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__clkbuf_1
X_24942_ _04289_ _04292_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__xnor2_2
X_20065_ _11612_ net190 _11518_ VGND VGND VPWR VPWR _11927_ sky130_fd_sc_hd__and3_1
X_24873_ _04072_ _04223_ _04224_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__o21ba_1
X_26612_ clknet_leaf_30_clk_sys _00229_ net621 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_23824_ _02992_ _03001_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__and2_1
X_26543_ clknet_leaf_69_clk_sys _00166_ net662 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_23755_ _03057_ _03058_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__nor2_1
X_20967_ net236 net231 VGND VGND VPWR VPWR _12814_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22706_ _02241_ _02256_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__xnor2_1
X_26474_ clknet_leaf_12_clk_sys _00105_ net604 VGND VGND VPWR VPWR top0.periodTop\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23686_ _03008_ _03043_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_49_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20898_ _12720_ _12721_ _12745_ _12687_ VGND VGND VPWR VPWR _12746_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25425_ _04768_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22637_ _01118_ _01776_ _02189_ net77 VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25356_ _04668_ _04700_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__xnor2_2
X_13370_ _05561_ _05562_ net52 _05518_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__o211a_1
X_22568_ _02051_ _02073_ _02074_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_24_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24307_ _03168_ _03169_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__nor2_1
X_21519_ net160 net155 VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__nand2_2
X_25287_ _04632_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_134_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22499_ net107 _01312_ _02020_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__nor3_1
X_27026_ clknet_leaf_15_clk_sys _00643_ net617 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_15040_ top0.pid_d.prev_int\[10\] _07139_ _07143_ net828 VGND VGND VPWR VPWR _00127_
+ sky130_fd_sc_hd__a22o_1
X_24238_ _03583_ _03585_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__or2_1
XFILLER_0_181_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24169_ _03398_ _03400_ _03406_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16991_ top0.pid_q.prev_error\[12\] top0.pid_q.curr_error\[12\] VGND VGND VPWR VPWR
+ _09046_ sky130_fd_sc_hd__xor2_1
X_15942_ _08031_ _08036_ VGND VGND VPWR VPWR _08037_ sky130_fd_sc_hd__xnor2_2
X_18730_ _10688_ _10706_ VGND VGND VPWR VPWR _10707_ sky130_fd_sc_hd__xnor2_4
X_18661_ _10637_ _10638_ VGND VGND VPWR VPWR _10639_ sky130_fd_sc_hd__xnor2_1
X_15873_ net443 _07873_ _07968_ VGND VGND VPWR VPWR _07969_ sky130_fd_sc_hd__o21a_1
X_14824_ _06982_ _06985_ _07023_ _06964_ VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__o22a_1
X_17612_ _09594_ _09597_ VGND VGND VPWR VPWR _09599_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18592_ _10561_ _10569_ VGND VGND VPWR VPWR _10571_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17543_ net412 net403 net358 VGND VGND VPWR VPWR _09530_ sky130_fd_sc_hd__o21ai_1
X_14755_ _06953_ _06956_ VGND VGND VPWR VPWR _06957_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13706_ net67 net63 _05586_ _05588_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__and4_1
XFILLER_0_86_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17474_ _09363_ _09459_ _09460_ VGND VGND VPWR VPWR _09461_ sky130_fd_sc_hd__or3_1
XFILLER_0_50_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14686_ net33 _05666_ VGND VGND VPWR VPWR _06890_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16425_ _08422_ _08423_ _08421_ VGND VGND VPWR VPWR _08514_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19213_ net440 _11159_ _11162_ _11120_ _11123_ VGND VGND VPWR VPWR _11163_ sky130_fd_sc_hd__a221o_1
X_13637_ _05828_ _05849_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__or2_1
XFILLER_0_184_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19144_ net402 _11096_ _11107_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__a21o_1
X_16356_ _08371_ _08373_ _08445_ VGND VGND VPWR VPWR _08446_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_41_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13568_ _05678_ _05679_ _05780_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15307_ net1026 _07372_ VGND VGND VPWR VPWR _07406_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19075_ net324 net1022 net362 _10956_ VGND VGND VPWR VPWR _11047_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16287_ _08270_ _08281_ _08268_ VGND VGND VPWR VPWR _08378_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_70_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13499_ _05509_ _05529_ _05711_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18026_ net321 net409 VGND VGND VPWR VPWR _10011_ sky130_fd_sc_hd__nand2_1
X_15238_ _07335_ _07336_ VGND VGND VPWR VPWR _07337_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15169_ net522 net471 VGND VGND VPWR VPWR _07268_ sky130_fd_sc_hd__nand2_2
XFILLER_0_2_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout208 top0.state\[0\] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__buf_2
Xfanout219 net220 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_2
X_19977_ _11632_ net183 VGND VGND VPWR VPWR _11845_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18928_ _10901_ _10902_ VGND VGND VPWR VPWR _10903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18859_ _10834_ _10758_ top0.pid_d.out\[10\] VGND VGND VPWR VPWR _10835_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_59_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21870_ _01418_ _01431_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_173_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20821_ _12411_ _12414_ VGND VGND VPWR VPWR _12670_ sky130_fd_sc_hd__nor2_1
XFILLER_0_194_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23540_ top0.a_in_matmul\[10\] top0.matmul0.a\[10\] _02926_ VGND VGND VPWR VPWR _02936_
+ sky130_fd_sc_hd__mux2_1
X_20752_ _11593_ net258 _12589_ VGND VGND VPWR VPWR _12601_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20683_ _12530_ _12519_ _12520_ VGND VGND VPWR VPWR _12532_ sky130_fd_sc_hd__nand3_2
X_23471_ net920 top0.matmul0.sin\[5\] _05461_ VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25210_ _03758_ _03981_ _03123_ _03889_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__and4_1
XFILLER_0_147_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22422_ net79 net87 VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__nand2_2
XFILLER_0_190_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26190_ _05324_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25141_ _04483_ _04488_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22353_ _01225_ _01328_ _01911_ _01408_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21304_ _13014_ _13146_ _13145_ _13104_ VGND VGND VPWR VPWR _13147_ sky130_fd_sc_hd__a2bb2o_1
X_25072_ _03343_ _04272_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__nor2_1
X_22284_ net115 _01211_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24023_ _02998_ _03000_ _03027_ _03028_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__o22a_1
X_21235_ _13062_ _13065_ _13074_ _13078_ VGND VGND VPWR VPWR _13079_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold240 top0.pid_d.curr_error\[0\] VGND VGND VPWR VPWR net940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 top0.matmul0.b\[10\] VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 top0.currT_r\[7\] VGND VGND VPWR VPWR net962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 spi0.data_packed\[37\] VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 top0.pid_q.prev_error\[0\] VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__dlygate4sd3_1
X_21166_ _12960_ VGND VGND VPWR VPWR _13011_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_48_clk_sys clknet_3_7__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_48_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
Xhold295 top0.pid_q.prev_int\[2\] VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_176_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20117_ _11413_ _11515_ VGND VGND VPWR VPWR _11974_ sky130_fd_sc_hd__nor2_1
X_25974_ top0.b_in_matmul\[3\] _05180_ _05165_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__mux2_1
X_21097_ _12677_ _12728_ _12727_ VGND VGND VPWR VPWR _12943_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_102_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24925_ _04271_ _04275_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__xnor2_2
X_20048_ _11907_ _11911_ VGND VGND VPWR VPWR _11912_ sky130_fd_sc_hd__xor2_1
XFILLER_0_176_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24856_ _04107_ _04108_ _04207_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23807_ _03161_ _03164_ VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__nor2_2
X_24787_ _04128_ _04139_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_197_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21999_ _01290_ _01293_ _01295_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__or3b_1
XFILLER_0_96_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14540_ _06697_ _06746_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__xor2_2
XFILLER_0_185_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26526_ clknet_leaf_63_clk_sys _00149_ net647 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_23738_ _03092_ _03095_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14471_ _06554_ _06608_ _06676_ _06677_ VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__a22o_1
X_26457_ clknet_leaf_57_clk_sys _00098_ net642 VGND VGND VPWR VPWR top0.kiq\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23669_ net569 net573 top0.matmul0.matmul_stage_inst.f\[1\] VGND VGND VPWR VPWR _03027_
+ sky130_fd_sc_hd__o21a_4
X_16210_ _08296_ _08301_ VGND VGND VPWR VPWR _08302_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25408_ _04748_ _04751_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__xnor2_1
X_13422_ net65 _05619_ _05628_ _05634_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17190_ _08399_ _09192_ _09200_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26388_ clknet_leaf_38_clk_sys _00029_ net677 VGND VGND VPWR VPWR top0.svm0.tC\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16141_ _08231_ _08233_ VGND VGND VPWR VPWR _08234_ sky130_fd_sc_hd__nand2_1
X_25339_ _04619_ _04624_ _04617_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__a21o_1
X_13353_ _05493_ _05494_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16072_ _08090_ _08149_ _08164_ VGND VGND VPWR VPWR _08165_ sky130_fd_sc_hd__o21ai_1
X_13284_ _05496_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27009_ clknet_leaf_23_clk_sys _00626_ net625 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19900_ net194 net184 VGND VGND VPWR VPWR _11774_ sky130_fd_sc_hd__or2_1
X_15023_ _07137_ VGND VGND VPWR VPWR _07138_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19831_ _11708_ _11709_ net248 VGND VGND VPWR VPWR _11710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19762_ net272 _11621_ _11644_ VGND VGND VPWR VPWR _11645_ sky130_fd_sc_hd__a21oi_1
X_16974_ top0.currT_r\[9\] _08997_ top0.currT_r\[10\] VGND VGND VPWR VPWR _09030_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18713_ net374 VGND VGND VPWR VPWR _10690_ sky130_fd_sc_hd__inv_2
X_15925_ net536 net443 VGND VGND VPWR VPWR _08020_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_189_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19693_ net182 _11578_ VGND VGND VPWR VPWR _11579_ sky130_fd_sc_hd__or2_1
XFILLER_0_190_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15856_ _07948_ _07951_ VGND VGND VPWR VPWR _07952_ sky130_fd_sc_hd__xnor2_1
X_18644_ _10458_ _10552_ net341 VGND VGND VPWR VPWR _10622_ sky130_fd_sc_hd__o21a_1
X_14807_ _06989_ _06990_ _07005_ _06993_ _07006_ VGND VGND VPWR VPWR _07007_ sky130_fd_sc_hd__o221a_1
X_18575_ _10550_ _10553_ VGND VGND VPWR VPWR _10554_ sky130_fd_sc_hd__xor2_1
X_15787_ net508 _07618_ _07619_ VGND VGND VPWR VPWR _07884_ sky130_fd_sc_hd__or3_1
XFILLER_0_118_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14738_ _06870_ _06901_ _06940_ VGND VGND VPWR VPWR _06941_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17526_ _09504_ _09512_ VGND VGND VPWR VPWR _09513_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_188_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17457_ _09438_ _09439_ _09441_ _09375_ _09443_ VGND VGND VPWR VPWR _09444_ sky130_fd_sc_hd__o221a_1
X_14669_ _06716_ _06871_ _06872_ VGND VGND VPWR VPWR _06873_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16408_ net456 net503 VGND VGND VPWR VPWR _08497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17388_ _09346_ _09347_ _09374_ VGND VGND VPWR VPWR _09375_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_43_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16339_ _08350_ _08360_ _08428_ VGND VGND VPWR VPWR _08429_ sky130_fd_sc_hd__o21a_1
X_19127_ net437 _05442_ _11094_ VGND VGND VPWR VPWR _11097_ sky130_fd_sc_hd__and3_2
XFILLER_0_131_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19058_ _10992_ _11030_ VGND VGND VPWR VPWR _11031_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18009_ net411 net319 VGND VGND VPWR VPWR _09994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21020_ _12782_ _12800_ VGND VGND VPWR VPWR _12867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_199_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22971_ top0.svm0.delta\[7\] _02480_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__xnor2_1
X_24710_ _04063_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__clkbuf_1
X_21922_ _01106_ _01107_ _01208_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25690_ net714 _04925_ _04957_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__a21o_1
X_24641_ _03882_ _03897_ _03994_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21853_ _01411_ _01410_ _01380_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20804_ _11673_ _12559_ VGND VGND VPWR VPWR _12653_ sky130_fd_sc_hd__nor2_1
X_24572_ _03925_ _03926_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__or2_1
XFILLER_0_171_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21784_ _01344_ _01345_ _01337_ _01340_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26311_ _05387_ VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23523_ _02927_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20735_ net295 net282 VGND VGND VPWR VPWR _12584_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27291_ clknet_3_3__leaf_clk_mosi _00905_ VGND VGND VPWR VPWR spi0.data_packed\[77\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26242_ spi0.data_packed\[19\] spi0.data_packed\[20\] net697 VGND VGND VPWR VPWR
+ _05353_ sky130_fd_sc_hd__mux2_1
X_23454_ _11515_ _02878_ net89 VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20666_ _12501_ _12513_ _12514_ VGND VGND VPWR VPWR _12515_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_80_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22405_ _01065_ net110 VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__nor2_1
X_26173_ spi0.data_packed\[14\] _05310_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__nor2_1
X_20597_ _12440_ _12445_ VGND VGND VPWR VPWR _12446_ sky130_fd_sc_hd__or2_1
X_23385_ _11513_ _02825_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_36_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25124_ _04387_ _04389_ _04381_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__o21a_1
X_22336_ _01867_ _01868_ _01871_ _01894_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__o31a_1
X_25055_ _04334_ _04399_ _04403_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22267_ _11674_ _01825_ _01826_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__and3_1
X_24006_ _03325_ _03106_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21218_ _13057_ _13059_ _13060_ _13061_ VGND VGND VPWR VPWR _13062_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22198_ net95 net104 VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__or2b_1
XFILLER_0_40_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21149_ _12980_ _12993_ VGND VGND VPWR VPWR _12994_ sky130_fd_sc_hd__xnor2_1
Xfanout550 net552 VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__buf_2
Xfanout561 top0.matmul0.matmul_stage_inst.state\[6\] VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__clkbuf_4
Xfanout572 net573 VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__clkbuf_4
X_13971_ net45 _05611_ _05612_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__and3_1
Xfanout583 net584 VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__clkbuf_4
X_25957_ _05167_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_45_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout594 net596 VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__clkbuf_4
X_15710_ _07527_ _07528_ _07531_ _07614_ _07694_ VGND VGND VPWR VPWR _07807_ sky130_fd_sc_hd__a221o_1
X_24908_ _04219_ _04220_ _04218_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__a21o_1
X_16690_ _08771_ _08774_ VGND VGND VPWR VPWR _08775_ sky130_fd_sc_hd__xor2_1
X_25888_ _05104_ _05105_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__nand2_1
X_15641_ net465 net520 VGND VGND VPWR VPWR _07739_ sky130_fd_sc_hd__nand2_2
X_24839_ _02982_ _04190_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__nor2_1
XFILLER_0_200_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18360_ _10339_ _10340_ VGND VGND VPWR VPWR _10341_ sky130_fd_sc_hd__nand2_1
X_15572_ _07663_ _07670_ VGND VGND VPWR VPWR _07671_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17311_ top0.matmul0.matmul_stage_inst.mult2\[9\] VGND VGND VPWR VPWR _09304_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14523_ _06616_ _06617_ VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__nand2_1
X_26509_ clknet_leaf_77_clk_sys net816 net631 VGND VGND VPWR VPWR top0.pid_d.prev_int\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18291_ net334 net376 VGND VGND VPWR VPWR _10273_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17242_ _09239_ _09244_ _09245_ VGND VGND VPWR VPWR _09246_ sky130_fd_sc_hd__a21oi_1
X_14454_ _06597_ _06600_ VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__nand2_2
XFILLER_0_154_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_54_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13405_ _05616_ _05617_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__and2_1
X_17173_ top0.pid_q.prev_int\[5\] _09172_ top0.pid_q.curr_int\[5\] VGND VGND VPWR
+ VPWR _09185_ sky130_fd_sc_hd__o21a_1
X_14385_ _06581_ _06593_ VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_181_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16124_ _08182_ _08216_ VGND VGND VPWR VPWR _08217_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13336_ _05541_ _05531_ _05532_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__or3_1
XFILLER_0_107_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16055_ _08137_ _08148_ VGND VGND VPWR VPWR _08149_ sky130_fd_sc_hd__xnor2_2
X_13267_ net42 _05478_ _05479_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__and3_1
X_15006_ _07128_ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__clkbuf_1
X_13198_ spi0.opcode\[1\] spi0.opcode\[5\] spi0.opcode\[6\] spi0.opcode\[7\] VGND
+ VGND VPWR VPWR _05428_ sky130_fd_sc_hd__or4_2
XFILLER_0_47_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19814_ _11692_ _11693_ VGND VGND VPWR VPWR _11694_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_63_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19745_ net174 _11608_ _11627_ _11628_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__a31o_1
X_16957_ _08900_ _09013_ top0.currT_r\[10\] VGND VGND VPWR VPWR _09014_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_155_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15908_ net493 _07227_ _07228_ VGND VGND VPWR VPWR _08003_ sky130_fd_sc_hd__a21o_2
X_19676_ _11561_ _11562_ net187 VGND VGND VPWR VPWR _11563_ sky130_fd_sc_hd__mux2_1
X_16888_ top0.pid_q.curr_error\[4\] _08939_ top0.pid_q.prev_error\[4\] VGND VGND VPWR
+ VPWR _08950_ sky130_fd_sc_hd__a21o_1
X_18627_ _10443_ _10604_ VGND VGND VPWR VPWR _10605_ sky130_fd_sc_hd__nor2_1
X_15839_ net536 net446 VGND VGND VPWR VPWR _07935_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18558_ net327 net373 VGND VGND VPWR VPWR _10537_ sky130_fd_sc_hd__nand2_2
XFILLER_0_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17509_ net353 _09494_ _09495_ net390 VGND VGND VPWR VPWR _09496_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18489_ _10465_ _10468_ VGND VGND VPWR VPWR _10469_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_72_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_13 _12739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20520_ _12279_ _12364_ _12367_ _12368_ VGND VGND VPWR VPWR _12369_ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_24 net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 _08403_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_46 net1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20451_ net302 _12284_ net275 VGND VGND VPWR VPWR _12300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23170_ _02641_ _06860_ _02645_ net930 VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__a22o_1
X_20382_ _12133_ _12148_ _12149_ VGND VGND VPWR VPWR _12231_ sky130_fd_sc_hd__and3b_1
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22121_ _01197_ _01257_ _01679_ _01682_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22052_ _01174_ _01613_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__xnor2_4
XPHY_EDGE_ROW_81_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21003_ _11689_ net238 VGND VGND VPWR VPWR _12850_ sky130_fd_sc_hd__or2_1
X_26860_ clknet_leaf_36_clk_sys _00477_ net678 VGND VGND VPWR VPWR top0.svm0.tA\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_25811_ _05036_ _05037_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26791_ clknet_leaf_1_clk_sys _00408_ net578 VGND VGND VPWR VPWR top0.cordic0.sin\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25742_ net778 _04925_ _04992_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22954_ top0.svm0.delta\[5\] VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap15 net16 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_97_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21905_ _01135_ _01464_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__nand2_1
X_25673_ net71 top0.matmul0.sin\[9\] VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__nand2_1
X_22885_ _02317_ top0.svm0.tB\[13\] _02403_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__a21o_1
XFILLER_0_168_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24624_ _03741_ _03974_ _03977_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__o21a_1
X_21836_ _01327_ _01378_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_195_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_90_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24555_ _03015_ _03016_ _03741_ _03742_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__o22a_1
XFILLER_0_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21767_ _01216_ _01328_ net147 VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23506_ _02918_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27274_ clknet_3_7__leaf_clk_mosi _00888_ VGND VGND VPWR VPWR spi0.data_packed\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_20718_ _12265_ _12504_ VGND VGND VPWR VPWR _12567_ sky130_fd_sc_hd__nor2_1
X_24486_ _03735_ _03748_ _03841_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__a21bo_1
X_21698_ net139 net131 VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26225_ _05344_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23437_ _11784_ _02872_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__nor2_1
X_20649_ net280 net270 net253 VGND VGND VPWR VPWR _12498_ sky130_fd_sc_hd__and3_1
XFILLER_0_190_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14170_ net852 _06280_ _06380_ _06381_ VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__a22o_1
X_26156_ _05297_ top0.cordic0.slte0.opB\[6\] _12006_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23368_ _02809_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__inv_2
X_25107_ _04347_ _04379_ _04377_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22319_ _01873_ _01878_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__xor2_1
X_26087_ _05267_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__clkbuf_1
X_23299_ _02725_ _02734_ _02745_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25038_ _04268_ _04301_ _04270_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_44_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17860_ _09845_ _09846_ VGND VGND VPWR VPWR _09847_ sky130_fd_sc_hd__xnor2_1
X_16811_ top0.kiq\[15\] _05448_ _08854_ VGND VGND VPWR VPWR _08879_ sky130_fd_sc_hd__and3_1
X_17791_ net409 net332 VGND VGND VPWR VPWR _09778_ sky130_fd_sc_hd__nand2_1
X_26989_ clknet_leaf_28_clk_sys _00606_ net622 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout380 top0.pid_d.mult0.a\[11\] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkbuf_4
Xfanout391 net392 VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__clkbuf_4
X_19530_ net182 VGND VGND VPWR VPWR _11420_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13954_ _06163_ _06123_ _06128_ _06138_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__or4_1
X_16742_ net445 _08822_ net500 VGND VGND VPWR VPWR _08826_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16673_ _07781_ net444 VGND VGND VPWR VPWR _08758_ sky130_fd_sc_hd__nand2_1
X_19461_ top0.pid_d.prev_int\[9\] VGND VGND VPWR VPWR _11357_ sky130_fd_sc_hd__inv_2
XFILLER_0_202_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13885_ _06096_ _06097_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__xor2_1
XFILLER_0_158_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18412_ _10391_ _10392_ VGND VGND VPWR VPWR _10393_ sky130_fd_sc_hd__or2b_1
XFILLER_0_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15624_ _07720_ _07721_ VGND VGND VPWR VPWR _07722_ sky130_fd_sc_hd__xnor2_1
X_19392_ top0.pid_d.curr_int\[0\] top0.pid_d.prev_int\[0\] VGND VGND VPWR VPWR _11297_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18343_ _10318_ _10324_ VGND VGND VPWR VPWR _10325_ sky130_fd_sc_hd__xnor2_1
X_15555_ _07650_ _07653_ VGND VGND VPWR VPWR _07654_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14506_ _06704_ _06712_ VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_189_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18274_ _10254_ _10255_ _10214_ _10209_ VGND VGND VPWR VPWR _10256_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_51_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15486_ _07564_ _07584_ VGND VGND VPWR VPWR _07585_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14437_ net30 _05579_ VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__nand2_1
X_17225_ top0.pid_q.curr_int\[12\] top0.pid_q.prev_int\[12\] _09230_ VGND VGND VPWR
+ VPWR _09231_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17156_ top0.pid_q.curr_int\[4\] _09141_ _09170_ _09136_ VGND VGND VPWR VPWR _00217_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14368_ _06523_ _06525_ VGND VGND VPWR VPWR _06577_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16107_ _08097_ _08104_ _08199_ VGND VGND VPWR VPWR _08200_ sky130_fd_sc_hd__a21o_1
X_13319_ top0.matmul0.beta_pass\[6\] _05434_ _05469_ _05463_ top0.c_out_calc\[6\]
+ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__a32o_2
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17087_ top0.pid_q.curr_error\[2\] _00011_ _09117_ VGND VGND VPWR VPWR _09120_ sky130_fd_sc_hd__and3_1
X_14299_ _06504_ _06508_ VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__xor2_2
XFILLER_0_123_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16038_ _08033_ _08035_ _08131_ VGND VGND VPWR VPWR _08132_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17989_ _09972_ _09974_ VGND VGND VPWR VPWR _09975_ sky130_fd_sc_hd__xnor2_1
X_19728_ _11576_ VGND VGND VPWR VPWR _11612_ sky130_fd_sc_hd__clkbuf_4
X_19659_ _11526_ _11546_ VGND VGND VPWR VPWR _11547_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22670_ _01643_ _01063_ _01980_ _02215_ _02221_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__o32a_1
XFILLER_0_177_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21621_ _01180_ _01181_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_158_Right_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24340_ _03213_ _03221_ _03220_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__a21oi_2
X_21552_ _01111_ _01113_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20503_ net294 _12326_ _12351_ _11438_ VGND VGND VPWR VPWR _12352_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24271_ _03628_ _03287_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_117_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21483_ net242 net236 net227 net219 VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26010_ net980 _05208_ _05196_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23222_ _02669_ _02672_ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__xnor2_1
X_20434_ _12266_ _12282_ VGND VGND VPWR VPWR _12283_ sky130_fd_sc_hd__xor2_4
X_23153_ net171 _02305_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20365_ _11525_ _12212_ _12213_ VGND VGND VPWR VPWR _12214_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22104_ _01195_ _01087_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23084_ _02339_ _02539_ _02583_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__or3_1
X_20296_ net258 _12101_ _12142_ _12143_ _12144_ VGND VGND VPWR VPWR _12145_ sky130_fd_sc_hd__a221o_1
X_22035_ _01289_ _01596_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__xnor2_1
X_26912_ clknet_leaf_0_clk_sys _00529_ net578 VGND VGND VPWR VPWR top0.matmul0.sin\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_26843_ clknet_leaf_45_clk_sys _00460_ net681 VGND VGND VPWR VPWR top0.svm0.delta\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_199_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26774_ clknet_leaf_4_clk_sys _00391_ net580 VGND VGND VPWR VPWR top0.cordic0.cos\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_23986_ _03343_ _03149_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__nor2_2
XFILLER_0_138_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25725_ net74 _04941_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__nand2_1
X_22937_ _02451_ VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_119_Left_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13670_ _05846_ _05882_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25656_ top0.matmul0.sin\[6\] _04926_ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__or2_2
X_22868_ _02332_ top0.svm0.tB\[4\] _02386_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__a21o_1
XFILLER_0_183_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24607_ _03961_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__clkbuf_1
X_21819_ net142 _01380_ _01280_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__a21oi_1
X_25587_ _04881_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22799_ _02317_ top0.svm0.tA\[13\] VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__or2_1
XFILLER_0_195_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15340_ _07437_ _07438_ VGND VGND VPWR VPWR _07439_ sky130_fd_sc_hd__xnor2_2
X_24538_ _03790_ _03792_ _03791_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27257_ clknet_3_3__leaf_clk_mosi _00871_ VGND VGND VPWR VPWR spi0.data_packed\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_15271_ net525 _07368_ _07369_ _07321_ VGND VGND VPWR VPWR _07370_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_149_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24469_ _03805_ _03806_ VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__nand2_2
X_17010_ net551 _09055_ _09063_ _08882_ VGND VGND VPWR VPWR _09064_ sky130_fd_sc_hd__a211o_1
X_14222_ _06425_ _06431_ _06432_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__and3_2
XFILLER_0_11_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26208_ spi0.data_packed\[2\] spi0.data_packed\[3\] net694 VGND VGND VPWR VPWR _05336_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_128_Left_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27188_ clknet_leaf_56_clk_sys _00802_ net666 VGND VGND VPWR VPWR top0.currT_r\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_62_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14153_ net64 _06268_ _06244_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__and3_1
X_26139_ _05284_ top0.cordic0.slte0.opB\[2\] _12006_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14084_ _06229_ _06231_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__nor2_1
X_18961_ _10805_ _10875_ _10933_ _10845_ _10934_ VGND VGND VPWR VPWR _10935_ sky130_fd_sc_hd__o221a_2
XFILLER_0_120_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17912_ _09894_ _09898_ _07710_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__o21a_1
X_18892_ _10865_ _10866_ VGND VGND VPWR VPWR _10867_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_96_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_96_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_17843_ _09828_ _09829_ VGND VGND VPWR VPWR _09830_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_137_Left_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17774_ _09757_ _09760_ VGND VGND VPWR VPWR _09761_ sky130_fd_sc_hd__xnor2_2
X_14986_ top0.svm0.delta\[0\] _07117_ VGND VGND VPWR VPWR _07118_ sky130_fd_sc_hd__or2_1
X_19513_ net441 _11402_ _11403_ net435 _11268_ VGND VGND VPWR VPWR _11404_ sky130_fd_sc_hd__a32o_1
X_16725_ net449 net452 net455 VGND VGND VPWR VPWR _08809_ sky130_fd_sc_hd__and3_1
X_13937_ _06148_ _06149_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19444_ top0.pid_d.prev_int\[7\] VGND VGND VPWR VPWR _11342_ sky130_fd_sc_hd__inv_2
X_13868_ _06074_ _06078_ _06079_ _06080_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16656_ top0.pid_q.out\[13\] _08739_ _08741_ VGND VGND VPWR VPWR _08742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15607_ top0.pid_q.curr_int\[0\] VGND VGND VPWR VPWR _07706_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19375_ net876 _11285_ _11288_ top0.pid_d.curr_error\[8\] VGND VGND VPWR VPWR _00318_
+ sky130_fd_sc_hd__a22o_1
X_13799_ _06011_ _06010_ net68 _05586_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__o211ai_4
X_16587_ _08593_ _08592_ _08594_ VGND VGND VPWR VPWR _08674_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18326_ _10215_ _10218_ _10307_ VGND VGND VPWR VPWR _10308_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_85_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15538_ _07575_ _07580_ VGND VGND VPWR VPWR _07637_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18257_ _10238_ _10239_ VGND VGND VPWR VPWR _10240_ sky130_fd_sc_hd__xor2_1
X_15469_ _07566_ _07567_ VGND VGND VPWR VPWR _07568_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_182_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17208_ _09215_ _09209_ top0.pid_q.curr_int\[10\] VGND VGND VPWR VPWR _09216_ sky130_fd_sc_hd__o21ba_1
X_18188_ _10169_ _10170_ VGND VGND VPWR VPWR _10171_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17139_ top0.pid_q.curr_int\[2\] VGND VGND VPWR VPWR _09155_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20150_ _12003_ VGND VGND VPWR VPWR _12004_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20081_ _11940_ _11941_ VGND VGND VPWR VPWR _11942_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23840_ _03196_ _03197_ VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__nor2_2
XFILLER_0_197_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23771_ _03125_ _03128_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__xnor2_2
X_20983_ _12826_ _12819_ VGND VGND VPWR VPWR _12830_ sky130_fd_sc_hd__nor2_1
X_25510_ top0.matmul0.matmul_stage_inst.mult1\[11\] _04604_ _03148_ VGND VGND VPWR
+ VPWR _04841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22722_ _02237_ _02255_ _02271_ _02222_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26490_ clknet_leaf_63_clk_sys _00010_ net656 VGND VGND VPWR VPWR top0.pid_q.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25441_ _04782_ _04783_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22653_ _02202_ _02204_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__nor2_1
XFILLER_0_192_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21604_ net94 VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__clkinv_4
X_25372_ _04668_ _04714_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__nand2_1
XFILLER_0_192_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22584_ _02077_ _02135_ _02137_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_62_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27111_ clknet_leaf_9_clk_sys _00001_ net595 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.start
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24323_ _03502_ _03158_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__nand2_2
XFILLER_0_133_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21535_ top0.cordic0.vec\[1\]\[4\] _01096_ _01088_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27042_ clknet_leaf_8_clk_sys _00659_ net597 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_24254_ _03610_ _03611_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21466_ net232 _12832_ _12815_ _12697_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_44_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23205_ net223 net217 net203 VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__mux2_2
XFILLER_0_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20417_ _12263_ _12264_ _12265_ _12262_ VGND VGND VPWR VPWR _12266_ sky130_fd_sc_hd__o2bb2a_4
X_24185_ _03045_ _03046_ _03063_ _03064_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21397_ _00916_ _00927_ _00962_ _00963_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__a31o_2
X_23136_ _02483_ _02625_ _02596_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__o21ai_1
X_20348_ net246 net238 VGND VGND VPWR VPWR _12197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23067_ net44 _02367_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__nand2_1
X_20279_ net276 net283 VGND VGND VPWR VPWR _12128_ sky130_fd_sc_hd__or2b_1
X_22018_ net151 _01338_ _01579_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__mux2_1
X_14840_ _07033_ _07035_ _07036_ _07037_ net20 VGND VGND VPWR VPWR _07038_ sky130_fd_sc_hd__o311a_1
X_26826_ clknet_leaf_46_clk_sys _00443_ net680 VGND VGND VPWR VPWR top0.svm0.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_14771_ _06957_ _06959_ VGND VGND VPWR VPWR _06972_ sky130_fd_sc_hd__or2_1
X_23969_ _03078_ _03322_ _03323_ _03324_ _03326_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__o2111ai_4
X_26757_ clknet_leaf_94_clk_sys _00374_ net591 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_187_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13722_ _05932_ _05933_ _05934_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__a21o_1
X_16510_ _08492_ _08540_ _08597_ VGND VGND VPWR VPWR _08598_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25708_ top0.matmul0.sin\[3\] _04969_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__xor2_1
X_17490_ net419 net333 net422 net330 VGND VGND VPWR VPWR _09477_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26688_ clknet_leaf_83_clk_sys _00305_ net649 VGND VGND VPWR VPWR top0.pid_d.curr_error\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_129_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13653_ net61 _05585_ _05588_ net63 VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__a22o_1
X_16441_ _08528_ _08523_ VGND VGND VPWR VPWR _08530_ sky130_fd_sc_hd__or2b_1
X_25639_ _04915_ _04916_ net69 VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16372_ _08142_ _08461_ VGND VGND VPWR VPWR _08462_ sky130_fd_sc_hd__xnor2_1
X_19160_ net370 _11095_ _11115_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_52_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13584_ _05789_ _05794_ _05796_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_186_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18111_ _10088_ _10094_ VGND VGND VPWR VPWR _10095_ sky130_fd_sc_hd__xnor2_2
X_15323_ net479 _07421_ VGND VGND VPWR VPWR _07422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19091_ net360 net316 _11008_ VGND VGND VPWR VPWR _11063_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18042_ net342 net380 VGND VGND VPWR VPWR _10027_ sky130_fd_sc_hd__nand2_1
X_15254_ _07309_ _07317_ VGND VGND VPWR VPWR _07353_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14205_ _06411_ _06412_ _06413_ _06414_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15185_ net528 net464 VGND VGND VPWR VPWR _07284_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14136_ _06200_ _06201_ _06347_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__a21oi_2
X_19993_ _11807_ VGND VGND VPWR VPWR _11860_ sky130_fd_sc_hd__inv_2
X_14067_ _06279_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__clkbuf_4
X_18944_ _10917_ _10918_ _10905_ VGND VGND VPWR VPWR _10919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18875_ _10848_ _10784_ _10849_ VGND VGND VPWR VPWR _10850_ sky130_fd_sc_hd__a21o_1
XFILLER_0_193_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17826_ _09645_ _09641_ VGND VGND VPWR VPWR _09813_ sky130_fd_sc_hd__or2b_1
XFILLER_0_179_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17757_ _09724_ _09743_ VGND VGND VPWR VPWR _09744_ sky130_fd_sc_hd__xnor2_1
X_14969_ _07106_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16708_ top0.pid_q.curr_int\[13\] _08740_ top0.pid_q.out\[13\] VGND VGND VPWR VPWR
+ _08793_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17688_ net413 net333 net339 net408 VGND VGND VPWR VPWR _09675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19427_ net431 _10333_ _11327_ net442 _11170_ VGND VGND VPWR VPWR _11328_ sky130_fd_sc_hd__a221o_1
X_16639_ _08694_ _08724_ VGND VGND VPWR VPWR _08725_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout19 spi0.data_packed\[14\] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19358_ _11283_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18309_ _10288_ _10290_ VGND VGND VPWR VPWR _10291_ sky130_fd_sc_hd__xor2_2
X_19289_ top0.matmul0.alpha_pass\[11\] _11221_ VGND VGND VPWR VPWR _11232_ sky130_fd_sc_hd__xor2_1
XFILLER_0_143_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21320_ net235 _13124_ VGND VGND VPWR VPWR _13162_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21251_ _12244_ _12669_ VGND VGND VPWR VPWR _13095_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20202_ _12047_ _12048_ _12049_ net269 _12050_ VGND VGND VPWR VPWR _12051_ sky130_fd_sc_hd__a221o_1
X_21182_ net246 _12985_ _13023_ _13024_ _13025_ VGND VGND VPWR VPWR _13026_ sky130_fd_sc_hd__a41o_1
XFILLER_0_25_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20133_ _11426_ net212 VGND VGND VPWR VPWR _11989_ sky130_fd_sc_hd__or2_1
X_25990_ top0.b_in_matmul\[7\] _05192_ _05165_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24941_ _04290_ _04291_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__xnor2_1
X_20064_ net190 _11902_ _11861_ VGND VGND VPWR VPWR _11926_ sky130_fd_sc_hd__o21ai_1
X_24872_ _04073_ _04074_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__nor2_1
X_23823_ _03177_ _03180_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__xnor2_2
X_26611_ clknet_leaf_84_clk_sys _00006_ net633 VGND VGND VPWR VPWR top0.pid_d.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26542_ clknet_leaf_51_clk_sys _00165_ net671 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23754_ _03061_ _03062_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__nor2_4
X_20966_ _12742_ _12810_ _12811_ _12813_ net715 VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22705_ _02222_ _02255_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__xor2_1
X_26473_ clknet_leaf_12_clk_sys _00104_ net603 VGND VGND VPWR VPWR top0.periodTop\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_23685_ _03012_ _03009_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_166_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20897_ _12678_ _12679_ _12685_ VGND VGND VPWR VPWR _12745_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_44_clk_sys clknet_3_7__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_44_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_25424_ top0.matmul0.matmul_stage_inst.mult2\[14\] _04767_ _03146_ VGND VGND VPWR
+ VPWR _04768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22636_ _01063_ _01118_ _01776_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25355_ _04697_ _04699_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__xnor2_1
X_22567_ _02098_ _02121_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24306_ _03660_ _03661_ _03662_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_23_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21518_ net142 VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__inv_2
X_25286_ _04039_ _04562_ _04631_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22498_ net112 _02020_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27025_ clknet_leaf_15_clk_sys _00642_ net617 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_24237_ _03566_ _03583_ _03585_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21449_ net1021 _00994_ _01014_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__or3b_1
XFILLER_0_142_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24168_ _03398_ _03400_ _03410_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23119_ _02485_ _02598_ _02612_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24099_ _03006_ _03185_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__nor2_2
X_16990_ _09043_ _09044_ net547 VGND VGND VPWR VPWR _09045_ sky130_fd_sc_hd__o21a_1
X_15941_ _08033_ _08035_ VGND VGND VPWR VPWR _08036_ sky130_fd_sc_hd__xor2_1
X_18660_ net323 net373 VGND VGND VPWR VPWR _10638_ sky130_fd_sc_hd__nand2_1
X_15872_ net443 _07873_ _07874_ VGND VGND VPWR VPWR _07968_ sky130_fd_sc_hd__a21bo_1
X_17611_ _09594_ _09597_ VGND VGND VPWR VPWR _09598_ sky130_fd_sc_hd__nor2_1
X_14823_ _06982_ _06983_ _07022_ _06952_ VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__o22a_1
XFILLER_0_153_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26809_ clknet_leaf_68_clk_sys _00426_ net662 VGND VGND VPWR VPWR top0.pid_q.prev_int\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_18591_ _10561_ _10569_ VGND VGND VPWR VPWR _10570_ sky130_fd_sc_hd__and2_1
XFILLER_0_192_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17542_ net407 net354 VGND VGND VPWR VPWR _09529_ sky130_fd_sc_hd__nand2_1
X_14754_ _06954_ _06955_ VGND VGND VPWR VPWR _06956_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13705_ _05914_ _05917_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__xnor2_2
X_14685_ net31 _05619_ VGND VGND VPWR VPWR _06889_ sky130_fd_sc_hd__nand2_1
X_17473_ net407 net400 VGND VGND VPWR VPWR _09460_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19212_ _11160_ _11161_ VGND VGND VPWR VPWR _11162_ sky130_fd_sc_hd__nor2_1
X_13636_ _05830_ _05848_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16424_ _08510_ _08512_ VGND VGND VPWR VPWR _08513_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19143_ top0.kid\[6\] _11098_ _11100_ top0.kpd\[6\] VGND VGND VPWR VPWR _11107_ sky130_fd_sc_hd__a22o_1
XFILLER_0_172_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13567_ net43 _05472_ _05678_ _05679_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__a22o_1
X_16355_ _08371_ _08373_ _08369_ VGND VGND VPWR VPWR _08445_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_82_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15306_ net479 _07404_ VGND VGND VPWR VPWR _07405_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16286_ _08362_ _08376_ VGND VGND VPWR VPWR _08377_ sky130_fd_sc_hd__xnor2_2
X_19074_ _11014_ _11039_ _11041_ _11045_ VGND VGND VPWR VPWR _11046_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_48_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13498_ _05509_ _05529_ _05557_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_140_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18025_ net325 net404 VGND VGND VPWR VPWR _10010_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15237_ net541 net462 VGND VGND VPWR VPWR _07336_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15168_ net520 net475 VGND VGND VPWR VPWR _07267_ sky130_fd_sc_hd__nand2_2
X_14119_ _06329_ _06330_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__xor2_2
XFILLER_0_10_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19976_ _11573_ _11510_ _11843_ VGND VGND VPWR VPWR _11844_ sky130_fd_sc_hd__o21ai_1
X_15099_ net525 net471 VGND VGND VPWR VPWR _07198_ sky130_fd_sc_hd__nand2_1
Xfanout209 top0.state\[0\] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18927_ _10766_ _10826_ _10824_ VGND VGND VPWR VPWR _10902_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_201_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18858_ top0.pid_d.curr_int\[10\] VGND VGND VPWR VPWR _10834_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17809_ net409 net404 net335 net337 VGND VGND VPWR VPWR _09796_ sky130_fd_sc_hd__nand4_1
XFILLER_0_94_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18789_ _10731_ _10741_ _10732_ VGND VGND VPWR VPWR _10765_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20820_ _12172_ _12173_ _12243_ VGND VGND VPWR VPWR _12669_ sky130_fd_sc_hd__or3_1
XFILLER_0_148_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20751_ _12589_ _12598_ _12599_ net288 VGND VGND VPWR VPWR _12600_ sky130_fd_sc_hd__a211o_1
XFILLER_0_106_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23470_ _02899_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__clkbuf_1
X_20682_ _12519_ _12520_ _12530_ VGND VGND VPWR VPWR _12531_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22421_ _01899_ _01932_ _01931_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_169_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25140_ _04484_ _04487_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22352_ _01225_ _01328_ _01311_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21303_ _13145_ _13104_ _13103_ VGND VGND VPWR VPWR _13146_ sky130_fd_sc_hd__o21bai_2
X_25071_ _03474_ _03936_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22283_ _01841_ _01842_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_131_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24022_ _03036_ _03037_ _03045_ _03046_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__o22a_1
Xhold230 top0.svm0.tA\[8\] VGND VGND VPWR VPWR net930 sky130_fd_sc_hd__dlygate4sd3_1
X_21234_ _12637_ _13077_ VGND VGND VPWR VPWR _13078_ sky130_fd_sc_hd__nand2_1
Xhold241 top0.pid_d.prev_int\[14\] VGND VGND VPWR VPWR net941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 top0.currT_r\[9\] VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold263 spi0.opcode\[7\] VGND VGND VPWR VPWR net963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _05370_ VGND VGND VPWR VPWR net974 sky130_fd_sc_hd__dlygate4sd3_1
X_21165_ _13008_ _13009_ VGND VGND VPWR VPWR _13010_ sky130_fd_sc_hd__xor2_2
Xhold285 top0.a_in_matmul\[8\] VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold296 top0.cordic0.sin\[12\] VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__dlygate4sd3_1
X_20116_ top0.cordic0.slte0.opA\[14\] _11972_ _11973_ _11971_ VGND VGND VPWR VPWR
+ _00374_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25973_ top0.matmul0.beta_pass\[3\] _05169_ _05179_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__a21o_1
X_21096_ _12941_ VGND VGND VPWR VPWR _12942_ sky130_fd_sc_hd__inv_2
X_24924_ _04273_ _04274_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__xnor2_1
X_20047_ _11896_ _11908_ _11909_ _11886_ _11910_ VGND VGND VPWR VPWR _11911_ sky130_fd_sc_hd__o221a_1
XFILLER_0_176_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24855_ _04107_ _04108_ _04109_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__a21o_1
XFILLER_0_197_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23806_ _03162_ _03163_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__nor2_1
X_24786_ _04136_ _04138_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__xnor2_2
X_21998_ _01555_ _01559_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__xnor2_2
X_23737_ _03063_ _03064_ _03093_ _03094_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__o22a_2
X_26525_ clknet_leaf_60_clk_sys _00148_ net651 VGND VGND VPWR VPWR top0.pid_q.out\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_200_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20949_ _11758_ _12785_ VGND VGND VPWR VPWR _12797_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14470_ _06676_ _06677_ _06553_ _06609_ VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_95_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23668_ _03022_ _03023_ _03024_ _03025_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__o22a_1
X_26456_ clknet_leaf_57_clk_sys _00097_ net664 VGND VGND VPWR VPWR top0.kiq\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13421_ _05633_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25407_ _04712_ _04750_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__xnor2_1
X_22619_ _02168_ _02170_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__nand2_1
X_26387_ clknet_leaf_39_clk_sys _00028_ net682 VGND VGND VPWR VPWR top0.svm0.tC\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_23599_ _02966_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16140_ _08232_ VGND VGND VPWR VPWR _08233_ sky130_fd_sc_hd__inv_2
X_25338_ _04673_ _04682_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__xnor2_2
X_13352_ net43 VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16071_ _08090_ _08149_ _08151_ VGND VGND VPWR VPWR _08164_ sky130_fd_sc_hd__a21bo_1
X_25269_ _04190_ _04131_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__nor2_2
X_13283_ _05495_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15022_ top0.pid_d.state\[0\] top0.pid_d.state\[3\] _07136_ VGND VGND VPWR VPWR _07137_
+ sky130_fd_sc_hd__or3_2
X_27008_ clknet_leaf_26_clk_sys _00625_ net625 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_19830_ _11435_ _11707_ VGND VGND VPWR VPWR _11709_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19761_ _11624_ _11626_ VGND VGND VPWR VPWR _11644_ sky130_fd_sc_hd__nand2_1
X_16973_ _09027_ _09028_ VGND VGND VPWR VPWR _09029_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18712_ net377 _10203_ _09364_ VGND VGND VPWR VPWR _10689_ sky130_fd_sc_hd__o21ai_1
X_15924_ _07933_ _07935_ _08018_ VGND VGND VPWR VPWR _08019_ sky130_fd_sc_hd__a21oi_2
X_19692_ _11416_ _11417_ _11572_ VGND VGND VPWR VPWR _11578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18643_ _10615_ _10620_ VGND VGND VPWR VPWR _10621_ sky130_fd_sc_hd__xnor2_1
X_15855_ _07949_ _07950_ VGND VGND VPWR VPWR _07951_ sky130_fd_sc_hd__xnor2_1
X_14806_ _06935_ _07004_ _07001_ VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18574_ _10484_ _10552_ VGND VGND VPWR VPWR _10553_ sky130_fd_sc_hd__xnor2_2
X_15786_ _07765_ _07770_ VGND VGND VPWR VPWR _07883_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17525_ _09508_ _09509_ _09511_ VGND VGND VPWR VPWR _09512_ sky130_fd_sc_hd__and3_1
X_14737_ _06870_ _06901_ _06866_ VGND VGND VPWR VPWR _06940_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_54_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17456_ _09442_ _09440_ _09373_ VGND VGND VPWR VPWR _09443_ sky130_fd_sc_hd__o21ai_1
X_14668_ _06831_ _06846_ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16407_ net450 net510 VGND VGND VPWR VPWR _08496_ sky130_fd_sc_hd__nand2_1
XFILLER_0_171_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13619_ _05826_ _05831_ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__xnor2_2
X_17387_ _09346_ _09347_ _09345_ VGND VGND VPWR VPWR _09374_ sky130_fd_sc_hd__o21a_1
X_14599_ _06740_ _06745_ _06800_ _06697_ VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__or4b_1
XFILLER_0_172_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19126_ _11095_ VGND VGND VPWR VPWR _11096_ sky130_fd_sc_hd__buf_2
XFILLER_0_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16338_ _08350_ _08360_ _08355_ VGND VGND VPWR VPWR _08428_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_70_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19057_ _11028_ _11029_ VGND VGND VPWR VPWR _11030_ sky130_fd_sc_hd__nor2_1
X_16269_ _08356_ _08359_ VGND VGND VPWR VPWR _08360_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18008_ net421 net313 VGND VGND VPWR VPWR _09993_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19959_ net183 _11808_ _11826_ _11828_ net181 VGND VGND VPWR VPWR _11829_ sky130_fd_sc_hd__a2111o_1
X_22970_ _02478_ _02474_ _02479_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__o21a_1
XFILLER_0_198_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21921_ _01457_ _01482_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__xnor2_2
X_24640_ _03882_ _03897_ _03879_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_171_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21852_ net141 _01412_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20803_ _11608_ _12278_ VGND VGND VPWR VPWR _12652_ sky130_fd_sc_hd__nand2_1
X_24571_ _03924_ _03921_ _03922_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__and3_1
X_21783_ net1031 _01342_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26310_ spi0.data_packed\[53\] spi0.data_packed\[54\] net700 VGND VGND VPWR VPWR
+ _05387_ sky130_fd_sc_hd__mux2_1
X_23522_ top0.a_in_matmul\[1\] top0.matmul0.a\[1\] _02926_ VGND VGND VPWR VPWR _02927_
+ sky130_fd_sc_hd__mux2_1
X_20734_ _12580_ _12582_ VGND VGND VPWR VPWR _12583_ sky130_fd_sc_hd__xnor2_2
X_27290_ clknet_3_3__leaf_clk_mosi _00904_ VGND VGND VPWR VPWR spi0.data_packed\[76\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26241_ _05352_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23453_ _02879_ _02877_ _02887_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__o21a_1
XFILLER_0_175_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20665_ _12503_ _12512_ VGND VGND VPWR VPWR _12514_ sky130_fd_sc_hd__nor2_1
XFILLER_0_190_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22404_ net134 _01957_ _01961_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26172_ spi0.data_packed\[6\] spi0.data_packed\[7\] _05303_ VGND VGND VPWR VPWR _05310_
+ sky130_fd_sc_hd__and3_1
X_23384_ _02796_ _02797_ _02807_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__or3_1
X_20596_ _12332_ _12444_ VGND VGND VPWR VPWR _12445_ sky130_fd_sc_hd__xnor2_2
X_25123_ _04471_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22335_ _01742_ _01893_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__nand2_1
X_25054_ _04251_ _04325_ _04334_ _04399_ _04330_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22266_ _01824_ _01822_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__nand2_1
X_24005_ _03069_ _03071_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__or2_2
X_21217_ _12646_ _12577_ VGND VGND VPWR VPWR _13061_ sky130_fd_sc_hd__nand2_1
X_22197_ net109 _01143_ _01757_ _01291_ _01116_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__a221o_2
XFILLER_0_40_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21148_ _12987_ _12992_ VGND VGND VPWR VPWR _12993_ sky130_fd_sc_hd__xnor2_1
Xfanout540 net541 VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__clkbuf_4
Xfanout551 net552 VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__buf_2
Xfanout562 net563 VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__clkbuf_4
X_13970_ _05541_ _05608_ _05609_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__or3_1
Xfanout573 top0.matmul0.matmul_stage_inst.state\[1\] VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__clkbuf_4
X_21079_ _12924_ _12851_ VGND VGND VPWR VPWR _12925_ sky130_fd_sc_hd__or2b_1
X_25956_ top0.matmul0.op_in\[1\] _12015_ _05165_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__mux2_1
Xfanout584 net585 VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__buf_2
Xfanout595 net596 VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__clkbuf_4
X_24907_ _04039_ _04067_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_100_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25887_ top0.matmul0.alpha_pass\[10\] net429 VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15640_ _07732_ _07737_ VGND VGND VPWR VPWR _07738_ sky130_fd_sc_hd__xnor2_2
X_24838_ _03090_ _03091_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__nor2_4
XFILLER_0_197_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15571_ _07665_ _07669_ VGND VGND VPWR VPWR _07670_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24769_ _04120_ _04121_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17310_ _09303_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__clkbuf_1
X_14522_ _06629_ _06632_ _06728_ VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__o21ai_2
X_26508_ clknet_leaf_77_clk_sys _00131_ net631 VGND VGND VPWR VPWR top0.pid_d.prev_int\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18290_ net331 net378 VGND VGND VPWR VPWR _10272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17241_ top0.pid_q.curr_int\[14\] top0.pid_q.prev_int\[14\] VGND VGND VPWR VPWR _09245_
+ sky130_fd_sc_hd__nor2_1
X_14453_ _06614_ _06660_ VGND VGND VPWR VPWR _06661_ sky130_fd_sc_hd__xnor2_4
X_26439_ clknet_leaf_80_clk_sys _00080_ net634 VGND VGND VPWR VPWR top0.kid\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13404_ top0.matmul0.beta_pass\[12\] _05435_ _05470_ _05464_ top0.c_out_calc\[12\]
+ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_126_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14384_ _06582_ _06592_ VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17172_ top0.pid_q.prev_int\[5\] _09172_ _09177_ top0.pid_q.prev_int\[6\] VGND VGND
+ VPWR VPWR _09184_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13335_ _05535_ _05547_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__xnor2_2
X_16123_ _08214_ _08215_ VGND VGND VPWR VPWR _08216_ sky130_fd_sc_hd__or2b_1
XFILLER_0_49_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13266_ top0.matmul0.beta_pass\[3\] _05434_ _05469_ _05463_ top0.c_out_calc\[3\]
+ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__a32oi_4
X_16054_ _08140_ _08147_ VGND VGND VPWR VPWR _08148_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15005_ spi0.data_packed\[8\] top0.periodTop\[8\] _07125_ VGND VGND VPWR VPWR _07128_
+ sky130_fd_sc_hd__mux2_1
X_13197_ top0.pid_d.iterate_enable VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19813_ _11676_ _11677_ _11513_ VGND VGND VPWR VPWR _11693_ sky130_fd_sc_hd__o21a_1
X_19744_ _11435_ _11621_ _11624_ _11626_ _11608_ VGND VGND VPWR VPWR _11628_ sky130_fd_sc_hd__a41oi_1
X_16956_ net429 _09012_ VGND VGND VPWR VPWR _09013_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15907_ net496 net492 VGND VGND VPWR VPWR _08002_ sky130_fd_sc_hd__or2_1
X_19675_ net128 net123 net121 net116 net199 net193 VGND VGND VPWR VPWR _11562_ sky130_fd_sc_hd__mux4_1
XFILLER_0_194_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16887_ top0.currT_r\[5\] _08948_ VGND VGND VPWR VPWR _08949_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18626_ _10439_ _10602_ _10603_ _10504_ VGND VGND VPWR VPWR _10604_ sky130_fd_sc_hd__o22a_1
XFILLER_0_154_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15838_ net448 net532 VGND VGND VPWR VPWR _07934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18557_ _10519_ _10535_ VGND VGND VPWR VPWR _10536_ sky130_fd_sc_hd__xnor2_4
X_15769_ _07864_ _07865_ VGND VGND VPWR VPWR _07866_ sky130_fd_sc_hd__nor2_1
X_17508_ net388 net357 VGND VGND VPWR VPWR _09495_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18488_ _10466_ _10467_ VGND VGND VPWR VPWR _10468_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17439_ _09418_ _09425_ VGND VGND VPWR VPWR _09426_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_14 _12739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_131_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_25 net1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_36 _10561_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 net687 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20450_ _12295_ _12298_ VGND VGND VPWR VPWR _12299_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19109_ top0.pid_d.out\[15\] _09339_ _11080_ _05443_ net435 VGND VGND VPWR VPWR _11081_
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_166_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20381_ _12228_ _12229_ VGND VGND VPWR VPWR _12230_ sky130_fd_sc_hd__and2_1
XFILLER_0_179_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22120_ _01667_ _01680_ _01681_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__or3b_1
XFILLER_0_42_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22051_ _01180_ _01181_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21002_ _12208_ _12848_ VGND VGND VPWR VPWR _12849_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25810_ _05035_ _05033_ _05034_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__and3_1
XFILLER_0_195_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26790_ clknet_leaf_1_clk_sys _00407_ net582 VGND VGND VPWR VPWR top0.cordic0.sin\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22953_ _02465_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__clkbuf_1
X_25741_ _04991_ _04912_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__and2b_1
XFILLER_0_69_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21904_ net151 net130 _01462_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__a21o_1
X_22884_ _02317_ top0.svm0.tB\[13\] _02401_ _02402_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__o22a_1
X_25672_ _04942_ _04943_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24623_ _03972_ _03973_ _03047_ _03827_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__a211o_1
X_21835_ _01390_ _01391_ _01396_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24554_ _03185_ _03908_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21766_ net133 net1031 VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__xor2_4
X_20717_ _12564_ _12565_ VGND VGND VPWR VPWR _12566_ sky130_fd_sc_hd__or2_1
X_23505_ top0.cordic0.cos\[7\] top0.matmul0.cos\[7\] _02915_ VGND VGND VPWR VPWR _02918_
+ sky130_fd_sc_hd__mux2_1
X_24485_ _03735_ _03748_ _03736_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__o21bai_1
X_27273_ clknet_3_7__leaf_clk_mosi _00887_ VGND VGND VPWR VPWR spi0.data_packed\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_21697_ net129 net113 VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__xnor2_4
X_23436_ _11649_ _02872_ _11954_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__a21o_1
X_26224_ spi0.data_packed\[10\] spi0.data_packed\[11\] net695 VGND VGND VPWR VPWR
+ _05344_ sky130_fd_sc_hd__mux2_1
X_20648_ net274 _12494_ _12496_ _12493_ VGND VGND VPWR VPWR _12497_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26155_ spi0.data_packed\[4\] _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23367_ _02807_ _02808_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__xnor2_2
X_20579_ _12056_ _12254_ VGND VGND VPWR VPWR _12428_ sky130_fd_sc_hd__xnor2_2
X_25106_ _04419_ _04454_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__xnor2_2
X_22318_ _01806_ _01874_ _01876_ _01877_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__a211o_1
X_26086_ top0.a_in_matmul\[13\] _05266_ _05164_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23298_ _02725_ _02734_ _01102_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__o21a_1
X_25037_ _04385_ _04386_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__and2_1
X_22249_ net210 _01738_ _01807_ _01808_ _01809_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__a32o_1
X_16810_ top0.pid_q.mult0.a\[14\] _08855_ _08858_ net803 _08878_ VGND VGND VPWR VPWR
+ _00163_ sky130_fd_sc_hd__a221o_1
X_17790_ net404 net336 VGND VGND VPWR VPWR _09777_ sky130_fd_sc_hd__nand2_1
X_26988_ clknet_leaf_28_clk_sys _00605_ net622 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout370 top0.pid_d.mult0.a\[14\] VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkbuf_4
Xfanout381 net382 VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__clkbuf_4
X_16741_ net445 _08703_ _08821_ _08822_ _08824_ VGND VGND VPWR VPWR _08825_ sky130_fd_sc_hd__a32o_1
Xfanout392 net394 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkbuf_4
X_13953_ _06163_ _06164_ _06165_ _06138_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__and4_1
X_25939_ _05146_ _05150_ _05151_ _02282_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__a31o_1
X_19460_ top0.pid_d.curr_int\[9\] _11290_ _11293_ _11356_ VGND VGND VPWR VPWR _00335_
+ sky130_fd_sc_hd__a22o_1
X_16672_ _08220_ _08756_ VGND VGND VPWR VPWR _08757_ sky130_fd_sc_hd__xnor2_1
X_13884_ _05565_ _05543_ _05545_ VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__or3_1
XFILLER_0_115_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18411_ _10381_ _10390_ VGND VGND VPWR VPWR _10392_ sky130_fd_sc_hd__or2_1
XFILLER_0_202_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15623_ net469 net518 VGND VGND VPWR VPWR _07721_ sky130_fd_sc_hd__nand2_1
X_19391_ top0.pid_d.curr_int\[0\] _11290_ _11293_ _11296_ VGND VGND VPWR VPWR _00326_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18342_ _10322_ _10323_ VGND VGND VPWR VPWR _10324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15554_ _07651_ _07652_ VGND VGND VPWR VPWR _07653_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14505_ _06706_ _06711_ VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_92_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_92_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_185_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18273_ net318 net365 VGND VGND VPWR VPWR _10255_ sky130_fd_sc_hd__and2_2
X_15485_ _07581_ _07583_ VGND VGND VPWR VPWR _07584_ sky130_fd_sc_hd__xnor2_1
X_17224_ top0.pid_q.curr_int\[12\] top0.pid_q.prev_int\[12\] _09225_ VGND VGND VPWR
+ VPWR _09230_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14436_ net23 _05586_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17155_ net543 _08075_ _09169_ VGND VGND VPWR VPWR _09170_ sky130_fd_sc_hd__a21o_1
X_14367_ _06494_ _06499_ _06575_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_25_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16106_ _08097_ _08104_ _08099_ VGND VGND VPWR VPWR _08199_ sky130_fd_sc_hd__o21ba_1
X_13318_ top0.matmul0.alpha_pass\[6\] _05434_ _05467_ VGND VGND VPWR VPWR _05531_
+ sky130_fd_sc_hd__and3_2
X_14298_ _06427_ _06428_ _06506_ _06507_ VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__o31ai_4
X_17086_ top0.pid_q.prev_error\[1\] _09115_ _09119_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16037_ _08033_ _08035_ _08031_ VGND VGND VPWR VPWR _08131_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_110_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13249_ net173 top0.svm0.state\[1\] top0.svm0.state\[0\] VGND VGND VPWR VPWR _05462_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_161_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17988_ _09885_ _09883_ _09973_ VGND VGND VPWR VPWR _09974_ sky130_fd_sc_hd__o21ai_2
X_19727_ _11610_ VGND VGND VPWR VPWR _11611_ sky130_fd_sc_hd__inv_2
X_16939_ top0.currT_r\[8\] _08984_ _08996_ VGND VGND VPWR VPWR _08997_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19658_ _11544_ _11545_ VGND VGND VPWR VPWR _11546_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18609_ _10443_ _10504_ _10586_ _10587_ VGND VGND VPWR VPWR _10588_ sky130_fd_sc_hd__a31o_1
XFILLER_0_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19589_ top0.cordic0.slte0.opB\[7\] top0.cordic0.slte0.opA\[7\] VGND VGND VPWR VPWR
+ _11478_ sky130_fd_sc_hd__xor2_1
X_21620_ _01180_ _01181_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21551_ net104 _01112_ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_145_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20502_ _11407_ _12065_ _12156_ net296 VGND VGND VPWR VPWR _12351_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24270_ _03293_ _03294_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__nand2_2
XFILLER_0_74_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21482_ net231 _01045_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23221_ _02670_ _02671_ _02660_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20433_ _12276_ _12281_ VGND VGND VPWR VPWR _12282_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23152_ _02637_ _02638_ _07117_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__a21oi_1
X_20364_ net296 net277 net269 VGND VGND VPWR VPWR _12213_ sky130_fd_sc_hd__or3b_1
XFILLER_0_113_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22103_ _01663_ _01660_ _01664_ _01653_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__a22oi_1
X_23083_ _02581_ _02582_ _02583_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__o21ai_1
X_20295_ net264 net261 VGND VGND VPWR VPWR _12144_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22034_ _01265_ _01279_ _01278_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__o21bai_2
X_26911_ clknet_leaf_109_clk_sys _00528_ net579 VGND VGND VPWR VPWR top0.matmul0.sin\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_26842_ clknet_leaf_44_clk_sys _00459_ net681 VGND VGND VPWR VPWR top0.svm0.delta\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_26773_ clknet_leaf_6_clk_sys _00390_ net590 VGND VGND VPWR VPWR top0.cordic0.cos\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_177_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23985_ _03024_ _03025_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__nor2_4
X_25724_ net856 _04964_ _04913_ _04980_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__a22o_1
X_22936_ _02449_ _02450_ _02347_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25655_ net799 _04925_ _04930_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_79_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22867_ _02332_ top0.svm0.tB\[4\] _02384_ top0.svm0.tB\[3\] _02385_ VGND VGND VPWR
+ VPWR _02386_ sky130_fd_sc_hd__o221a_1
XFILLER_0_167_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24606_ top0.matmul0.matmul_stage_inst.mult2\[3\] _03960_ _03642_ VGND VGND VPWR
+ VPWR _03961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21818_ net135 net121 VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22798_ _02317_ top0.svm0.tA\[13\] VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__and2_1
X_25586_ top0.matmul0.a\[15\] top0.matmul0.matmul_stage_inst.e\[15\] _04878_ VGND
+ VGND VPWR VPWR _04881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24537_ _03790_ _03792_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__and2_1
X_21749_ _01310_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_164_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27256_ clknet_3_2__leaf_clk_mosi _00870_ VGND VGND VPWR VPWR spi0.data_packed\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_15270_ net525 net479 VGND VGND VPWR VPWR _07369_ sky130_fd_sc_hd__nand2_1
X_24468_ _03690_ _03822_ _03823_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14221_ _06427_ _06428_ _06429_ _06430_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__o22ai_2
X_26207_ _05335_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__clkbuf_1
X_23419_ _11514_ _02856_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24399_ _03658_ _03755_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__xnor2_1
X_27187_ clknet_leaf_56_clk_sys _00801_ net666 VGND VGND VPWR VPWR top0.currT_r\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_46_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14152_ _06360_ _06361_ _06362_ _06363_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__o22a_1
XFILLER_0_151_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26138_ spi0.data_packed\[0\] _05283_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14083_ _06285_ _06294_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__xnor2_4
X_18960_ _10805_ _10875_ _10887_ _10723_ VGND VGND VPWR VPWR _10934_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26069_ top0.matmul0.alpha_pass\[9\] _05237_ _05253_ VGND VGND VPWR VPWR _05254_
+ sky130_fd_sc_hd__a21o_1
X_17911_ top0.pid_d.out\[0\] _07138_ _09897_ net434 VGND VGND VPWR VPWR _09898_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_39_clk_sys clknet_3_7__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_39_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18891_ net374 net312 VGND VGND VPWR VPWR _10866_ sky130_fd_sc_hd__nand2_1
X_17842_ net322 net417 VGND VGND VPWR VPWR _09829_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17773_ _09758_ _09759_ VGND VGND VPWR VPWR _09760_ sky130_fd_sc_hd__xnor2_1
X_14985_ _07116_ VGND VGND VPWR VPWR _07117_ sky130_fd_sc_hd__buf_2
XFILLER_0_195_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19512_ _11401_ _11399_ _11400_ VGND VGND VPWR VPWR _11403_ sky130_fd_sc_hd__nand3_1
X_16724_ _08769_ _08774_ _08807_ VGND VGND VPWR VPWR _08808_ sky130_fd_sc_hd__o21a_1
X_13936_ net60 _05726_ _05727_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19443_ _11340_ VGND VGND VPWR VPWR _11341_ sky130_fd_sc_hd__buf_2
X_16655_ top0.pid_q.curr_int\[13\] _08740_ VGND VGND VPWR VPWR _08741_ sky130_fd_sc_hd__xor2_1
X_13867_ _05922_ _05949_ _06075_ _06077_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__a31o_1
XFILLER_0_201_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15606_ _07704_ VGND VGND VPWR VPWR _07705_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19374_ net880 _11285_ _11288_ top0.pid_d.curr_error\[7\] VGND VGND VPWR VPWR _00317_
+ sky130_fd_sc_hd__a22o_1
X_16586_ _08668_ _08672_ VGND VGND VPWR VPWR _08673_ sky130_fd_sc_hd__xnor2_1
X_13798_ _06005_ _06006_ _05517_ VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__o21a_1
X_18325_ _10215_ _10218_ _10216_ VGND VGND VPWR VPWR _10307_ sky130_fd_sc_hd__a21bo_1
X_15537_ _07630_ _07635_ VGND VGND VPWR VPWR _07636_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18256_ _10135_ _10145_ _10144_ VGND VGND VPWR VPWR _10239_ sky130_fd_sc_hd__a21o_1
X_15468_ net531 net460 VGND VGND VPWR VPWR _07567_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17207_ top0.pid_q.prev_int\[10\] VGND VGND VPWR VPWR _09215_ sky130_fd_sc_hd__inv_2
X_14419_ _06623_ _06626_ VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__xnor2_2
X_18187_ net334 net378 VGND VGND VPWR VPWR _10170_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15399_ net541 _07484_ net472 VGND VGND VPWR VPWR _07498_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17138_ _09147_ _09148_ _09153_ VGND VGND VPWR VPWR _09154_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17069_ top0.pid_q.curr_error\[11\] _09100_ _09102_ _09036_ VGND VGND VPWR VPWR _00192_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20080_ top0.cordic0.slte0.opA\[10\] _11932_ _11931_ VGND VGND VPWR VPWR _11941_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_176_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_191_Right_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23770_ _03126_ _03127_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__nor2_1
X_20982_ _12826_ _12827_ _12828_ VGND VGND VPWR VPWR _12829_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22721_ _02237_ _02240_ _02255_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25440_ _04562_ _04631_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22652_ _02202_ _02204_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__and2_1
XFILLER_0_178_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21603_ _01163_ _01164_ net90 VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__mux2_2
X_25371_ _04668_ _04714_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22583_ _02079_ _02086_ _02124_ _02136_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27110_ clknet_leaf_11_clk_sys _00016_ net601 VGND VGND VPWR VPWR top0.matmul0.state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_24322_ _03677_ _03166_ _03678_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__o21ai_4
X_21534_ net146 _01090_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24253_ _03511_ _03516_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__xor2_1
X_27041_ clknet_leaf_8_clk_sys _00658_ net597 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_21465_ _12769_ _12761_ _12820_ _11759_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23204_ _02652_ _02655_ _11420_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__mux2_1
X_20416_ net298 net294 VGND VGND VPWR VPWR _12265_ sky130_fd_sc_hd__or2b_1
XFILLER_0_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24184_ _03015_ _03016_ _03076_ _03077_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__o22a_1
XFILLER_0_102_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21396_ _00954_ _00956_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23135_ top0.svm0.delta\[11\] _02622_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__or2_1
X_20347_ _12186_ _12191_ _12193_ _12195_ VGND VGND VPWR VPWR _12196_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_109_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_40_clk_sys clknet_3_7__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_40_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_23066_ net46 _02540_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20278_ _11672_ _12126_ VGND VGND VPWR VPWR _12127_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_101_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22017_ net153 net135 VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__xor2_1
XFILLER_0_41_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26825_ clknet_leaf_46_clk_sys _00442_ net680 VGND VGND VPWR VPWR top0.svm0.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_14770_ net857 _06279_ _06971_ _05465_ VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__a22o_1
X_26756_ clknet_leaf_5_clk_sys _00373_ net590 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23968_ _03325_ _03254_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__nor2_2
X_13721_ _05932_ _05933_ net54 _05495_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__o211a_1
X_25707_ top0.matmul0.sin\[1\] top0.matmul0.sin\[0\] top0.matmul0.sin\[2\] net72 VGND
+ VGND VPWR VPWR _04969_ sky130_fd_sc_hd__o31a_1
XFILLER_0_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22919_ _02298_ net555 _02297_ _02435_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__a31o_1
X_26687_ clknet_leaf_83_clk_sys _00304_ net646 VGND VGND VPWR VPWR top0.pid_d.curr_error\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_23899_ _03250_ _03113_ VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__nor2_2
XFILLER_0_195_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16440_ _08523_ _08528_ VGND VGND VPWR VPWR _08529_ sky130_fd_sc_hd__and2b_1
X_13652_ _05810_ _05864_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25638_ top0.matmul0.sin\[1\] top0.matmul0.sin\[0\] top0.matmul0.sin\[2\] top0.matmul0.sin\[3\]
+ _04884_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__o311a_1
XFILLER_0_112_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16371_ _08339_ _08346_ _08460_ VGND VGND VPWR VPWR _08461_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13583_ _05795_ _05789_ _05793_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__o21a_1
XFILLER_0_137_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25569_ top0.matmul0.a\[7\] top0.matmul0.matmul_stage_inst.e\[7\] _04867_ VGND VGND
+ VPWR VPWR _04872_ sky130_fd_sc_hd__mux2_1
X_18110_ _10092_ _10093_ VGND VGND VPWR VPWR _10094_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15322_ net1026 _07404_ VGND VGND VPWR VPWR _07421_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19090_ _11052_ _11061_ VGND VGND VPWR VPWR _11062_ sky130_fd_sc_hd__xor2_1
XFILLER_0_136_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18041_ top0.pid_d.mult0.b\[5\] net383 VGND VGND VPWR VPWR _10026_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27239_ clknet_3_7__leaf_clk_mosi _00853_ VGND VGND VPWR VPWR spi0.data_packed\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_15253_ _07332_ _07349_ _07330_ VGND VGND VPWR VPWR _07352_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_163_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14204_ _06411_ _06412_ _06413_ _06414_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__or4_4
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15184_ net531 net462 VGND VGND VPWR VPWR _07283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14135_ _06200_ _06201_ _06198_ VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19992_ _11856_ _11858_ _11859_ net981 VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14066_ _06277_ _06278_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__nand2_4
XFILLER_0_39_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18943_ _10828_ _10829_ net435 VGND VGND VPWR VPWR _10918_ sky130_fd_sc_hd__nor3b_1
X_18874_ _10848_ _10784_ _10769_ VGND VGND VPWR VPWR _10849_ sky130_fd_sc_hd__o21ba_1
X_17825_ _09810_ _09635_ _09811_ VGND VGND VPWR VPWR _09812_ sky130_fd_sc_hd__o21a_1
Xhold1 spi0.cs_sync\[0\] VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17756_ _09726_ _09737_ VGND VGND VPWR VPWR _09743_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_178_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14968_ spi0.data_packed\[26\] top0.kiq\[10\] _07097_ VGND VGND VPWR VPWR _07106_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16707_ top0.pid_q.out\[14\] _07704_ VGND VGND VPWR VPWR _08792_ sky130_fd_sc_hd__nor2_1
X_13919_ _05725_ _05728_ top0.periodTop_r\[0\] _06131_ VGND VGND VPWR VPWR _06132_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17687_ _09670_ _09673_ VGND VGND VPWR VPWR _09674_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14899_ spi0.data_packed\[57\] top0.kpq\[9\] _07064_ VGND VGND VPWR VPWR _07070_
+ sky130_fd_sc_hd__mux2_1
X_19426_ _11325_ _11326_ VGND VGND VPWR VPWR _11327_ sky130_fd_sc_hd__xnor2_1
X_16638_ _08716_ _08723_ VGND VGND VPWR VPWR _08724_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19357_ _05449_ _11282_ VGND VGND VPWR VPWR _11283_ sky130_fd_sc_hd__and2_1
X_16569_ _08571_ _08574_ _08655_ _07213_ net459 VGND VGND VPWR VPWR _08656_ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18308_ net364 _10289_ VGND VGND VPWR VPWR _10290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19288_ net437 _11229_ _11230_ VGND VGND VPWR VPWR _11231_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18239_ _10200_ _10221_ VGND VGND VPWR VPWR _10222_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21250_ _13079_ _13092_ _13093_ _12666_ VGND VGND VPWR VPWR _13094_ sky130_fd_sc_hd__a211oi_2
X_20201_ net276 net269 VGND VGND VPWR VPWR _12050_ sky130_fd_sc_hd__nor2_1
X_21181_ _12985_ _13019_ VGND VGND VPWR VPWR _13025_ sky130_fd_sc_hd__and2b_1
XFILLER_0_13_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20132_ _11986_ _11987_ _11936_ VGND VGND VPWR VPWR _11988_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24940_ _03254_ _03900_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__nor2_1
X_20063_ top0.cordic0.slte0.opA\[9\] _11918_ _11920_ VGND VGND VPWR VPWR _11925_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_110_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24871_ _04073_ _04074_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__and2_1
X_26610_ clknet_leaf_80_clk_sys _00005_ net633 VGND VGND VPWR VPWR top0.pid_d.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_197_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23822_ _03178_ _03179_ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26541_ clknet_leaf_60_clk_sys _00164_ net653 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[15\]
+ sky130_fd_sc_hd__dfrtp_2
X_23753_ _03087_ _03100_ _03110_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__o21bai_1
X_20965_ _12812_ VGND VGND VPWR VPWR _12813_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_200_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22704_ _02250_ _02253_ _02254_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__o21ai_2
X_26472_ clknet_leaf_12_clk_sys _00103_ net603 VGND VGND VPWR VPWR top0.periodTop\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23684_ _03038_ _03039_ _03041_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__o21a_2
X_20896_ _12743_ VGND VGND VPWR VPWR _12744_ sky130_fd_sc_hd__buf_1
XFILLER_0_193_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_156_Left_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25423_ _04754_ _04766_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__xnor2_1
X_22635_ _01221_ _02187_ _01166_ _01118_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__a211o_1
XFILLER_0_192_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25354_ _04522_ _04698_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22566_ _02119_ _02120_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24305_ _03291_ _03229_ _03230_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__and3b_1
X_21517_ net139 net131 VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__nor2_2
XFILLER_0_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25285_ _04371_ _03056_ _03363_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22497_ _02017_ _02022_ _02052_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__a21o_1
X_27024_ clknet_leaf_18_clk_sys _00641_ net612 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24236_ _03584_ _03589_ _03590_ _03593_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__a22o_1
X_21448_ _01002_ _01013_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_160_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24167_ _03478_ _03489_ _03524_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__a21o_1
X_21379_ _00940_ _00946_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_165_Left_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23118_ _02483_ _02612_ _02596_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__o21ai_1
X_24098_ _03379_ _03383_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__xnor2_4
X_23049_ net36 _02542_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__nor2_1
X_15940_ _07948_ _07950_ _08034_ VGND VGND VPWR VPWR _08035_ sky130_fd_sc_hd__a21oi_2
X_15871_ _07828_ _07830_ _07966_ VGND VGND VPWR VPWR _07967_ sky130_fd_sc_hd__a21oi_1
X_17610_ _09555_ _09596_ VGND VGND VPWR VPWR _09597_ sky130_fd_sc_hd__xnor2_1
X_14822_ _06981_ _06984_ VGND VGND VPWR VPWR _07022_ sky130_fd_sc_hd__nor2_1
XFILLER_0_192_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26808_ clknet_leaf_68_clk_sys _00425_ net662 VGND VGND VPWR VPWR top0.pid_q.prev_int\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18590_ _10562_ _10568_ VGND VGND VPWR VPWR _10569_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17541_ _09521_ _09527_ VGND VGND VPWR VPWR _09528_ sky130_fd_sc_hd__nor2_1
X_14753_ net25 _05726_ _05727_ VGND VGND VPWR VPWR _06955_ sky130_fd_sc_hd__and3_2
X_26739_ clknet_leaf_96_clk_sys _00356_ net587 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[14\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_58_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_174_Left_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13704_ _05915_ _05916_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__or2_1
X_17472_ _09351_ net390 VGND VGND VPWR VPWR _09459_ sky130_fd_sc_hd__nand2_1
X_14684_ net37 _06351_ VGND VGND VPWR VPWR _06888_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19211_ top0.matmul0.alpha_pass\[4\] _11150_ VGND VGND VPWR VPWR _11161_ sky130_fd_sc_hd__and2_1
X_16423_ net498 _08511_ VGND VGND VPWR VPWR _08512_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13635_ _05832_ _05844_ _05847_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__a21oi_2
X_19142_ net405 _11096_ _11106_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__a21o_1
X_16354_ _08364_ _08375_ _08443_ VGND VGND VPWR VPWR _08444_ sky130_fd_sc_hd__o21a_1
X_13566_ _05696_ _05698_ _05778_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__a21bo_1
X_15305_ net533 _07403_ VGND VGND VPWR VPWR _07404_ sky130_fd_sc_hd__and2_1
X_19073_ _11043_ _11044_ _10999_ VGND VGND VPWR VPWR _11045_ sky130_fd_sc_hd__mux2_1
X_16285_ _08364_ _08375_ VGND VGND VPWR VPWR _08376_ sky130_fd_sc_hd__xor2_1
X_13497_ _05693_ _05709_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18024_ _09918_ _09929_ _10008_ VGND VGND VPWR VPWR _10009_ sky130_fd_sc_hd__o21ai_2
X_15236_ net537 net464 VGND VGND VPWR VPWR _07335_ sky130_fd_sc_hd__nand2_2
XFILLER_0_2_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_183_Left_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15167_ _07201_ _07264_ _07265_ VGND VGND VPWR VPWR _07266_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_50_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14118_ net30 _05520_ _05521_ VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__and3_2
X_19975_ _11484_ _11504_ _11509_ net189 _11410_ VGND VGND VPWR VPWR _11843_ sky130_fd_sc_hd__a2111o_1
X_15098_ net528 net470 VGND VGND VPWR VPWR _07197_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14049_ _06164_ _06165_ _06161_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__a21oi_1
X_18926_ _10900_ VGND VGND VPWR VPWR _10901_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18857_ top0.pid_d.out\[11\] _07138_ VGND VGND VPWR VPWR _10833_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17808_ _09791_ _09794_ VGND VGND VPWR VPWR _09795_ sky130_fd_sc_hd__xnor2_2
X_18788_ _10684_ _10752_ _10751_ VGND VGND VPWR VPWR _10764_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_192_Left_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17739_ _09701_ _09725_ VGND VGND VPWR VPWR _09726_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_173_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20750_ _12589_ _12598_ net258 VGND VGND VPWR VPWR _12599_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19409_ top0.pid_d.curr_int\[3\] top0.pid_d.prev_int\[3\] VGND VGND VPWR VPWR _11312_
+ sky130_fd_sc_hd__xnor2_1
X_20681_ net274 _12524_ _12528_ _12529_ VGND VGND VPWR VPWR _12530_ sky130_fd_sc_hd__a211o_1
XFILLER_0_175_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22420_ _01953_ _01977_ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22351_ _01225_ _01327_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21302_ _13016_ VGND VGND VPWR VPWR _13145_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25070_ _04410_ _04418_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__xnor2_2
X_22282_ _01225_ _01328_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_198_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24021_ _02982_ _03161_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__nor2_2
XFILLER_0_130_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21233_ _12605_ _13076_ VGND VGND VPWR VPWR _13077_ sky130_fd_sc_hd__xnor2_1
Xhold220 top0.cordic0.sin\[5\] VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 top0.pid_d.curr_error\[10\] VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 spi0.data_packed\[43\] VGND VGND VPWR VPWR net942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 spi0.data_packed\[38\] VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 top0.pid_d.prev_int\[4\] VGND VGND VPWR VPWR net964 sky130_fd_sc_hd__dlygate4sd3_1
X_21164_ _12939_ _12951_ _12938_ VGND VGND VPWR VPWR _13009_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold275 spi0.data_packed\[35\] VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 net1 VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__clkbuf_2
Xhold286 top0.pid_d.curr_error\[2\] VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 top0.matmul0.state\[0\] VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20115_ top0.cordic0.slte0.opA\[14\] _11857_ VGND VGND VPWR VPWR _11973_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21095_ _12806_ _12878_ VGND VGND VPWR VPWR _12941_ sky130_fd_sc_hd__or2_1
X_25972_ top0.pid_q.out\[3\] _12032_ _05014_ spi0.data_packed\[51\] VGND VGND VPWR
+ VPWR _05179_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24923_ _03496_ _04182_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__nor2_1
X_20046_ top0.cordic0.slte0.opA\[7\] _11895_ VGND VGND VPWR VPWR _11910_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24854_ _04100_ _04204_ _04205_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__a21o_1
XFILLER_0_197_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23805_ net568 top0.matmul0.matmul_stage_inst.b\[13\] top0.matmul0.matmul_stage_inst.a\[13\]
+ net564 VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__a22o_2
XFILLER_0_198_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24785_ _04137_ _03971_ _03970_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__a21bo_1
X_21997_ _01557_ _01558_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26524_ clknet_leaf_66_clk_sys _00147_ net660 VGND VGND VPWR VPWR top0.pid_q.out\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_23736_ net567 net560 top0.matmul0.matmul_stage_inst.e\[10\] VGND VGND VPWR VPWR
+ _03094_ sky130_fd_sc_hd__o21a_2
X_20948_ _11758_ _12785_ VGND VGND VPWR VPWR _12796_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26455_ clknet_leaf_57_clk_sys _00096_ net642 VGND VGND VPWR VPWR top0.kiq\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23667_ net570 top0.matmul0.matmul_stage_inst.b\[9\] top0.matmul0.matmul_stage_inst.a\[9\]
+ net566 VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__a22o_4
X_20879_ _12722_ _12723_ _12726_ VGND VGND VPWR VPWR _12728_ sky130_fd_sc_hd__a21o_1
X_25406_ _04382_ _04749_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__xnor2_2
X_13420_ _05630_ _05631_ _05632_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22618_ _02171_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__inv_2
X_26386_ clknet_leaf_41_clk_sys _00027_ net682 VGND VGND VPWR VPWR top0.svm0.tC\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_193_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23598_ top0.matmul0.alpha_pass\[6\] _09284_ net559 VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25337_ _04680_ _04681_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__and2b_1
X_13351_ _05560_ _05563_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22549_ net119 _01069_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16070_ _08088_ _08161_ _08162_ VGND VGND VPWR VPWR _08163_ sky130_fd_sc_hd__a21oi_1
X_25268_ _04097_ _04288_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__nor2_2
X_13282_ _05493_ _05494_ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__nor2_1
X_27007_ clknet_leaf_26_clk_sys _00624_ net627 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_15021_ net431 net441 VGND VGND VPWR VPWR _07136_ sky130_fd_sc_hd__or2_2
X_24219_ _03114_ _03161_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25199_ _04477_ _04478_ _04545_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16972_ top0.pid_q.prev_error\[11\] top0.pid_q.curr_error\[11\] VGND VGND VPWR VPWR
+ _09028_ sky130_fd_sc_hd__xor2_1
X_19760_ _11640_ _11642_ VGND VGND VPWR VPWR _11643_ sky130_fd_sc_hd__xnor2_2
X_15923_ _07933_ _07935_ _07934_ VGND VGND VPWR VPWR _08018_ sky130_fd_sc_hd__o21a_1
X_18711_ _10255_ _10687_ _10615_ _10620_ VGND VGND VPWR VPWR _10688_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19691_ _11573_ _11415_ _11574_ _11575_ _11576_ VGND VGND VPWR VPWR _11577_ sky130_fd_sc_hd__a221o_1
XFILLER_0_200_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18642_ _10618_ _10619_ VGND VGND VPWR VPWR _10620_ sky130_fd_sc_hd__xnor2_1
X_15854_ net461 net519 VGND VGND VPWR VPWR _07950_ sky130_fd_sc_hd__nand2_1
X_14805_ _06935_ _07004_ _06989_ VGND VGND VPWR VPWR _07005_ sky130_fd_sc_hd__o21a_1
XFILLER_0_189_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18573_ _10472_ _10474_ _10551_ VGND VGND VPWR VPWR _10552_ sky130_fd_sc_hd__a21oi_2
X_15785_ _07867_ _07881_ VGND VGND VPWR VPWR _07882_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17524_ _09418_ _09421_ _09510_ VGND VGND VPWR VPWR _09511_ sky130_fd_sc_hd__or3_1
X_14736_ _06900_ _06938_ VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17455_ _09379_ _09384_ _09375_ VGND VGND VPWR VPWR _09442_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14667_ _06831_ _06846_ VGND VGND VPWR VPWR _06871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16406_ _08416_ _08418_ _08494_ VGND VGND VPWR VPWR _08495_ sky130_fd_sc_hd__a21oi_2
X_13618_ _05815_ _05821_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__xor2_1
XFILLER_0_145_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17386_ _09369_ _09372_ VGND VGND VPWR VPWR _09373_ sky130_fd_sc_hd__xnor2_2
X_14598_ _06697_ _06740_ VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__xor2_1
XFILLER_0_116_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19125_ _05430_ _11094_ VGND VGND VPWR VPWR _11095_ sky130_fd_sc_hd__nor2_4
X_16337_ _08415_ _08426_ VGND VGND VPWR VPWR _08427_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13549_ net32 _05682_ _05687_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19056_ _10993_ _11027_ VGND VGND VPWR VPWR _11029_ sky130_fd_sc_hd__and2_1
X_16268_ _08357_ _08358_ VGND VGND VPWR VPWR _08359_ sky130_fd_sc_hd__xor2_1
XFILLER_0_112_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18007_ _09935_ _09936_ _09991_ VGND VGND VPWR VPWR _09992_ sky130_fd_sc_hd__a21bo_1
X_15219_ _07309_ _07312_ _07317_ VGND VGND VPWR VPWR _07318_ sky130_fd_sc_hd__o21a_1
XFILLER_0_164_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16199_ _08287_ net500 net476 VGND VGND VPWR VPWR _08291_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19958_ _11654_ _11510_ _11633_ _11827_ VGND VGND VPWR VPWR _11828_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_87_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_87_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_184_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18909_ _10881_ _10883_ net320 VGND VGND VPWR VPWR _10884_ sky130_fd_sc_hd__o21ai_1
X_19889_ _11761_ _11763_ VGND VGND VPWR VPWR _11764_ sky130_fd_sc_hd__xor2_2
X_21920_ net165 _01459_ _01481_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21851_ _01410_ _01411_ _01412_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20802_ net254 _12559_ VGND VGND VPWR VPWR _12651_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24570_ _03921_ _03922_ _03924_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__a21oi_1
X_21782_ net1031 _01342_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__nor2_1
XFILLER_0_188_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23521_ _05460_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__clkbuf_4
X_20733_ _12570_ _12581_ VGND VGND VPWR VPWR _12582_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26240_ spi0.data_packed\[18\] spi0.data_packed\[19\] net697 VGND VGND VPWR VPWR
+ _05352_ sky130_fd_sc_hd__mux2_1
X_20664_ _12503_ _12512_ VGND VGND VPWR VPWR _12513_ sky130_fd_sc_hd__nand2_1
X_23452_ net88 _02878_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22403_ top0.cordic0.vec\[1\]\[10\] _01259_ _01958_ _01959_ _01960_ VGND VGND VPWR
+ VPWR _01961_ sky130_fd_sc_hd__a41o_1
X_23383_ net187 _02822_ _02823_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26171_ _05309_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__clkbuf_1
X_20595_ net281 _12443_ VGND VGND VPWR VPWR _12444_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25122_ top0.matmul0.matmul_stage_inst.mult2\[9\] _04470_ _03642_ VGND VGND VPWR
+ VPWR _04471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22334_ _01867_ _01868_ _01892_ _01745_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_171_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_3__f_clk_sys clknet_0_clk_sys VGND VGND VPWR VPWR clknet_3_3__leaf_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25053_ _04402_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22265_ _01824_ _01822_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24004_ _03353_ _03358_ _03361_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__a21o_1
X_21216_ _12646_ _12577_ VGND VGND VPWR VPWR _13060_ sky130_fd_sc_hd__or2_1
X_22196_ net109 net119 VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__or2b_1
XFILLER_0_130_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21147_ _12990_ _12991_ VGND VGND VPWR VPWR _12992_ sky130_fd_sc_hd__xnor2_1
Xfanout530 top0.pid_q.mult0.a\[4\] VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__clkbuf_2
Xfanout541 net542 VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__clkbuf_4
Xfanout552 top0.pid_q.state\[2\] VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__clkbuf_2
Xfanout563 top0.matmul0.matmul_stage_inst.state\[5\] VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__clkbuf_4
X_25955_ _05166_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__clkbuf_1
X_21078_ _11726_ net226 VGND VGND VPWR VPWR _12924_ sky130_fd_sc_hd__nor2_1
Xfanout574 top0.matmul0.matmul_stage_inst.state\[1\] VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__clkbuf_4
Xfanout585 net586 VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__buf_2
X_24906_ _03976_ _04254_ _04255_ _03827_ _04256_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__o221a_4
Xfanout596 net597 VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__buf_2
X_20029_ _11657_ _11893_ _11796_ _11518_ VGND VGND VPWR VPWR _11894_ sky130_fd_sc_hd__o211ai_1
X_25886_ _05103_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_197_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24837_ _03343_ _03200_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15570_ net480 _07668_ VGND VGND VPWR VPWR _07669_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24768_ _04118_ _04119_ _04105_ _04106_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_96_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14521_ _06629_ _06632_ _06634_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__a21bo_1
X_26507_ clknet_leaf_77_clk_sys _00130_ net631 VGND VGND VPWR VPWR top0.pid_d.prev_int\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23719_ _03067_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24699_ _03928_ _04051_ _04052_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17240_ top0.pid_q.curr_int\[14\] top0.pid_q.prev_int\[14\] VGND VGND VPWR VPWR _09244_
+ sky130_fd_sc_hd__nand2_1
X_14452_ _06652_ _06659_ VGND VGND VPWR VPWR _06660_ sky130_fd_sc_hd__xor2_2
X_26438_ clknet_leaf_79_clk_sys _00079_ net634 VGND VGND VPWR VPWR top0.kid\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13403_ top0.matmul0.alpha_pass\[12\] _05435_ _05474_ VGND VGND VPWR VPWR _05616_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_148_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17171_ _08235_ _09176_ _09183_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__o21ai_1
X_14383_ _06590_ _06591_ VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__xor2_4
XFILLER_0_181_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26369_ _05416_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16122_ _08184_ _08213_ VGND VGND VPWR VPWR _08215_ sky130_fd_sc_hd__nand2_1
X_13334_ _05540_ _05546_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16053_ _08146_ VGND VGND VPWR VPWR _08147_ sky130_fd_sc_hd__inv_2
X_13265_ top0.matmul0.alpha_pass\[3\] _05466_ _05474_ VGND VGND VPWR VPWR _05478_
+ sky130_fd_sc_hd__nand3_2
XFILLER_0_150_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15004_ _07127_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__clkbuf_1
X_13196_ net744 _05422_ state\[0\] _05426_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__a22o_1
X_19812_ _11448_ _11691_ _11675_ VGND VGND VPWR VPWR _11692_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19743_ _11621_ _11624_ _11626_ _11526_ VGND VGND VPWR VPWR _11627_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16955_ top0.currT_r\[9\] _08997_ _09011_ VGND VGND VPWR VPWR _09012_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_159_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15906_ _07919_ _07925_ _07924_ VGND VGND VPWR VPWR _08001_ sky130_fd_sc_hd__o21a_1
X_16886_ _05439_ _08947_ VGND VGND VPWR VPWR _08948_ sky130_fd_sc_hd__nand2_1
X_19674_ net150 net144 net138 net133 net199 net193 VGND VGND VPWR VPWR _11561_ sky130_fd_sc_hd__mux4_1
XFILLER_0_189_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18625_ _10440_ _10579_ VGND VGND VPWR VPWR _10603_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15837_ net538 net443 VGND VGND VPWR VPWR _07933_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_59_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18556_ _10533_ _10534_ VGND VGND VPWR VPWR _10535_ sky130_fd_sc_hd__or2b_2
X_15768_ _07861_ _07863_ VGND VGND VPWR VPWR _07865_ sky130_fd_sc_hd__and2_1
X_14719_ net31 _05666_ VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__nand2_1
X_17507_ _09493_ net385 VGND VGND VPWR VPWR _09494_ sky130_fd_sc_hd__nor2_1
X_18487_ net323 net379 VGND VGND VPWR VPWR _10467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15699_ top0.pid_q.out\[1\] top0.pid_q.curr_int\[1\] VGND VGND VPWR VPWR _07797_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_131_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17438_ _09421_ _09424_ VGND VGND VPWR VPWR _09425_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_15 _12739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_26 net1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_184_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_37 _11094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 net687 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17369_ _09355_ VGND VGND VPWR VPWR _09356_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19108_ _11029_ _11077_ _10992_ VGND VGND VPWR VPWR _11080_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_103_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20380_ _12227_ _12218_ _12219_ VGND VGND VPWR VPWR _12229_ sky130_fd_sc_hd__nand3_1
XFILLER_0_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19039_ _11003_ _11011_ VGND VGND VPWR VPWR _11012_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_24_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22050_ _01590_ _01611_ _01605_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21001_ _12846_ _12847_ VGND VGND VPWR VPWR _12848_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25740_ _04989_ net73 top0.matmul0.sin\[13\] VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__mux2_1
X_22952_ _02463_ _02464_ _02332_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__mux2_1
Xmax_cap17 _05430_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
X_21903_ _01462_ _01463_ _01464_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__a21o_1
X_25671_ _04883_ top0.matmul0.sin\[9\] _04941_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__nand3_1
X_22883_ _02374_ top0.svm0.tB\[12\] VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__and2_1
XFILLER_0_179_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24622_ _03742_ _03827_ _03741_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__a21oi_2
X_21834_ _01333_ _01395_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_167_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24553_ _03741_ _03827_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__nor2_2
X_21765_ net133 net1031 VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_66_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23504_ _02917_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__clkbuf_1
X_20716_ _11673_ _12561_ _12563_ VGND VGND VPWR VPWR _12565_ sky130_fd_sc_hd__and3_1
X_27272_ clknet_3_7__leaf_clk_mosi _00886_ VGND VGND VPWR VPWR spi0.data_packed\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24484_ _03816_ _03839_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__xnor2_2
X_21696_ _01197_ _01257_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__or2_1
XFILLER_0_163_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26223_ _05343_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__clkbuf_1
X_23435_ _02868_ _02871_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__xor2_1
X_20647_ _12495_ net263 _12490_ VGND VGND VPWR VPWR _12496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_191_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26154_ spi0.data_packed\[3\] _05292_ net18 VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20578_ _12342_ _12426_ VGND VGND VPWR VPWR _12427_ sky130_fd_sc_hd__xnor2_2
X_23366_ _02796_ _02797_ _11513_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__o21ai_1
X_25105_ _04452_ _04453_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__and2b_1
X_22317_ net210 VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26085_ top0.matmul0.alpha_pass\[13\] _05237_ _05265_ VGND VGND VPWR VPWR _05266_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23297_ _02741_ _02743_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__xnor2_2
X_25036_ _04382_ _04384_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__nand2_1
X_22248_ _01684_ _01737_ _01738_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_44_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22179_ net745 _12813_ _01740_ _12963_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__a22o_1
X_26987_ clknet_leaf_27_clk_sys _00604_ net615 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[3\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout360 net361 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkbuf_4
Xfanout371 net372 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__buf_2
XFILLER_0_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16740_ _08287_ net445 _08823_ VGND VGND VPWR VPWR _08824_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout382 net384 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_4
X_13952_ _06121_ _06122_ _06119_ _06120_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__a211o_1
X_25938_ top0.matmul0.alpha_pass\[14\] net428 VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__nor2_1
Xfanout393 net394 VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkbuf_4
X_16671_ _08453_ _08720_ net498 _08447_ VGND VGND VPWR VPWR _08756_ sky130_fd_sc_hd__o211a_1
X_13883_ _05573_ _05538_ _05539_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__nor3_1
X_25869_ top0.matmul0.alpha_pass\[9\] top0.matmul0.beta_pass\[9\] VGND VGND VPWR VPWR
+ _05088_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_201_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18410_ _10381_ _10390_ VGND VGND VPWR VPWR _10391_ sky130_fd_sc_hd__and2_1
X_15622_ net474 net514 VGND VGND VPWR VPWR _07720_ sky130_fd_sc_hd__nand2_1
XFILLER_0_198_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19390_ net431 _09892_ _09893_ _11295_ VGND VGND VPWR VPWR _11296_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18341_ _10319_ _10321_ VGND VGND VPWR VPWR _10323_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_186_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15553_ net451 net538 VGND VGND VPWR VPWR _07652_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14504_ _06707_ _06710_ VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__xnor2_2
X_18272_ net406 _09353_ _10074_ _10253_ VGND VGND VPWR VPWR _10254_ sky130_fd_sc_hd__a31o_1
X_15484_ _07286_ _07291_ _07582_ VGND VGND VPWR VPWR _07583_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17223_ _09222_ _09192_ _09228_ _09135_ _09229_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__a221o_1
X_14435_ net28 _06640_ VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__nand2_1
XFILLER_0_181_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17154_ net553 _09167_ _09168_ net548 _08942_ VGND VGND VPWR VPWR _09169_ sky130_fd_sc_hd__a32o_1
X_14366_ _06494_ _06499_ _06492_ VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16105_ _08189_ _08197_ VGND VGND VPWR VPWR _08198_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13317_ net48 VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17085_ top0.pid_q.curr_error\[1\] _00011_ _09117_ VGND VGND VPWR VPWR _09119_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_172_Right_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14297_ _06425_ _06505_ VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16036_ _08049_ _08129_ VGND VGND VPWR VPWR _08130_ sky130_fd_sc_hd__xnor2_1
X_13248_ _05461_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17987_ _09885_ _09883_ _09888_ VGND VGND VPWR VPWR _09973_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19726_ net277 _11602_ VGND VGND VPWR VPWR _11610_ sky130_fd_sc_hd__and2_1
XFILLER_0_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16938_ top0.currT_r\[8\] _08984_ _08985_ VGND VGND VPWR VPWR _08996_ sky130_fd_sc_hd__o21a_1
X_19657_ _11543_ _11531_ _11533_ _11534_ VGND VGND VPWR VPWR _11545_ sky130_fd_sc_hd__nand4_1
X_16869_ top0.currT_r\[3\] _08917_ _08931_ VGND VGND VPWR VPWR _08932_ sky130_fd_sc_hd__o21a_1
XFILLER_0_189_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18608_ _10585_ _10505_ _10582_ _10438_ VGND VGND VPWR VPWR _10587_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_88_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19588_ _11474_ _11475_ _11476_ VGND VGND VPWR VPWR _11477_ sky130_fd_sc_hd__or3b_1
XFILLER_0_75_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18539_ net385 _09518_ _09494_ _10074_ VGND VGND VPWR VPWR _10518_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21550_ net115 net109 VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__and2b_2
XFILLER_0_63_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20501_ net302 _12349_ VGND VGND VPWR VPWR _12350_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21481_ net242 _01006_ net218 VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_173_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20432_ _12279_ _12280_ VGND VGND VPWR VPWR _12281_ sky130_fd_sc_hd__xnor2_1
X_23220_ net165 _11519_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__nor2_1
XFILLER_0_200_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23151_ top0.svm0.delta\[15\] _02636_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__or2_1
X_20363_ net271 net277 VGND VGND VPWR VPWR _12212_ sky130_fd_sc_hd__or2b_1
XFILLER_0_101_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22102_ _01660_ _01640_ _01645_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__mux2_1
X_23082_ top0.periodTop_r\[4\] top0.svm0.counter\[4\] VGND VGND VPWR VPWR _02583_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20294_ net261 net269 VGND VGND VPWR VPWR _12143_ sky130_fd_sc_hd__or2b_1
XFILLER_0_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26910_ clknet_leaf_110_clk_sys _00527_ net579 VGND VGND VPWR VPWR top0.matmul0.sin\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_22033_ _01355_ _01275_ _01594_ net162 VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26841_ clknet_leaf_45_clk_sys _00458_ net681 VGND VGND VPWR VPWR top0.svm0.delta\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_26772_ clknet_leaf_7_clk_sys _00389_ net593 VGND VGND VPWR VPWR top0.cordic0.cos\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_23984_ _03336_ _03340_ _03341_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__a21o_2
XFILLER_0_199_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25723_ top0.matmul0.sin\[8\] _04979_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__xnor2_1
X_22935_ _02440_ _02448_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25654_ net71 _04928_ _04929_ net73 _04878_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__a221o_1
X_22866_ top0.svm0.tB\[3\] _02384_ _02339_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24605_ _03863_ _03959_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__xnor2_1
X_21817_ _01328_ _01378_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__xnor2_2
X_25585_ _04880_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22797_ top0.svm0.counter\[13\] VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24536_ _03801_ _03802_ VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__or2_1
X_21748_ net136 VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27255_ clknet_3_2__leaf_clk_mosi _00869_ VGND VGND VPWR VPWR spi0.data_packed\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_24467_ _03572_ _03687_ _03689_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__and3_1
X_21679_ _01232_ _01235_ _01240_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14220_ _06427_ _06428_ _06429_ _06430_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26206_ spi0.data_packed\[1\] spi0.data_packed\[2\] net695 VGND VGND VPWR VPWR _05335_
+ sky130_fd_sc_hd__mux2_1
X_23418_ _02846_ _02848_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__or2_1
X_27186_ clknet_leaf_57_clk_sys _00800_ net645 VGND VGND VPWR VPWR top0.currT_r\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_184_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24398_ _03663_ _03754_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14151_ _06119_ _06120_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__nor2_1
X_26137_ net18 spi0.data_packed\[15\] VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23349_ _11526_ _02792_ net176 VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14082_ _06288_ _06293_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_131_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26068_ top0.pid_d.out\[9\] _05232_ _05233_ spi0.data_packed\[73\] VGND VGND VPWR
+ VPWR _05253_ sky130_fd_sc_hd__a22o_1
X_25019_ _04279_ _04281_ _04280_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__a21o_1
X_17910_ _09896_ _09895_ top0.pid_d.out\[0\] VGND VGND VPWR VPWR _09897_ sky130_fd_sc_hd__mux2_1
X_18890_ net371 net314 VGND VGND VPWR VPWR _10865_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17841_ net326 net414 VGND VGND VPWR VPWR _09828_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14984_ _06276_ _07114_ _07115_ VGND VGND VPWR VPWR _07116_ sky130_fd_sc_hd__mux2_1
X_17772_ net379 net355 VGND VGND VPWR VPWR _09759_ sky130_fd_sc_hd__nand2_1
Xfanout190 top0.cordic0.gm0.iter\[2\] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
X_19511_ _11399_ _11400_ _11401_ VGND VGND VPWR VPWR _11402_ sky130_fd_sc_hd__a21o_1
X_13935_ net56 _05723_ _05724_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__and3_1
X_16723_ _08769_ _08774_ _08771_ VGND VGND VPWR VPWR _08807_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19442_ net431 _11292_ VGND VGND VPWR VPWR _11340_ sky130_fd_sc_hd__and2_1
X_16654_ _08619_ _08626_ _08618_ VGND VGND VPWR VPWR _08740_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_159_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13866_ _05922_ _05949_ _06075_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__or3_1
XFILLER_0_88_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15605_ _07703_ VGND VGND VPWR VPWR _07704_ sky130_fd_sc_hd__buf_2
X_16585_ _08670_ _08671_ VGND VGND VPWR VPWR _08672_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19373_ net879 _11285_ _11288_ top0.pid_d.curr_error\[6\] VGND VGND VPWR VPWR _00316_
+ sky130_fd_sc_hd__a22o_1
X_13797_ _06005_ _06006_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__and2_1
XFILLER_0_186_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18324_ _10202_ _10220_ _10305_ VGND VGND VPWR VPWR _10306_ sky130_fd_sc_hd__a21oi_2
X_15536_ _07632_ _07634_ VGND VGND VPWR VPWR _07635_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18255_ _10131_ _10147_ _10237_ VGND VGND VPWR VPWR _10238_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_84_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15467_ net528 net462 VGND VGND VPWR VPWR _07566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17206_ _08550_ _09192_ _09214_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14418_ _06624_ _06625_ VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18186_ net331 net382 VGND VGND VPWR VPWR _10169_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15398_ net541 top0.pid_q.mult0.a\[1\] net472 VGND VGND VPWR VPWR _07497_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17137_ top0.pid_q.prev_int\[2\] VGND VGND VPWR VPWR _09153_ sky130_fd_sc_hd__inv_2
X_14349_ _06513_ _06528_ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17068_ _09108_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16019_ _08109_ _08112_ VGND VGND VPWR VPWR _08113_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19709_ net182 net188 _11427_ net179 VGND VGND VPWR VPWR _11594_ sky130_fd_sc_hd__a31o_1
X_20981_ net225 net222 _12817_ VGND VGND VPWR VPWR _12828_ sky130_fd_sc_hd__and3_1
XFILLER_0_170_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_69_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22720_ net733 _12004_ _12740_ _02270_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__a31o_1
XFILLER_0_192_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22651_ _02144_ _02143_ _02163_ _02203_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__a31o_1
XFILLER_0_165_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21602_ net110 net96 _01163_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__a21oi_1
X_25370_ _04521_ _04697_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__xor2_1
XFILLER_0_63_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22582_ _02080_ _02123_ _02122_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24321_ _03677_ _03166_ _03154_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_8_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21533_ _01088_ _01092_ _01094_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_161_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27040_ clknet_leaf_7_clk_sys _00657_ net593 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_24252_ _03482_ _03520_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21464_ net231 _12770_ _12814_ _12769_ _11759_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_78_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23203_ _02653_ _02654_ _11409_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__mux2_1
X_20415_ net295 net298 VGND VGND VPWR VPWR _12264_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_16_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24183_ _03185_ _03114_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__nor2_1
X_21395_ _00954_ _00956_ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23134_ net959 _02623_ _02624_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20346_ _12176_ _12178_ _12194_ VGND VGND VPWR VPWR _12195_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23065_ _05565_ top0.svm0.counter\[8\] VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__nand2_1
X_20277_ net267 top0.cordic0.vec\[0\]\[8\] VGND VGND VPWR VPWR _12126_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_102_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22016_ net136 _01512_ _01319_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26824_ clknet_leaf_37_clk_sys net707 net679 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_87_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26755_ clknet_leaf_5_clk_sys _00372_ net590 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_23967_ _03250_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__buf_4
XFILLER_0_168_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13720_ net50 _05484_ _05486_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__and3_1
X_25706_ net871 _04964_ _04936_ _04968_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__a22o_1
X_22918_ _02298_ _02434_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26686_ clknet_leaf_83_clk_sys _00303_ net647 VGND VGND VPWR VPWR top0.pid_d.curr_error\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_23898_ _03249_ _03253_ _03255_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13651_ _05811_ _05812_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__xor2_1
X_25637_ _04914_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__inv_2
X_22849_ top0.svm0.tA\[8\] _02366_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16370_ _08339_ _08346_ _08337_ VGND VGND VPWR VPWR _08460_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13582_ _05710_ _05712_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__and2_1
XFILLER_0_155_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25568_ _04871_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15321_ _07373_ _07419_ VGND VGND VPWR VPWR _07420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24519_ _03057_ _03058_ _03196_ _03197_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25499_ _04835_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18040_ net346 net375 VGND VGND VPWR VPWR _10025_ sky130_fd_sc_hd__nand2_2
XFILLER_0_109_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27238_ clknet_3_7__leaf_clk_mosi _00852_ VGND VGND VPWR VPWR spi0.data_packed\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_15252_ _07332_ _07349_ VGND VGND VPWR VPWR _07351_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14203_ _06288_ _06293_ _06285_ VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27169_ clknet_leaf_32_clk_sys _00783_ net664 VGND VGND VPWR VPWR top0.periodTop_r\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_15183_ net535 net460 VGND VGND VPWR VPWR _07282_ sky130_fd_sc_hd__nand2_2
XFILLER_0_201_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14134_ _06181_ _06203_ _06345_ VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19991_ _11431_ _11856_ net177 VGND VGND VPWR VPWR _11859_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14065_ top0.svm0.state\[1\] top0.svm0.state\[0\] net171 VGND VGND VPWR VPWR _06278_
+ sky130_fd_sc_hd__a21o_1
X_18942_ net435 _10828_ _10829_ VGND VGND VPWR VPWR _10917_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18873_ _10772_ VGND VGND VPWR VPWR _10848_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17824_ _09647_ _09684_ VGND VGND VPWR VPWR _09811_ sky130_fd_sc_hd__or2b_1
XFILLER_0_146_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2 spi0.cs_sync\[1\] VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__dlygate4sd3_1
X_14967_ _07105_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__clkbuf_1
X_17755_ _09513_ _09456_ _09741_ VGND VGND VPWR VPWR _09742_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_159_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16706_ _08745_ _08790_ VGND VGND VPWR VPWR _08791_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_199_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13918_ _05721_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__buf_4
X_17686_ _09671_ _09672_ VGND VGND VPWR VPWR _09673_ sky130_fd_sc_hd__xnor2_1
X_14898_ _07069_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19425_ top0.pid_d.curr_int\[5\] top0.pid_d.prev_int\[5\] VGND VGND VPWR VPWR _11326_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16637_ _08717_ _08722_ VGND VGND VPWR VPWR _08723_ sky130_fd_sc_hd__xnor2_1
X_13849_ net62 _06047_ _06045_ _06023_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19356_ top0.pid_d.curr_error\[12\] _11243_ _11276_ VGND VGND VPWR VPWR _11282_ sky130_fd_sc_hd__mux2_1
X_16568_ net501 _08654_ net459 VGND VGND VPWR VPWR _08655_ sky130_fd_sc_hd__or3b_1
XFILLER_0_71_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18307_ net344 net348 VGND VGND VPWR VPWR _10289_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15519_ net492 net506 VGND VGND VPWR VPWR _07618_ sky130_fd_sc_hd__nand2_1
X_16499_ _08579_ _08586_ VGND VGND VPWR VPWR _08587_ sky130_fd_sc_hd__xnor2_2
X_19287_ _11227_ _11228_ VGND VGND VPWR VPWR _11230_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18238_ _10202_ _10220_ VGND VGND VPWR VPWR _10221_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18169_ _10151_ _10152_ VGND VGND VPWR VPWR _10153_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20200_ net283 net276 VGND VGND VPWR VPWR _12049_ sky130_fd_sc_hd__and2b_2
X_21180_ _11689_ _12982_ VGND VGND VPWR VPWR _13024_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20131_ top0.cordic0.slte0.opA\[14\] _11775_ _11967_ VGND VGND VPWR VPWR _11987_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20062_ top0.cordic0.slte0.opA\[9\] _11918_ VGND VGND VPWR VPWR _11924_ sky130_fd_sc_hd__and2_1
X_24870_ _04218_ _04221_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_174_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23821_ _02994_ _02996_ _02989_ _02991_ VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__o22a_1
XFILLER_0_139_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26540_ clknet_leaf_60_clk_sys _00163_ net653 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[14\]
+ sky130_fd_sc_hd__dfrtp_2
X_23752_ _03102_ _03109_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__xnor2_4
X_20964_ _12003_ _12035_ VGND VGND VPWR VPWR _12812_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22703_ _02250_ _02253_ _01948_ _01248_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__o2bb2a_1
X_26471_ clknet_leaf_12_clk_sys _00102_ net603 VGND VGND VPWR VPWR top0.periodTop\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_23683_ _03010_ _03040_ _03038_ _03039_ VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20895_ top0.cordic0.domain\[0\] net211 VGND VGND VPWR VPWR _12743_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25422_ _04759_ _04761_ _04765_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22634_ _01213_ _01063_ net78 VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__a21o_1
XFILLER_0_193_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25353_ _04516_ _04642_ _04571_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__a21o_1
XFILLER_0_192_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22565_ _01948_ _02025_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24304_ _03229_ _03230_ _03291_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__a21bo_1
X_21516_ net143 net139 VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__nor2b_4
X_25284_ _04541_ _04542_ _04629_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22496_ _02017_ _02022_ _02028_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27023_ clknet_leaf_15_clk_sys _00640_ net614 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_24235_ _03591_ _03592_ _03588_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21447_ _01011_ _01012_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24166_ _03511_ _03516_ _03520_ _03522_ _03523_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_43_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21378_ _00944_ _00945_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__xor2_1
X_23117_ top0.svm0.delta\[6\] _02609_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__or2_1
X_20329_ _12175_ _12150_ _12151_ _12177_ VGND VGND VPWR VPWR _12178_ sky130_fd_sc_hd__nand4_2
X_24097_ _03454_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23048_ top0.svm0.counter\[15\] _06777_ _02543_ top0.svm0.counter\[14\] VGND VGND
+ VPWR VPWR _02549_ sky130_fd_sc_hd__or4b_1
X_15870_ _07828_ _07830_ _07826_ VGND VGND VPWR VPWR _07966_ sky130_fd_sc_hd__o21a_1
X_14821_ _07019_ _07020_ VGND VGND VPWR VPWR _07021_ sky130_fd_sc_hd__nand2_1
X_26807_ clknet_leaf_69_clk_sys _00424_ net662 VGND VGND VPWR VPWR top0.pid_q.prev_int\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_24999_ _02982_ _04272_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14752_ net23 _05723_ _05724_ VGND VGND VPWR VPWR _06954_ sky130_fd_sc_hd__and3_1
X_17540_ _09522_ _09523_ _09526_ VGND VGND VPWR VPWR _09527_ sky130_fd_sc_hd__a21o_1
X_26738_ clknet_leaf_101_clk_sys _00355_ net587 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[13\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_98_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13703_ _05607_ _05543_ _05545_ net61 _05585_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__o311a_1
XFILLER_0_6_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17471_ _09375_ _09379_ _09457_ VGND VGND VPWR VPWR _09458_ sky130_fd_sc_hd__o21ai_1
X_14683_ net31 _06881_ _06883_ _05731_ _06886_ VGND VGND VPWR VPWR _06887_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26669_ clknet_leaf_82_clk_sys _00286_ net646 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19210_ top0.matmul0.alpha_pass\[4\] _11150_ VGND VGND VPWR VPWR _11160_ sky130_fd_sc_hd__nor2_1
X_13634_ _05832_ _05844_ _05846_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__o21a_1
X_16422_ net461 net466 VGND VGND VPWR VPWR _08511_ sky130_fd_sc_hd__xor2_1
XFILLER_0_157_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16353_ _08364_ _08375_ _08362_ VGND VGND VPWR VPWR _08443_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_6_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19141_ top0.kid\[5\] _11098_ _11100_ top0.kpd\[5\] VGND VGND VPWR VPWR _11106_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13565_ net49 net46 _05585_ _05587_ _05697_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__a41o_1
XFILLER_0_27_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15304_ net487 _07401_ _07402_ VGND VGND VPWR VPWR _07403_ sky130_fd_sc_hd__a21o_1
X_19072_ _11042_ _11014_ _11016_ _11040_ VGND VGND VPWR VPWR _11044_ sky130_fd_sc_hd__o2bb2a_1
X_16284_ _08369_ _08374_ VGND VGND VPWR VPWR _08375_ sky130_fd_sc_hd__xnor2_2
X_13496_ _05695_ _05708_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18023_ _09918_ _09929_ _09916_ VGND VGND VPWR VPWR _10008_ sky130_fd_sc_hd__a21o_1
X_15235_ _07304_ _07319_ VGND VGND VPWR VPWR _07334_ sky130_fd_sc_hd__nor2_1
X_15166_ _07203_ _07208_ VGND VGND VPWR VPWR _07265_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14117_ _05500_ _05468_ _05471_ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__nor3_2
XFILLER_0_201_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15097_ _07191_ _07195_ VGND VGND VPWR VPWR _07196_ sky130_fd_sc_hd__xnor2_1
X_19974_ top0.cordic0.slte0.opA\[3\] _11841_ _11842_ _11840_ VGND VGND VPWR VPWR _00363_
+ sky130_fd_sc_hd__a22o_1
X_14048_ _06161_ _06164_ _06165_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__and3_1
X_18925_ _10892_ _10899_ VGND VGND VPWR VPWR _10900_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18856_ net435 _09339_ _10831_ VGND VGND VPWR VPWR _10832_ sky130_fd_sc_hd__and3_1
XFILLER_0_197_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17807_ _09792_ _09793_ VGND VGND VPWR VPWR _09794_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18787_ _10763_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__clkbuf_1
X_15999_ net532 top0.pid_q.mult0.b\[15\] VGND VGND VPWR VPWR _08093_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_55_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17738_ _09699_ _09704_ VGND VGND VPWR VPWR _09725_ sky130_fd_sc_hd__xor2_1
XFILLER_0_194_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17669_ net404 net337 VGND VGND VPWR VPWR _09656_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19408_ _11308_ _11310_ VGND VGND VPWR VPWR _11311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20680_ net263 _12525_ VGND VGND VPWR VPWR _12529_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19339_ net438 _11123_ VGND VGND VPWR VPWR _11276_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_83_clk_sys clknet_3_4__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_83_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22350_ _01845_ _01901_ _01906_ net97 _01908_ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21301_ _13143_ VGND VGND VPWR VPWR _13144_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22281_ _01311_ _01075_ _01840_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24020_ _03335_ _03377_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21232_ _12583_ _13075_ VGND VGND VPWR VPWR _13076_ sky130_fd_sc_hd__xnor2_1
Xhold210 top0.pid_d.curr_error\[13\] VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 top0.c_out_calc\[15\] VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold232 top0.cordic0.slte0.opA\[8\] VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 top0.matmul0.b\[15\] VGND VGND VPWR VPWR net943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold254 _05372_ VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 top0.b_in_matmul\[5\] VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__dlygate4sd3_1
X_21163_ _12965_ _13007_ VGND VGND VPWR VPWR _13008_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_141_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold276 top0.pid_q.prev_int\[7\] VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 top0.matmul0.a\[3\] VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout701 net513 VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__buf_4
Xhold298 top0.b_in_matmul\[1\] VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__dlygate4sd3_1
X_20114_ net1014 _11971_ net177 VGND VGND VPWR VPWR _11972_ sky130_fd_sc_hd__o21ai_1
X_25971_ _05178_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__clkbuf_1
X_21094_ _12938_ _12939_ VGND VGND VPWR VPWR _12940_ sky130_fd_sc_hd__or2b_1
X_24922_ _03474_ _04272_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__nor2_1
X_20045_ _11880_ _11908_ VGND VGND VPWR VPWR _11909_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24853_ _03313_ _03889_ _04099_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23804_ net572 top0.matmul0.matmul_stage_inst.d\[13\] top0.matmul0.matmul_stage_inst.c\[13\]
+ net556 VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__a22o_2
XFILLER_0_198_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24784_ _03990_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__inv_2
X_21996_ _01175_ _01455_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_197_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26523_ clknet_leaf_61_clk_sys _00146_ net651 VGND VGND VPWR VPWR top0.pid_q.out\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_178_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23735_ net570 net575 top0.matmul0.matmul_stage_inst.f\[10\] VGND VGND VPWR VPWR
+ _03093_ sky130_fd_sc_hd__o21a_2
XFILLER_0_96_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20947_ _12783_ _12708_ VGND VGND VPWR VPWR _12795_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26454_ clknet_leaf_55_clk_sys _00095_ net668 VGND VGND VPWR VPWR top0.kiq\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_23666_ net574 top0.matmul0.matmul_stage_inst.d\[9\] top0.matmul0.matmul_stage_inst.c\[9\]
+ net558 VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__a22o_4
XFILLER_0_37_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20878_ _12722_ _12723_ _12726_ VGND VGND VPWR VPWR _12727_ sky130_fd_sc_hd__and3_1
X_25405_ _04411_ _04694_ _04646_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22617_ _02168_ _02170_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__nor2_2
X_26385_ clknet_leaf_41_clk_sys _00026_ net685 VGND VGND VPWR VPWR top0.svm0.tC\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23597_ _02965_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25336_ _04675_ _04679_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__or2_1
X_13350_ _05561_ _05562_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__xor2_1
XFILLER_0_180_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22548_ net119 net104 _01069_ _02102_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_134_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25267_ _03200_ _04518_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__nor2_2
XFILLER_0_162_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13281_ top0.matmul0.beta_pass\[2\] _05466_ _05470_ _05463_ top0.c_out_calc\[2\]
+ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__a32o_1
X_22479_ _02011_ _02035_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__xnor2_2
X_27006_ clknet_leaf_25_clk_sys _00623_ net627 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_15020_ _07135_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24218_ _03572_ _03323_ _03561_ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25198_ _04477_ _04478_ _04476_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24149_ _03491_ _03492_ VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__xnor2_1
X_16971_ _09025_ _09019_ _09026_ VGND VGND VPWR VPWR _09027_ sky130_fd_sc_hd__a21o_1
X_18710_ net377 _09518_ _10074_ _10612_ VGND VGND VPWR VPWR _10687_ sky130_fd_sc_hd__a22o_1
X_15922_ _08013_ _08016_ VGND VGND VPWR VPWR _08017_ sky130_fd_sc_hd__xnor2_1
X_19690_ _11420_ VGND VGND VPWR VPWR _11576_ sky130_fd_sc_hd__clkbuf_4
X_18641_ net390 net309 VGND VGND VPWR VPWR _10619_ sky130_fd_sc_hd__nand2_1
X_15853_ net458 net521 VGND VGND VPWR VPWR _07949_ sky130_fd_sc_hd__nand2_1
X_14804_ _06943_ _06949_ VGND VGND VPWR VPWR _07004_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18572_ _10472_ _10474_ _10473_ VGND VGND VPWR VPWR _10551_ sky130_fd_sc_hd__o21a_1
X_15784_ _07869_ _07880_ VGND VGND VPWR VPWR _07881_ sky130_fd_sc_hd__xor2_1
XFILLER_0_54_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17523_ _09413_ _09424_ VGND VGND VPWR VPWR _09510_ sky130_fd_sc_hd__nand2_1
X_14735_ _06913_ _06937_ VGND VGND VPWR VPWR _06938_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14666_ top0.periodTop_r\[9\] _06867_ _06868_ _06869_ VGND VGND VPWR VPWR _06870_
+ sky130_fd_sc_hd__a31o_1
X_17454_ _09440_ VGND VGND VPWR VPWR _09441_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13617_ _05596_ _05829_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__xnor2_4
X_16405_ _08416_ _08418_ _08417_ VGND VGND VPWR VPWR _08494_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14597_ _06800_ _06794_ _06801_ VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__a21oi_1
X_17385_ _09370_ _09371_ VGND VGND VPWR VPWR _09372_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19124_ top0.pid_d.state\[0\] net433 _07136_ VGND VGND VPWR VPWR _11094_ sky130_fd_sc_hd__nor3_4
X_16336_ _08420_ _08425_ VGND VGND VPWR VPWR _08426_ sky130_fd_sc_hd__xor2_1
X_13548_ net32 _05682_ _05687_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16267_ net456 net510 VGND VGND VPWR VPWR _08358_ sky130_fd_sc_hd__nand2_1
X_19055_ _10993_ _11027_ VGND VGND VPWR VPWR _11028_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13479_ _05685_ _05691_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18006_ _09935_ _09936_ _09937_ VGND VGND VPWR VPWR _09991_ sky130_fd_sc_hd__o21ai_1
X_15218_ _07313_ _07316_ VGND VGND VPWR VPWR _07317_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16198_ net473 net501 VGND VGND VPWR VPWR _08290_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15149_ _07245_ _07246_ _07247_ VGND VGND VPWR VPWR _07248_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19957_ net185 _11510_ _11657_ VGND VGND VPWR VPWR _11827_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18908_ _10712_ _10882_ _10710_ VGND VGND VPWR VPWR _10883_ sky130_fd_sc_hd__a21oi_1
X_19888_ _11515_ _11762_ VGND VGND VPWR VPWR _11763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18839_ _10813_ _10814_ VGND VGND VPWR VPWR _10815_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21850_ _01380_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20801_ _12552_ _12555_ VGND VGND VPWR VPWR _12650_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21781_ net130 net121 net1031 _01342_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__and4_1
XFILLER_0_72_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23520_ _02925_ VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__clkbuf_1
X_20732_ _12253_ _12572_ VGND VGND VPWR VPWR _12581_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_186_Right_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23451_ _02879_ _02878_ _02877_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__a21o_1
X_20663_ _12305_ _12510_ _12511_ VGND VGND VPWR VPWR _12512_ sky130_fd_sc_hd__or3b_2
XFILLER_0_163_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22402_ _01259_ _01954_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__and2b_1
XFILLER_0_34_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26170_ _05308_ top0.cordic0.slte0.opB\[9\] _12006_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__mux2_1
X_23382_ net215 _11448_ _11730_ _02713_ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__a22o_1
X_20594_ _12057_ _12284_ _12441_ net302 _12442_ VGND VGND VPWR VPWR _12443_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25121_ _04404_ _04469_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__xnor2_1
X_22333_ _01867_ _01869_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25052_ top0.matmul0.matmul_stage_inst.mult2\[8\] _04401_ _03642_ VGND VGND VPWR
+ VPWR _04402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22264_ _01066_ net96 VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__nand2_1
X_24003_ _03302_ _03360_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__xnor2_4
X_21215_ _12544_ _12545_ _13058_ VGND VGND VPWR VPWR _13059_ sky130_fd_sc_hd__or3_1
XFILLER_0_143_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22195_ net78 net89 VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__xor2_2
X_21146_ _12180_ _12824_ VGND VGND VPWR VPWR _12991_ sky130_fd_sc_hd__or2_1
Xfanout520 net521 VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__clkbuf_4
Xfanout531 net533 VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__buf_4
Xfanout542 top0.pid_q.mult0.a\[0\] VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__clkbuf_4
X_25954_ top0.matmul0.op_in\[0\] _05162_ _05165_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__mux2_1
X_21077_ _12697_ _12851_ _12922_ VGND VGND VPWR VPWR _12923_ sky130_fd_sc_hd__or3_1
Xfanout553 top0.pid_q.state\[1\] VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__clkbuf_4
Xfanout564 top0.matmul0.matmul_stage_inst.state\[4\] VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__buf_4
Xfanout575 top0.matmul0.matmul_stage_inst.state\[1\] VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__clkbuf_2
Xfanout586 net606 VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__clkbuf_2
X_24905_ _04252_ _04174_ _04253_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__a21o_1
Xfanout597 net598 VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__clkbuf_2
X_20028_ _11892_ _11824_ VGND VGND VPWR VPWR _11893_ sky130_fd_sc_hd__nor2_1
X_25885_ top0.matmul0.alpha_pass\[9\] top0.matmul0.beta_pass\[9\] VGND VGND VPWR VPWR
+ _05103_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24836_ _03474_ _04097_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24767_ _04105_ _04106_ _04118_ _04119_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_14_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21979_ _01493_ _01514_ _01519_ _01530_ _01540_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__a221o_1
X_14520_ _06714_ _06726_ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23718_ _03066_ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__clkbuf_4
X_26506_ clknet_leaf_78_clk_sys _00129_ net639 VGND VGND VPWR VPWR top0.pid_d.prev_int\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24698_ _03931_ _04050_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14451_ _06654_ _06658_ VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23649_ _02993_ _02995_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__nor2_2
X_26437_ clknet_leaf_79_clk_sys _00078_ net632 VGND VGND VPWR VPWR top0.kid\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13402_ _05606_ _05614_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_181_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17170_ top0.pid_q.curr_int\[6\] _09141_ _09182_ _09136_ VGND VGND VPWR VPWR _09183_
+ sky130_fd_sc_hd__a22oi_1
X_14382_ _06437_ net1015 net23 VGND VGND VPWR VPWR _06591_ sky130_fd_sc_hd__and3b_1
X_26368_ spi0.opcode\[2\] spi0.opcode\[3\] net691 VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16121_ _08184_ _08213_ VGND VGND VPWR VPWR _08214_ sky130_fd_sc_hd__nor2_1
X_25319_ _04382_ _04647_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__nand2_2
X_13333_ _05541_ _05543_ _05545_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__or3_1
XFILLER_0_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26299_ _05381_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16052_ _08143_ _08145_ VGND VGND VPWR VPWR _08146_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13264_ net43 _05475_ _05476_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_23_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15003_ spi0.data_packed\[7\] top0.periodTop\[7\] _07125_ VGND VGND VPWR VPWR _07127_
+ sky130_fd_sc_hd__mux2_1
X_13195_ _05425_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19811_ _11535_ _11536_ _11654_ VGND VGND VPWR VPWR _11691_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_31_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_31_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_102_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19742_ _11619_ _11610_ _11625_ VGND VGND VPWR VPWR _11626_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_198_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16954_ top0.currT_r\[9\] _08997_ top0.matmul0.beta_pass\[9\] VGND VGND VPWR VPWR
+ _09011_ sky130_fd_sc_hd__a21bo_1
X_15905_ _07928_ _07962_ _07999_ VGND VGND VPWR VPWR _08000_ sky130_fd_sc_hd__o21ai_4
X_19673_ net186 net180 VGND VGND VPWR VPWR _11560_ sky130_fd_sc_hd__nor2_4
X_16885_ top0.matmul0.beta_pass\[5\] _08946_ VGND VGND VPWR VPWR _08947_ sky130_fd_sc_hd__xnor2_1
X_18624_ _10579_ VGND VGND VPWR VPWR _10602_ sky130_fd_sc_hd__inv_2
X_15836_ _07838_ _07842_ _07931_ VGND VGND VPWR VPWR _07932_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_32_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18555_ _10529_ _10532_ VGND VGND VPWR VPWR _10534_ sky130_fd_sc_hd__nand2_1
X_15767_ _07861_ _07863_ VGND VGND VPWR VPWR _07864_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17506_ net390 VGND VGND VPWR VPWR _09493_ sky130_fd_sc_hd__inv_2
X_14718_ net25 _05619_ VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__nand2_1
X_18486_ net320 net381 VGND VGND VPWR VPWR _10466_ sky130_fd_sc_hd__nand2_1
X_15698_ top0.pid_q.out\[0\] top0.pid_q.curr_int\[0\] VGND VGND VPWR VPWR _07796_
+ sky130_fd_sc_hd__nand2_1
X_17437_ _09380_ _09422_ _09423_ VGND VGND VPWR VPWR _09424_ sky130_fd_sc_hd__a21oi_2
X_14649_ _06758_ _06788_ _06853_ VGND VGND VPWR VPWR _06854_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_170_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_16 _12812_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_27 net1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_38 net1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_166_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17368_ net353 VGND VGND VPWR VPWR _09355_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19107_ _11028_ _11077_ VGND VGND VPWR VPWR _11079_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16319_ _08406_ _08407_ VGND VGND VPWR VPWR _08409_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17299_ _09292_ _09288_ _09293_ VGND VGND VPWR VPWR _09294_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_41_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19038_ _10772_ _11010_ VGND VGND VPWR VPWR _11011_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21000_ net271 net251 VGND VGND VPWR VPWR _12847_ sky130_fd_sc_hd__xor2_2
XFILLER_0_195_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22951_ _02440_ _02462_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_50_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21902_ net145 net122 VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__nand2_2
X_25670_ top0.matmul0.sin\[9\] _04941_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__or2_2
X_22882_ _02374_ top0.svm0.tB\[12\] _02399_ _02400_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__o22a_1
X_24621_ _03315_ _03974_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21833_ _01178_ _01394_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24552_ _03760_ _03761_ _03906_ VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21764_ _01325_ _01301_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23503_ net1008 top0.matmul0.cos\[6\] _02915_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__mux2_1
X_27271_ clknet_3_7__leaf_clk_mosi _00885_ VGND VGND VPWR VPWR spi0.data_packed\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_20715_ _12561_ _12563_ _11673_ VGND VGND VPWR VPWR _12564_ sky130_fd_sc_hd__a21oi_1
X_24483_ _03820_ _03838_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21695_ _01247_ _01256_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26222_ spi0.data_packed\[9\] spi0.data_packed\[10\] net695 VGND VGND VPWR VPWR _05343_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23434_ _02869_ _02870_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20646_ net274 net263 VGND VGND VPWR VPWR _12495_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26153_ _05295_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__clkbuf_1
X_23365_ net216 _02806_ _11560_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20577_ _12355_ _12425_ VGND VGND VPWR VPWR _12426_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25104_ _04449_ _04451_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22316_ _01806_ _01875_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__nor2_1
X_26084_ top0.pid_d.out\[13\] _12031_ _05013_ spi0.data_packed\[77\] VGND VGND VPWR
+ VPWR _05265_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23296_ _11512_ _02742_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__nand2_1
X_25035_ _04382_ _04384_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__or2_1
X_22247_ net210 _01684_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22178_ _01684_ _01739_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__xnor2_1
X_21129_ _12915_ _12973_ _12917_ VGND VGND VPWR VPWR _12974_ sky130_fd_sc_hd__o21ba_1
X_26986_ clknet_leaf_27_clk_sys _00603_ net621 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[2\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout350 net351 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__buf_2
Xfanout361 top0.pid_d.mult0.b\[0\] VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__buf_4
XFILLER_0_108_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout372 top0.pid_d.mult0.a\[13\] VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkbuf_4
X_13951_ _06126_ _06127_ _06124_ _06125_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__a211o_1
X_25937_ top0.matmul0.alpha_pass\[15\] top0.matmul0.beta_pass\[15\] VGND VGND VPWR
+ VPWR _05150_ sky130_fd_sc_hd__xnor2_1
Xfanout383 net384 VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__buf_4
Xfanout394 top0.pid_d.mult0.a\[8\] VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__buf_2
X_13882_ _06094_ _05534_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__nor2_1
X_16670_ _08750_ _08754_ VGND VGND VPWR VPWR _08755_ sky130_fd_sc_hd__xnor2_1
X_25868_ _05031_ _05086_ _05087_ _05028_ net801 VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15621_ net477 net512 VGND VGND VPWR VPWR _07719_ sky130_fd_sc_hd__nand2_2
X_24819_ _04078_ _04086_ _04081_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_154_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25799_ _05027_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18340_ _10319_ _10321_ VGND VGND VPWR VPWR _10322_ sky130_fd_sc_hd__or2_1
X_15552_ net454 net536 VGND VGND VPWR VPWR _07651_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14503_ _06708_ _06709_ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__xor2_2
X_18271_ _09353_ _09364_ VGND VGND VPWR VPWR _10253_ sky130_fd_sc_hd__nor2_1
X_15483_ _07286_ _07291_ _07288_ VGND VGND VPWR VPWR _07582_ sky130_fd_sc_hd__o21a_1
XFILLER_0_189_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17222_ top0.pid_q.curr_int\[12\] _09140_ _09192_ _08679_ VGND VGND VPWR VPWR _09229_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14434_ _06639_ _06641_ VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14365_ _06565_ _06573_ VGND VGND VPWR VPWR _06574_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_4_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17153_ _09165_ _09166_ VGND VGND VPWR VPWR _09168_ sky130_fd_sc_hd__nand2_1
X_13316_ _05512_ _05516_ _05528_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__o21a_1
X_16104_ _08191_ _08196_ VGND VGND VPWR VPWR _08197_ sky130_fd_sc_hd__xnor2_1
X_17084_ net984 _09115_ _09118_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__a21o_1
X_14296_ _06425_ _06505_ VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16035_ _08123_ _08128_ VGND VGND VPWR VPWR _08129_ sky130_fd_sc_hd__xnor2_1
X_13247_ _05460_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17986_ _09971_ VGND VGND VPWR VPWR _09972_ sky130_fd_sc_hd__inv_2
X_19725_ net277 _11602_ VGND VGND VPWR VPWR _11609_ sky130_fd_sc_hd__nor2_1
X_16937_ net461 _08890_ _08995_ _08930_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19656_ _11531_ _11533_ _11534_ _11543_ VGND VGND VPWR VPWR _11544_ sky130_fd_sc_hd__a31o_1
X_16868_ top0.currT_r\[3\] _08917_ top0.matmul0.beta_pass\[3\] VGND VGND VPWR VPWR
+ _08931_ sky130_fd_sc_hd__a21bo_1
X_18607_ _10438_ _10580_ _10582_ VGND VGND VPWR VPWR _10586_ sky130_fd_sc_hd__o21ai_1
X_15819_ net499 _07914_ VGND VGND VPWR VPWR _07915_ sky130_fd_sc_hd__nand2_1
X_19587_ top0.cordic0.slte0.opA\[16\] top0.cordic0.slte0.opA\[17\] VGND VGND VPWR
+ VPWR _11476_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16799_ top0.kiq\[9\] _08863_ _08866_ VGND VGND VPWR VPWR _08873_ sky130_fd_sc_hd__and3_1
XFILLER_0_181_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18538_ _10514_ _10515_ VGND VGND VPWR VPWR _10517_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18469_ net317 _10447_ _10448_ _10208_ VGND VGND VPWR VPWR _10449_ sky130_fd_sc_hd__a22o_1
X_20500_ _11438_ _12142_ _12347_ _12348_ VGND VGND VPWR VPWR _12349_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21480_ _12968_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_16_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20431_ _12042_ _12127_ VGND VGND VPWR VPWR _12280_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_43_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23150_ top0.svm0.delta\[15\] _02636_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__nand2_1
X_20362_ _12209_ _12204_ _12205_ VGND VGND VPWR VPWR _12211_ sky130_fd_sc_hd__and3_1
XFILLER_0_141_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22101_ _01647_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23081_ _05735_ _02339_ _02538_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__and3_1
X_20293_ net290 net282 VGND VGND VPWR VPWR _12142_ sky130_fd_sc_hd__nand2_2
XFILLER_0_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22032_ _01177_ _01306_ _01593_ net146 VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26840_ clknet_leaf_46_clk_sys _00457_ net676 VGND VGND VPWR VPWR top0.svm0.counter\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_138_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23983_ _03337_ _03338_ _03339_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__and3_1
X_26771_ clknet_leaf_6_clk_sys _00388_ net590 VGND VGND VPWR VPWR top0.cordic0.cos\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22934_ _02306_ _02448_ _02309_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__a21o_1
X_25722_ top0.matmul0.sin\[7\] _04931_ net74 VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22865_ _02347_ top0.svm0.tB\[2\] _02383_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__o21a_1
X_25653_ net71 top0.matmul0.sin\[5\] VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24604_ _03957_ _03958_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__nand2_1
X_21816_ net135 _01338_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__xnor2_4
X_25584_ top0.matmul0.a\[14\] top0.matmul0.matmul_stage_inst.e\[14\] _04878_ VGND
+ VGND VPWR VPWR _04880_ sky130_fd_sc_hd__mux2_1
X_22796_ _02315_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24535_ _03060_ _03889_ _03801_ _03802_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21747_ net164 _01302_ _01305_ _01308_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__a211o_1
XFILLER_0_182_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24466_ _03572_ _03687_ _03689_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27254_ clknet_3_2__leaf_clk_mosi _00868_ VGND VGND VPWR VPWR spi0.data_packed\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21678_ _01234_ _01236_ _01239_ _01232_ _01233_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__o32a_1
XFILLER_0_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23417_ net215 _02687_ _11730_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26205_ _05334_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__clkbuf_1
X_20629_ _12277_ _12327_ net306 VGND VGND VPWR VPWR _12478_ sky130_fd_sc_hd__mux2_1
X_27185_ clknet_leaf_58_clk_sys _00799_ net644 VGND VGND VPWR VPWR top0.currT_r\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_24397_ _03676_ _03753_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14150_ _06360_ _06249_ _06361_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__o21a_1
X_26136_ spi0.data_packed\[31\] _05275_ _05277_ net802 VGND VGND VPWR VPWR _00812_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23348_ _02785_ _02791_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14081_ _06289_ _06292_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__xnor2_2
X_26067_ _05252_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__clkbuf_1
X_23279_ _02651_ _02726_ _11572_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__mux2_1
X_25018_ _04364_ _04367_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__xnor2_2
X_17840_ net329 net408 VGND VGND VPWR VPWR _09827_ sky130_fd_sc_hd__nand2_2
X_17771_ net375 net361 VGND VGND VPWR VPWR _09758_ sky130_fd_sc_hd__nand2_1
X_14983_ net171 VGND VGND VPWR VPWR _07115_ sky130_fd_sc_hd__inv_2
X_26969_ clknet_leaf_30_clk_sys _00586_ net623 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[1\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout180 top0.cordic0.gm0.iter\[4\] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_4
Xfanout191 net193 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_4
X_19510_ top0.pid_d.curr_int\[15\] top0.pid_d.prev_int\[15\] VGND VGND VPWR VPWR _11401_
+ sky130_fd_sc_hd__xor2_1
X_16722_ _08750_ _08754_ _08777_ _08801_ _08805_ VGND VGND VPWR VPWR _08806_ sky130_fd_sc_hd__o311a_1
X_13934_ net64 _05721_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19441_ top0.pid_d.curr_int\[7\] _11290_ _11293_ _11339_ VGND VGND VPWR VPWR _00333_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16653_ top0.pid_q.out\[13\] _07704_ VGND VGND VPWR VPWR _08739_ sky130_fd_sc_hd__nor2_1
X_13865_ _05957_ _06075_ _06077_ _05922_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15604_ top0.pid_q.state\[0\] net546 _07698_ VGND VGND VPWR VPWR _07703_ sky130_fd_sc_hd__or3_1
X_19372_ net884 _11285_ _11288_ top0.pid_d.curr_error\[5\] VGND VGND VPWR VPWR _00315_
+ sky130_fd_sc_hd__a22o_1
X_16584_ _08312_ _08589_ VGND VGND VPWR VPWR _08671_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13796_ _05999_ _06002_ _06008_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18323_ _10202_ _10220_ _10200_ VGND VGND VPWR VPWR _10305_ sky130_fd_sc_hd__o21a_1
X_15535_ _07556_ _07561_ _07633_ VGND VGND VPWR VPWR _07634_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18254_ _10131_ _10147_ _10133_ VGND VGND VPWR VPWR _10237_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15466_ net526 net464 VGND VGND VPWR VPWR _07565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17205_ top0.pid_q.curr_int\[10\] _09140_ _09213_ _09135_ VGND VGND VPWR VPWR _09214_
+ sky130_fd_sc_hd__a22o_1
X_14417_ _05500_ _05731_ VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18185_ net338 net376 VGND VGND VPWR VPWR _10168_ sky130_fd_sc_hd__nand2_2
XFILLER_0_170_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15397_ _07494_ _07495_ _07440_ VGND VGND VPWR VPWR _07496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17136_ top0.pid_q.curr_int\[2\] _09141_ _09152_ _09136_ VGND VGND VPWR VPWR _00215_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14348_ _06554_ _06556_ VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__xnor2_2
X_14279_ net45 _05723_ _05724_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__and3_1
X_17067_ net1018 _09107_ VGND VGND VPWR VPWR _09108_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16018_ _08110_ _08111_ VGND VGND VPWR VPWR _08112_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17969_ _09951_ _09954_ VGND VGND VPWR VPWR _09955_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19708_ _11592_ VGND VGND VPWR VPWR _11593_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20980_ _12817_ _12820_ VGND VGND VPWR VPWR _12827_ sky130_fd_sc_hd__or2_1
XFILLER_0_192_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19639_ net306 net300 VGND VGND VPWR VPWR _11527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22650_ _02143_ _02163_ _01948_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21601_ net105 net86 VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22581_ _02079_ _02134_ _02124_ _02086_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24320_ _03139_ _03141_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__and2_1
X_21532_ _01093_ _01088_ _01090_ _01091_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24251_ _03600_ _03605_ _03608_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21463_ _11759_ _01027_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23202_ net306 net300 net286 net277 net197 net188 VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__mux4_1
X_20414_ net302 _12262_ VGND VGND VPWR VPWR _12263_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24182_ _03505_ _03508_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_160_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21394_ net771 _12034_ _12037_ _00961_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__a31o_1
X_23133_ _02508_ _02598_ _02622_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__and3_1
X_20345_ _12163_ _12164_ VGND VGND VPWR VPWR _12194_ sky130_fd_sc_hd__or2_2
XFILLER_0_3_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23064_ net170 _02540_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__xor2_1
XFILLER_0_105_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20276_ net304 _12121_ _12124_ VGND VGND VPWR VPWR _12125_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22015_ _01296_ _01297_ _01575_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_78_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_78_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_26823_ clknet_leaf_37_clk_sys net709 net679 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfrtp_1
X_26754_ clknet_leaf_6_clk_sys _00371_ net591 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_23966_ _03121_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__clkbuf_4
X_25705_ top0.matmul0.sin\[2\] _04967_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__xnor2_1
X_22917_ net555 _06277_ net172 VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23897_ _03250_ _03106_ _03254_ _03252_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__o22a_1
X_26685_ clknet_leaf_62_clk_sys _00302_ net646 VGND VGND VPWR VPWR top0.pid_d.curr_error\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_22848_ top0.svm0.tA\[8\] _02366_ _02367_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__o21a_1
X_13650_ _05861_ _05862_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__xnor2_2
X_25636_ top0.matmul0.sin\[1\] top0.matmul0.sin\[0\] top0.matmul0.sin\[2\] top0.matmul0.sin\[3\]
+ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__or4_4
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13581_ _05710_ _05712_ _05793_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22779_ top0.svm0.counter\[4\] net170 _02299_ _02302_ VGND VGND VPWR VPWR _02303_
+ sky130_fd_sc_hd__or4_1
XFILLER_0_151_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25567_ top0.matmul0.a\[6\] top0.matmul0.matmul_stage_inst.e\[6\] _04867_ VGND VGND
+ VPWR VPWR _04871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15320_ net1026 net487 _07372_ VGND VGND VPWR VPWR _07419_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24518_ _03252_ _03825_ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25498_ top0.matmul0.matmul_stage_inst.mult1\[5\] _04154_ _04829_ VGND VGND VPWR
+ VPWR _04835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27237_ clknet_3_7__leaf_clk_mosi _00851_ VGND VGND VPWR VPWR spi0.data_packed\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_15251_ _07330_ _07332_ _07349_ VGND VGND VPWR VPWR _07350_ sky130_fd_sc_hd__nand3_1
XFILLER_0_191_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24449_ net570 net574 top0.matmul0.matmul_stage_inst.f\[15\] VGND VGND VPWR VPWR
+ _03805_ sky130_fd_sc_hd__o21ai_2
X_14202_ _06288_ _06293_ VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__and2_1
X_15182_ _07266_ _07280_ VGND VGND VPWR VPWR _07281_ sky130_fd_sc_hd__xnor2_4
X_27168_ clknet_leaf_32_clk_sys _00782_ net664 VGND VGND VPWR VPWR top0.periodTop_r\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_14133_ _06181_ _06203_ _06238_ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26119_ spi0.data_packed\[16\] _05279_ _05280_ net907 VGND VGND VPWR VPWR _00797_
+ sky130_fd_sc_hd__a22o_1
X_19990_ top0.cordic0.slte0.opA\[4\] _11857_ VGND VGND VPWR VPWR _11858_ sky130_fd_sc_hd__nor2_1
X_27099_ clknet_leaf_20_clk_sys _00716_ net610 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.a\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14064_ _06276_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__clkbuf_4
X_18941_ _10912_ _10915_ VGND VGND VPWR VPWR _10916_ sky130_fd_sc_hd__xnor2_1
X_18872_ _10723_ _10843_ _10844_ _10786_ _10846_ VGND VGND VPWR VPWR _10847_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_20_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17823_ _09684_ _09647_ VGND VGND VPWR VPWR _09810_ sky130_fd_sc_hd__and2b_1
Xhold3 top0.kpq\[13\] VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__dlygate4sd3_1
X_17754_ _09513_ _09456_ _09467_ VGND VGND VPWR VPWR _09741_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_6_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14966_ spi0.data_packed\[25\] top0.kiq\[9\] _07097_ VGND VGND VPWR VPWR _07105_
+ sky130_fd_sc_hd__mux2_1
X_16705_ _08787_ _08789_ VGND VGND VPWR VPWR _08790_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13917_ _05742_ _06129_ _05748_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__o21ai_4
X_17685_ net393 net345 VGND VGND VPWR VPWR _09672_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14897_ spi0.data_packed\[56\] top0.kpq\[8\] _07064_ VGND VGND VPWR VPWR _07069_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19424_ top0.pid_d.prev_int\[4\] _11318_ _11324_ VGND VGND VPWR VPWR _11325_ sky130_fd_sc_hd__o21a_1
XFILLER_0_162_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16636_ _08527_ _08721_ VGND VGND VPWR VPWR _08722_ sky130_fd_sc_hd__xnor2_2
X_13848_ _06053_ _06060_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19355_ net760 _11275_ _11281_ _11232_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16567_ net461 net466 VGND VGND VPWR VPWR _08654_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13779_ _05991_ _05987_ _05989_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__or3_1
X_18306_ net341 net369 VGND VGND VPWR VPWR _10288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15518_ net486 net508 VGND VGND VPWR VPWR _07617_ sky130_fd_sc_hd__nand2_2
X_19286_ _11227_ _11228_ VGND VGND VPWR VPWR _11229_ sky130_fd_sc_hd__nand2_1
X_16498_ _08582_ _08585_ VGND VGND VPWR VPWR _08586_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18237_ _10215_ _10219_ VGND VGND VPWR VPWR _10220_ sky130_fd_sc_hd__xnor2_2
X_15449_ _07273_ _07271_ _07278_ VGND VGND VPWR VPWR _07548_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18168_ _10042_ _10048_ VGND VGND VPWR VPWR _10152_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17119_ _07697_ net543 VGND VGND VPWR VPWR _09138_ sky130_fd_sc_hd__and2b_1
X_18099_ net421 net310 VGND VGND VPWR VPWR _10083_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20130_ top0.cordic0.slte0.opA\[14\] _11775_ VGND VGND VPWR VPWR _11986_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20061_ _11494_ net1013 _11921_ _11923_ VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23820_ _02985_ _02987_ _02979_ _02980_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__o22a_1
XFILLER_0_174_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23751_ _03105_ _03108_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__xnor2_2
X_20963_ _12739_ net1021 _12809_ VGND VGND VPWR VPWR _12811_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_174_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22702_ _02192_ _02251_ _02252_ _02195_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__o22ai_2
X_23682_ _02984_ _02986_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__or2_1
X_26470_ clknet_leaf_12_clk_sys _00101_ net618 VGND VGND VPWR VPWR top0.periodTop\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20894_ _11433_ _11648_ VGND VGND VPWR VPWR _12742_ sky130_fd_sc_hd__nor2_2
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25421_ _04663_ _04758_ _04756_ _04764_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__o22a_1
XFILLER_0_166_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22633_ _02140_ _02165_ _02185_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__o21ai_2
X_25352_ _04690_ _04696_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22564_ _02101_ _02118_ VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24303_ _03290_ _03287_ _03659_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21515_ _01074_ _01076_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__xnor2_2
X_25283_ _04541_ _04542_ _04540_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22495_ _02030_ _02034_ _02050_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24234_ _03565_ _03583_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27022_ clknet_leaf_16_clk_sys _00639_ net612 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_21446_ _01004_ _01010_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24165_ _03518_ _03519_ _03521_ _03513_ _03482_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__o221a_1
XFILLER_0_142_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21377_ net223 _12815_ _11789_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__a21o_1
X_23116_ net955 _02610_ _02611_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__a21o_1
X_20328_ _11787_ _12165_ VGND VGND VPWR VPWR _12177_ sky130_fd_sc_hd__xnor2_1
X_24096_ _03378_ _03453_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__xor2_2
XFILLER_0_31_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23047_ _02536_ _02537_ _02546_ _02547_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__a22o_1
X_20259_ net290 net284 VGND VGND VPWR VPWR _12108_ sky130_fd_sc_hd__nor2b_4
X_14820_ _07018_ _07013_ VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__or2b_1
X_26806_ clknet_leaf_70_clk_sys _00423_ net662 VGND VGND VPWR VPWR top0.pid_q.prev_int\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_24998_ _03496_ _03826_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14751_ net31 _06824_ VGND VGND VPWR VPWR _06953_ sky130_fd_sc_hd__nand2_1
X_26737_ clknet_leaf_101_clk_sys _00354_ net587 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_23949_ _03304_ _03305_ _03060_ _03306_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__a31o_1
X_13702_ _05657_ _05822_ _05588_ net64 VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17470_ _09375_ _09379_ _09373_ VGND VGND VPWR VPWR _09457_ sky130_fd_sc_hd__a21bo_1
X_14682_ _05626_ _06832_ _06884_ net25 _06885_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__o221a_1
XFILLER_0_168_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26668_ clknet_leaf_82_clk_sys _00285_ net647 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_16421_ net458 net501 VGND VGND VPWR VPWR _08510_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13633_ _05576_ _05845_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__xnor2_1
X_25619_ net746 _04896_ _04891_ _04901_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__o22a_1
XFILLER_0_184_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26599_ clknet_leaf_68_clk_sys _00222_ net662 VGND VGND VPWR VPWR top0.pid_q.curr_int\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19140_ net410 _11096_ _11105_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16352_ _08427_ _08441_ VGND VGND VPWR VPWR _08442_ sky130_fd_sc_hd__xnor2_2
X_13564_ _05773_ _05776_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_137_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15303_ net1026 net527 net495 net491 VGND VGND VPWR VPWR _07402_ sky130_fd_sc_hd__and4_1
XFILLER_0_137_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19071_ _11014_ _11042_ _11039_ VGND VGND VPWR VPWR _11043_ sky130_fd_sc_hd__o21a_1
X_13495_ _05700_ _05707_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__xnor2_1
X_16283_ _08371_ _08373_ VGND VGND VPWR VPWR _08374_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18022_ _10001_ _10006_ VGND VGND VPWR VPWR _10007_ sky130_fd_sc_hd__xnor2_2
X_15234_ _07176_ _07185_ VGND VGND VPWR VPWR _07333_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15165_ _07203_ _07208_ VGND VGND VPWR VPWR _07264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14116_ _06209_ _06326_ _06327_ _06215_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_50_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15096_ _07193_ _07194_ VGND VGND VPWR VPWR _07195_ sky130_fd_sc_hd__xor2_1
X_19973_ top0.cordic0.slte0.opA\[3\] _11785_ VGND VGND VPWR VPWR _11842_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18924_ _10897_ _10898_ VGND VGND VPWR VPWR _10899_ sky130_fd_sc_hd__and2b_1
X_14047_ _06258_ _06259_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__or2_2
XFILLER_0_66_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18855_ _10764_ _10830_ VGND VGND VPWR VPWR _10831_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17806_ net393 top0.pid_d.mult0.b\[4\] VGND VGND VPWR VPWR _09793_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18786_ _05449_ _10762_ VGND VGND VPWR VPWR _10763_ sky130_fd_sc_hd__and2_1
X_15998_ _08012_ _08037_ _08091_ VGND VGND VPWR VPWR _08092_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_94_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_167_Right_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17737_ _09719_ _09722_ _09723_ VGND VGND VPWR VPWR _09724_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14949_ spi0.data_packed\[17\] top0.kiq\[1\] _07086_ VGND VGND VPWR VPWR _07096_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17668_ _09610_ _09653_ _09654_ VGND VGND VPWR VPWR _09655_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_134_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19407_ _11307_ _11301_ _11302_ _11309_ VGND VGND VPWR VPWR _11310_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16619_ _08701_ _08704_ VGND VGND VPWR VPWR _08705_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17599_ net345 net426 _09585_ VGND VGND VPWR VPWR _09586_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_26_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_26_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19338_ _11273_ VGND VGND VPWR VPWR _11275_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19269_ _11125_ _11209_ _11212_ _11213_ _07800_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__o311a_1
XFILLER_0_5_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21300_ _13016_ _13103_ VGND VGND VPWR VPWR _13143_ sky130_fd_sc_hd__nand2_1
XFILLER_0_198_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22280_ net139 net123 _01217_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21231_ _12643_ _12618_ VGND VGND VPWR VPWR _13075_ sky130_fd_sc_hd__and2_1
Xhold200 top0.periodTop\[10\] VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold211 top0.pid_d.curr_int\[7\] VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold222 top0.currT_r\[12\] VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 top0.svm0.delta\[7\] VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold244 spi0.data_packed\[34\] VGND VGND VPWR VPWR net944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 top0.svm0.delta\[6\] VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21162_ _12998_ _13006_ VGND VGND VPWR VPWR _13007_ sky130_fd_sc_hd__xnor2_2
Xhold266 top0.b_in_matmul\[6\] VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 top0.pid_q.prev_int\[3\] VGND VGND VPWR VPWR net977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 top0.pid_q.prev_int\[10\] VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__dlygate4sd3_1
X_20113_ _11967_ _11970_ VGND VGND VPWR VPWR _11971_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold299 top0.cordic0.sin\[9\] VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout702 net29 VGND VGND VPWR VPWR net1030 sky130_fd_sc_hd__buf_4
X_25970_ top0.b_in_matmul\[2\] _05177_ _05165_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21093_ _12935_ _12937_ VGND VGND VPWR VPWR _12939_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24921_ _03198_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__buf_4
X_20044_ top0.cordic0.slte0.opA\[7\] _11895_ VGND VGND VPWR VPWR _11908_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24852_ _03313_ _03889_ _04099_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__a21o_1
X_23803_ _03149_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24783_ _04130_ _04135_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__xnor2_1
X_21995_ _01378_ _01392_ _01556_ _01372_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__o22a_2
X_26522_ clknet_leaf_66_clk_sys _00145_ net660 VGND VGND VPWR VPWR top0.pid_q.out\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_23734_ _03088_ _03089_ _03090_ _03091_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__o22a_2
X_20946_ _12784_ _12788_ _12789_ _12791_ _12793_ VGND VGND VPWR VPWR _12794_ sky130_fd_sc_hd__o221a_1
XFILLER_0_163_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26453_ clknet_leaf_55_clk_sys _00094_ net668 VGND VGND VPWR VPWR top0.kiq\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_23665_ net565 net557 top0.matmul0.matmul_stage_inst.e\[3\] VGND VGND VPWR VPWR _03023_
+ sky130_fd_sc_hd__o21a_1
X_20877_ _12724_ _12682_ _12725_ _12165_ VGND VGND VPWR VPWR _12726_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25404_ _04739_ _04747_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22616_ _02098_ _02119_ _02169_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__o21ai_2
X_26384_ clknet_leaf_41_clk_sys _00025_ net684 VGND VGND VPWR VPWR top0.svm0.tC\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_23596_ net76 _09278_ net559 VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25335_ _04675_ _04679_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22547_ net77 _01924_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_174_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13280_ top0.matmul0.alpha_pass\[2\] _05466_ _05474_ VGND VGND VPWR VPWR _05493_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25266_ _04570_ _04574_ _04611_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__o21ai_2
X_22478_ _02030_ _02034_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27005_ clknet_leaf_25_clk_sys _00622_ net627 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_24217_ _03561_ _03574_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21429_ _00984_ _00986_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__nor2_1
X_25197_ _04540_ _04543_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24148_ _03157_ _03060_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24079_ _03312_ _03321_ _03327_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__a21oi_1
X_16970_ _09025_ _09019_ top0.pid_q.prev_error\[10\] VGND VGND VPWR VPWR _09026_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_120_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15921_ _08014_ _08015_ VGND VGND VPWR VPWR _08016_ sky130_fd_sc_hd__xnor2_1
X_18640_ _10616_ _10617_ VGND VGND VPWR VPWR _10618_ sky130_fd_sc_hd__xnor2_1
X_15852_ net467 net515 VGND VGND VPWR VPWR _07948_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14803_ _06989_ _06994_ _07002_ _06935_ VGND VGND VPWR VPWR _07003_ sky130_fd_sc_hd__o22a_1
X_18571_ _10469_ _10478_ _10477_ VGND VGND VPWR VPWR _10550_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_118_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15783_ _07871_ _07879_ VGND VGND VPWR VPWR _07880_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17522_ _09424_ _09505_ VGND VGND VPWR VPWR _09509_ sky130_fd_sc_hd__or2_1
X_14734_ _06935_ _06936_ VGND VGND VPWR VPWR _06937_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17453_ _09379_ _09384_ VGND VGND VPWR VPWR _09440_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14665_ _06823_ _06826_ VGND VGND VPWR VPWR _06869_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16404_ _08142_ _08461_ VGND VGND VPWR VPWR _08493_ sky130_fd_sc_hd__nor2_1
X_13616_ _05578_ _05594_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__xor2_2
XFILLER_0_27_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17384_ net408 net347 VGND VGND VPWR VPWR _09371_ sky130_fd_sc_hd__nand2_1
X_14596_ _06800_ _06793_ VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19123_ _11093_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__clkbuf_1
X_16335_ _08421_ _08424_ VGND VGND VPWR VPWR _08425_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13547_ _05756_ _05759_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_42_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19054_ _10994_ _11026_ VGND VGND VPWR VPWR _11027_ sky130_fd_sc_hd__xnor2_2
X_16266_ net449 net516 VGND VGND VPWR VPWR _08357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13478_ _05686_ _05690_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_140_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18005_ _09986_ _09989_ VGND VGND VPWR VPWR _09990_ sky130_fd_sc_hd__xnor2_2
X_15217_ _07314_ _07315_ VGND VGND VPWR VPWR _07316_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16197_ net503 net497 _08288_ net473 VGND VGND VPWR VPWR _08289_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15148_ _07222_ _07245_ _07226_ net520 VGND VGND VPWR VPWR _07247_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19956_ net189 _11823_ _11807_ _11825_ VGND VGND VPWR VPWR _11826_ sky130_fd_sc_hd__a31o_1
X_15079_ net535 net465 VGND VGND VPWR VPWR _07178_ sky130_fd_sc_hd__nand2_1
X_18907_ net323 _10790_ net368 VGND VGND VPWR VPWR _10882_ sky130_fd_sc_hd__or3_1
X_19887_ _11728_ _11732_ _11740_ VGND VGND VPWR VPWR _11762_ sky130_fd_sc_hd__or3_1
X_18838_ net391 _09692_ _10228_ VGND VGND VPWR VPWR _10814_ sky130_fd_sc_hd__or3_2
XFILLER_0_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18769_ _10662_ _10663_ _10745_ VGND VGND VPWR VPWR _10746_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20800_ _12575_ _12578_ _12546_ VGND VGND VPWR VPWR _12649_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21780_ net129 net113 VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20731_ _12561_ _12563_ VGND VGND VPWR VPWR _12580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23450_ _01230_ _11519_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__nor2_1
X_20662_ _12465_ _12509_ VGND VGND VPWR VPWR _12511_ sky130_fd_sc_hd__nand2_1
X_22401_ _01217_ _01917_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__or2_1
X_23381_ _11789_ _11629_ _02712_ _11560_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__a2bb2o_1
X_20593_ net298 _12057_ VGND VGND VPWR VPWR _12442_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25120_ _04467_ _04468_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22332_ _01886_ _01887_ _01890_ _01802_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25051_ _04331_ _04400_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__xnor2_1
X_22263_ _01769_ _01822_ net77 VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24002_ _03306_ _03303_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__xor2_2
X_21214_ _12660_ _12575_ VGND VGND VPWR VPWR _13058_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22194_ net149 _01751_ _01754_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_130_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21145_ _12988_ _12989_ _12699_ net231 _12814_ VGND VGND VPWR VPWR _12990_ sky130_fd_sc_hd__a221o_1
Xwire1 _11850_ VGND VGND VPWR VPWR net1012 sky130_fd_sc_hd__clkbuf_1
Xfanout510 top0.pid_q.mult0.a\[11\] VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__buf_4
Xfanout521 top0.pid_q.mult0.a\[7\] VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__buf_4
Xfanout532 net533 VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__clkbuf_2
X_25953_ _05164_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__clkbuf_4
X_21076_ net234 _12696_ VGND VGND VPWR VPWR _12922_ sky130_fd_sc_hd__nor2_1
Xfanout543 top0.pid_q.state\[5\] VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__clkbuf_4
Xfanout554 top0.pid_q.state\[1\] VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__buf_2
Xfanout565 top0.matmul0.matmul_stage_inst.state\[4\] VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__buf_2
X_24904_ _04252_ _03741_ _03742_ _04254_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__o22a_1
Xfanout576 net577 VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__buf_4
X_20027_ net201 _11612_ VGND VGND VPWR VPWR _11892_ sky130_fd_sc_hd__nor2_1
Xfanout587 net589 VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__clkbuf_4
X_25884_ _05088_ _05096_ _05101_ top0.matmul0.alpha_pass\[8\] _05436_ VGND VGND VPWR
+ VPWR _05102_ sky130_fd_sc_hd__o221ai_4
Xfanout598 net605 VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24835_ _04091_ _04092_ _04186_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__o21a_1
XFILLER_0_201_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24766_ _04116_ _04117_ _04111_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21978_ _01493_ _01531_ _01533_ _01536_ _01539_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__a32o_1
X_26505_ clknet_leaf_81_clk_sys _00128_ net638 VGND VGND VPWR VPWR top0.pid_d.prev_int\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_23717_ _03073_ _03074_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__and2_2
XFILLER_0_56_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20929_ _12126_ _12776_ net284 VGND VGND VPWR VPWR _12777_ sky130_fd_sc_hd__mux2_1
X_24697_ _03931_ _04050_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14450_ _06656_ _06657_ VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26436_ clknet_leaf_79_clk_sys _00077_ net632 VGND VGND VPWR VPWR top0.kid\[9\] sky130_fd_sc_hd__dfrtp_1
X_23648_ _03004_ _03005_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__nor2_4
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13401_ _05610_ _05613_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__xnor2_4
X_14381_ _06587_ _06589_ VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_14_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26367_ _05415_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23579_ _02956_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16120_ _08198_ _08212_ VGND VGND VPWR VPWR _08213_ sky130_fd_sc_hd__xnor2_1
X_25318_ _04651_ _04652_ _04662_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_187_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13332_ _05544_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__buf_6
XFILLER_0_36_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26298_ spi0.data_packed\[47\] spi0.data_packed\[48\] net697 VGND VGND VPWR VPWR
+ _05381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16051_ _08055_ _08057_ _08144_ VGND VGND VPWR VPWR _08145_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_33_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25249_ _04525_ _04528_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13263_ top0.matmul0.beta_pass\[4\] _05434_ _05470_ _05463_ top0.c_out_calc\[4\]
+ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15002_ _07126_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13194_ spi0.opcode\[1\] spi0.opcode\[5\] _05423_ _05424_ VGND VGND VPWR VPWR _05425_
+ sky130_fd_sc_hd__nand4_4
X_19810_ _11680_ _11683_ _11673_ VGND VGND VPWR VPWR _11690_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16953_ _08882_ _09002_ _09009_ _09010_ _08889_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__o311a_1
X_19741_ net277 _11602_ _11619_ _11584_ net286 VGND VGND VPWR VPWR _11625_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_60_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15904_ _07928_ _07962_ _07930_ VGND VGND VPWR VPWR _07999_ sky130_fd_sc_hd__a21bo_1
X_19672_ _11422_ _11557_ _11558_ net84 VGND VGND VPWR VPWR _11559_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16884_ _08944_ top0.currT_r\[4\] _08945_ VGND VGND VPWR VPWR _08946_ sky130_fd_sc_hd__a21o_1
XFILLER_0_189_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18623_ _10579_ _10600_ _10421_ _10507_ VGND VGND VPWR VPWR _10601_ sky130_fd_sc_hd__o211a_1
X_15835_ _07838_ _07842_ _07839_ VGND VGND VPWR VPWR _07931_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_154_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18554_ _10529_ _10532_ VGND VGND VPWR VPWR _10533_ sky130_fd_sc_hd__nor2_1
X_15766_ _07749_ _07750_ _07862_ VGND VGND VPWR VPWR _07863_ sky130_fd_sc_hd__o21a_1
X_17505_ _09480_ _09491_ VGND VGND VPWR VPWR _09492_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14717_ net34 _06351_ VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__nand2_1
X_18485_ net327 net376 VGND VGND VPWR VPWR _10465_ sky130_fd_sc_hd__nand2_2
X_15697_ _07712_ _07794_ VGND VGND VPWR VPWR _07795_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17436_ net333 net422 net427 net330 VGND VGND VPWR VPWR _09423_ sky130_fd_sc_hd__a22oi_1
X_14648_ _06758_ _06788_ _06785_ VGND VGND VPWR VPWR _06853_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_17 top0.periodTop_r\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 net496 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17367_ net407 _09353_ VGND VGND VPWR VPWR _09354_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_39 net1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14579_ _06759_ _06784_ VGND VGND VPWR VPWR _06785_ sky130_fd_sc_hd__xor2_2
X_19106_ _11037_ _11028_ _11077_ VGND VGND VPWR VPWR _11078_ sky130_fd_sc_hd__or3_1
X_16318_ _08406_ _08407_ VGND VGND VPWR VPWR _08408_ sky130_fd_sc_hd__nand2_1
X_17298_ _09292_ _09288_ top0.matmul0.matmul_stage_inst.mult1\[7\] VGND VGND VPWR
+ VPWR _09293_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19037_ _11008_ _11009_ VGND VGND VPWR VPWR _11010_ sky130_fd_sc_hd__xor2_2
XFILLER_0_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16249_ net468 net473 net477 VGND VGND VPWR VPWR _08340_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_189_Left_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19939_ net195 _11410_ VGND VGND VPWR VPWR _11810_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22950_ _02306_ _02462_ _02309_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__a21o_1
X_21901_ net151 net130 _01135_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__a21o_1
X_22881_ top0.svm0.tB\[11\] _02398_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24620_ _03972_ _03973_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__nand2_2
X_21832_ _01392_ _01393_ net163 VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24551_ _03502_ _03758_ _03760_ _03761_ VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__a22o_1
X_21763_ net166 net158 VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20714_ _12560_ _12562_ _12559_ VGND VGND VPWR VPWR _12563_ sky130_fd_sc_hd__o21ai_1
X_23502_ _02916_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__clkbuf_1
X_27270_ clknet_3_6__leaf_clk_mosi _00884_ VGND VGND VPWR VPWR spi0.data_packed\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_24482_ _03835_ _03837_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__xnor2_2
X_21694_ _01252_ _01254_ _01255_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26221_ _05342_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__clkbuf_1
X_20645_ net263 _12490_ _12493_ VGND VGND VPWR VPWR _12494_ sky130_fd_sc_hd__mux2_1
X_23433_ top0.cordic0.vec\[1\]\[14\] _02858_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23364_ _02687_ _02688_ _11654_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__mux2_1
X_26152_ _05294_ top0.cordic0.slte0.opB\[5\] _12006_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__mux2_1
X_20576_ _12259_ _12421_ _12423_ _12424_ VGND VGND VPWR VPWR _12425_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25103_ _04449_ _04451_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22315_ _01738_ _01739_ _01684_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__mux2_1
X_23295_ _02659_ _02669_ _02730_ _02731_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__or4_1
X_26083_ _05264_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25034_ _04262_ _04266_ _04383_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__o21a_1
X_22246_ _01684_ _01737_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22177_ _01737_ _01738_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__nand2_1
X_21128_ net255 _12785_ VGND VGND VPWR VPWR _12973_ sky130_fd_sc_hd__nor2_1
X_26985_ clknet_leaf_27_clk_sys _00602_ net621 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout340 net342 VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout351 top0.pid_d.mult0.b\[2\] VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__clkbuf_4
Xfanout362 net367 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__buf_4
X_13950_ _06155_ _06160_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__xnor2_1
X_25936_ net916 _05028_ _05031_ _05149_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__a22o_1
Xfanout373 top0.pid_d.mult0.a\[13\] VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_4
X_21059_ net262 _12208_ VGND VGND VPWR VPWR _12905_ sky130_fd_sc_hd__nand2_1
Xfanout384 top0.pid_d.mult0.a\[10\] VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__buf_2
Xfanout395 net397 VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__buf_2
XFILLER_0_198_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13881_ net41 VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__inv_1
X_25867_ _05082_ _05085_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__or2_1
X_15620_ _07636_ _07658_ _07717_ VGND VGND VPWR VPWR _07718_ sky130_fd_sc_hd__a21o_1
X_24818_ _04088_ _04123_ _04169_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_201_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25798_ _05024_ _05026_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15551_ net457 net531 VGND VGND VPWR VPWR _07650_ sky130_fd_sc_hd__nand2_1
X_24749_ _04098_ _04101_ VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14502_ net31 _05639_ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__nand2_2
XFILLER_0_167_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18270_ _10165_ _10250_ _10251_ VGND VGND VPWR VPWR _10252_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15482_ _07575_ _07580_ VGND VGND VPWR VPWR _07581_ sky130_fd_sc_hd__xnor2_1
X_17221_ net551 _09050_ _09227_ net553 VGND VGND VPWR VPWR _09228_ sky130_fd_sc_hd__a22o_1
X_14433_ net30 _06640_ _06583_ _05579_ net33 VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__a32o_1
XFILLER_0_181_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26419_ clknet_leaf_60_clk_sys _00060_ net650 VGND VGND VPWR VPWR top0.kpq\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17152_ _09165_ _09166_ VGND VGND VPWR VPWR _09167_ sky130_fd_sc_hd__or2_1
X_14364_ _06567_ _06572_ VGND VGND VPWR VPWR _06573_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16103_ _08192_ _08195_ VGND VGND VPWR VPWR _08196_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_135_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13315_ _05512_ _05516_ _05527_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17083_ top0.pid_q.curr_error\[0\] _00011_ _09117_ VGND VGND VPWR VPWR _09118_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14295_ _06429_ _06430_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16034_ _08124_ _08127_ VGND VGND VPWR VPWR _08128_ sky130_fd_sc_hd__xnor2_1
X_13246_ top0.matmul0.state\[0\] top0.matmul0.start VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__nand2_4
XFILLER_0_126_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17985_ _09960_ _09970_ VGND VGND VPWR VPWR _09971_ sky130_fd_sc_hd__xnor2_1
X_16936_ top0.pid_q.state\[3\] _08987_ _08994_ _08882_ VGND VGND VPWR VPWR _08995_
+ sky130_fd_sc_hd__a211o_1
X_19724_ net273 VGND VGND VPWR VPWR _11608_ sky130_fd_sc_hd__inv_6
XFILLER_0_189_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16867_ net483 _08890_ _08929_ _08930_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__o211a_1
X_19655_ _11540_ _11542_ VGND VGND VPWR VPWR _11543_ sky130_fd_sc_hd__xor2_2
XFILLER_0_189_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15818_ net496 net492 VGND VGND VPWR VPWR _07914_ sky130_fd_sc_hd__xor2_4
X_18606_ _10443_ VGND VGND VPWR VPWR _10585_ sky130_fd_sc_hd__inv_2
X_19586_ top0.cordic0.slte0.opB\[11\] top0.cordic0.slte0.opA\[11\] VGND VGND VPWR
+ VPWR _11475_ sky130_fd_sc_hd__and2b_1
X_16798_ net1028 _08856_ _08859_ net827 _08872_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__a221o_1
XFILLER_0_189_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18537_ _10514_ _10515_ VGND VGND VPWR VPWR _10516_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15749_ _07182_ _07840_ _07844_ _07845_ VGND VGND VPWR VPWR _07846_ sky130_fd_sc_hd__o211a_1
XFILLER_0_176_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18468_ net385 net317 VGND VGND VPWR VPWR _10448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17419_ _09391_ _09405_ VGND VGND VPWR VPWR _09406_ sky130_fd_sc_hd__or2_1
X_18399_ _10369_ _10379_ VGND VGND VPWR VPWR _10380_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20430_ _12056_ _12278_ VGND VGND VPWR VPWR _12279_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_67_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20361_ _12204_ _12205_ _12209_ VGND VGND VPWR VPWR _12210_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22100_ _01646_ _01648_ _01661_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23080_ _05735_ _02580_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20292_ _12096_ _12140_ _11672_ VGND VGND VPWR VPWR _12141_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_197_Left_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22031_ _01592_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26770_ clknet_leaf_4_clk_sys _00387_ net580 VGND VGND VPWR VPWR top0.cordic0.cos\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_23982_ _03337_ _03338_ _03339_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__a21o_1
X_25721_ net792 _04964_ _04913_ _04978_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__a22o_1
X_22933_ _02446_ _02447_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__or2b_1
XFILLER_0_98_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25652_ _04926_ _04927_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__nand2_1
X_22864_ _02352_ top0.svm0.tB\[1\] top0.svm0.tB\[2\] _02347_ _02382_ VGND VGND VPWR
+ VPWR _02383_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24603_ _03954_ _03956_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__or2_1
X_21815_ net135 net122 VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25583_ _04879_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22795_ _02313_ top0.svm0.tA\[15\] VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24534_ _03888_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__clkbuf_4
X_21746_ net154 _01306_ _01307_ net159 VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27253_ clknet_3_2__leaf_clk_mosi _00867_ VGND VGND VPWR VPWR spi0.data_packed\[39\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_74_clk_sys clknet_3_5__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_74_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_109_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24465_ _03740_ _03744_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21677_ _11444_ _01237_ _01238_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__and3_1
XFILLER_0_188_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26204_ spi0.data_packed\[0\] spi0.data_packed\[1\] net694 VGND VGND VPWR VPWR _05334_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23416_ net103 _02853_ _02854_ _02852_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20628_ _12473_ _12464_ VGND VGND VPWR VPWR _12477_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27184_ clknet_leaf_59_clk_sys _00798_ net644 VGND VGND VPWR VPWR top0.currT_r\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_24396_ _03751_ _03752_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26135_ spi0.data_packed\[30\] _05275_ _05277_ top0.currT_r\[14\] VGND VGND VPWR
+ VPWR _00811_ sky130_fd_sc_hd__a22o_1
X_20559_ _12170_ _12407_ VGND VGND VPWR VPWR _12408_ sky130_fd_sc_hd__xnor2_2
X_23347_ _02788_ _02790_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__xor2_4
XFILLER_0_184_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14080_ _06290_ _06291_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__xor2_1
X_26066_ net985 _05251_ _05230_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23278_ net286 net278 net272 net265 net204 net196 VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__mux4_1
X_25017_ _04365_ _04366_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__xnor2_1
X_22229_ net77 _01785_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_201_Left_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17770_ net424 net319 VGND VGND VPWR VPWR _09757_ sky130_fd_sc_hd__nand2_1
X_14982_ top0.start_svm _07113_ VGND VGND VPWR VPWR _07114_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26968_ clknet_leaf_30_clk_sys _00585_ net623 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout170 top0.svm0.counter\[7\] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout181 top0.cordic0.gm0.iter\[4\] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_4
X_16721_ _08803_ _08804_ _08749_ VGND VGND VPWR VPWR _08805_ sky130_fd_sc_hd__mux2_1
Xfanout192 net193 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_195_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13933_ _06144_ _06145_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25919_ _08899_ _05129_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__nor2_1
X_26899_ clknet_leaf_108_clk_sys _00516_ net581 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19440_ top0.pid_d.state\[5\] _10508_ _11338_ net442 _11189_ VGND VGND VPWR VPWR
+ _11339_ sky130_fd_sc_hd__a221o_1
X_16652_ _08690_ _08737_ VGND VGND VPWR VPWR _08738_ sky130_fd_sc_hd__xnor2_2
X_13864_ _05878_ _06076_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15603_ _07697_ _07701_ VGND VGND VPWR VPWR _07702_ sky130_fd_sc_hd__nor2_1
XFILLER_0_201_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19371_ net878 _11285_ _11288_ top0.pid_d.curr_error\[4\] VGND VGND VPWR VPWR _00314_
+ sky130_fd_sc_hd__a22o_1
X_16583_ _08588_ _08590_ _08669_ VGND VGND VPWR VPWR _08670_ sky130_fd_sc_hd__a21oi_2
X_13795_ _06004_ _06007_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18322_ _10270_ _10303_ VGND VGND VPWR VPWR _10304_ sky130_fd_sc_hd__xnor2_1
X_15534_ _07556_ _07561_ _07554_ VGND VGND VPWR VPWR _07633_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18253_ _10222_ _10235_ VGND VGND VPWR VPWR _10236_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15465_ _07549_ _07563_ VGND VGND VPWR VPWR _07564_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17204_ net554 _09211_ _09212_ _09023_ VGND VGND VPWR VPWR _09213_ sky130_fd_sc_hd__a31o_1
X_14416_ net39 _05625_ VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18184_ _10151_ _10152_ _10166_ VGND VGND VPWR VPWR _10167_ sky130_fd_sc_hd__a21o_1
X_15396_ net472 _07407_ VGND VGND VPWR VPWR _07495_ sky130_fd_sc_hd__nor2_1
X_17135_ net543 _07895_ _09151_ net553 _08913_ VGND VGND VPWR VPWR _09152_ sky130_fd_sc_hd__a221o_1
X_14347_ _06487_ _06530_ _06555_ VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_163_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17066_ _09016_ top0.pid_q.curr_error\[10\] _09096_ VGND VGND VPWR VPWR _09107_ sky130_fd_sc_hd__mux2_1
X_14278_ net51 _05721_ VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__nand2_2
XFILLER_0_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16017_ net467 net510 VGND VGND VPWR VPWR _08111_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13229_ _05450_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17968_ _09848_ _09952_ _09953_ VGND VGND VPWR VPWR _09954_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19707_ net277 VGND VGND VPWR VPWR _11592_ sky130_fd_sc_hd__inv_2
X_16919_ _08977_ _08978_ VGND VGND VPWR VPWR _08979_ sky130_fd_sc_hd__nand2_1
X_17899_ _09754_ _09755_ _09775_ VGND VGND VPWR VPWR _09886_ sky130_fd_sc_hd__and3_1
X_19638_ _11430_ VGND VGND VPWR VPWR _11526_ sky130_fd_sc_hd__buf_4
XFILLER_0_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19569_ top0.cordic0.slte0.opA\[3\] _11456_ VGND VGND VPWR VPWR _11458_ sky130_fd_sc_hd__nor2_1
X_21600_ _01141_ _01145_ _01161_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22580_ _02123_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21531_ net148 net141 VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__or2b_1
XFILLER_0_16_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24250_ _03603_ _03602_ _03606_ _03553_ _03607_ VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21462_ _01026_ _12764_ _12770_ net231 VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_161_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20413_ net275 _12108_ VGND VGND VPWR VPWR _12262_ sky130_fd_sc_hd__xnor2_4
X_23201_ net297 net291 net272 net266 net197 net188 VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__mux4_1
X_24181_ _03455_ _03525_ _03534_ _03538_ VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__a31o_1
X_21393_ _00959_ _00960_ _12740_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__a21oi_1
X_23132_ _02483_ _02622_ _02596_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__o21ai_1
X_20344_ _12187_ _12192_ VGND VGND VPWR VPWR _12193_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23063_ net42 top0.svm0.counter\[9\] VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__xor2_1
XFILLER_0_144_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20275_ net283 _12100_ _12122_ _12123_ VGND VGND VPWR VPWR _12124_ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22014_ _01296_ _01297_ _01575_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26822_ clknet_leaf_38_clk_sys net705 net677 VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26753_ clknet_leaf_93_clk_sys _00370_ net591 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_98_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23965_ _03120_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__clkbuf_4
X_25704_ _04884_ _04905_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__or2_1
X_22916_ top0.svm0.calc_ready _02297_ _02433_ net706 _02309_ VGND VGND VPWR VPWR _00441_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_169_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26684_ clknet_leaf_62_clk_sys _00301_ net646 VGND VGND VPWR VPWR top0.pid_d.curr_error\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_23896_ _03251_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25635_ net859 _04904_ _04911_ _04913_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22847_ top0.svm0.counter\[8\] VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13580_ _05790_ _05792_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__xor2_1
X_25566_ _04870_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__clkbuf_1
X_22778_ _02300_ _02301_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24517_ _03869_ _03870_ _03871_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__o21a_1
X_21729_ net131 net126 VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__nand2_1
X_25497_ _04834_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27236_ clknet_3_7__leaf_clk_mosi _00850_ VGND VGND VPWR VPWR spi0.data_packed\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_15250_ _07333_ _07343_ _07348_ VGND VGND VPWR VPWR _07349_ sky130_fd_sc_hd__a21o_1
X_24448_ _03800_ _03803_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14201_ _06409_ _06410_ _06310_ VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_163_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27167_ clknet_leaf_32_clk_sys _00781_ net618 VGND VGND VPWR VPWR top0.periodTop_r\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_15181_ _07271_ _07279_ VGND VGND VPWR VPWR _07280_ sky130_fd_sc_hd__xnor2_4
X_24379_ _03133_ _03226_ _03225_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_2_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14132_ _06303_ _06343_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__xnor2_4
X_26118_ net737 _05279_ _05280_ net24 VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__a22o_1
XFILLER_0_201_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27098_ clknet_leaf_20_clk_sys _00715_ net609 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.a\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14063_ top0.svm0.state\[1\] top0.svm0.state\[0\] VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__or2_1
X_18940_ _10836_ _10913_ _10914_ VGND VGND VPWR VPWR _10915_ sky130_fd_sc_hd__o21ai_2
X_26049_ top0.matmul0.alpha_pass\[4\] _05237_ _05238_ VGND VGND VPWR VPWR _05239_
+ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18871_ _10786_ _10844_ _10806_ _10845_ VGND VGND VPWR VPWR _10846_ sky130_fd_sc_hd__a211o_1
XFILLER_0_101_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17822_ _09756_ _09808_ VGND VGND VPWR VPWR _09809_ sky130_fd_sc_hd__xnor2_2
Xhold4 net4 VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14965_ _07104_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__clkbuf_1
X_17753_ _09724_ _09738_ _09739_ VGND VGND VPWR VPWR _09740_ sky130_fd_sc_hd__a21o_1
X_13916_ _05743_ _05744_ _05745_ _05746_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__a2bb2oi_1
X_16704_ _08788_ VGND VGND VPWR VPWR _08789_ sky130_fd_sc_hd__inv_2
X_17684_ net399 net342 VGND VGND VPWR VPWR _09671_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14896_ _07068_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16635_ net498 _08720_ VGND VGND VPWR VPWR _08721_ sky130_fd_sc_hd__and2_1
X_19423_ top0.pid_d.prev_int\[4\] _11318_ top0.pid_d.curr_int\[4\] VGND VGND VPWR
+ VPWR _11324_ sky130_fd_sc_hd__a21o_1
X_13847_ _06056_ _06059_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16566_ _08643_ _08652_ VGND VGND VPWR VPWR _08653_ sky130_fd_sc_hd__xor2_2
X_19354_ net931 _11275_ _11281_ _11223_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__a22o_1
X_13778_ _05985_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18305_ _10172_ _10180_ _10181_ VGND VGND VPWR VPWR _10287_ sky130_fd_sc_hd__o21ai_2
X_15517_ _07532_ _07615_ VGND VGND VPWR VPWR _07616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19285_ top0.pid_d.prev_error\[11\] top0.pid_d.curr_error\[11\] VGND VGND VPWR VPWR
+ _11228_ sky130_fd_sc_hd__xnor2_1
X_16497_ _08527_ _08584_ VGND VGND VPWR VPWR _08585_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_139_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18236_ _10216_ _10218_ VGND VGND VPWR VPWR _10219_ sky130_fd_sc_hd__xnor2_1
X_15448_ _07533_ _07534_ _07545_ VGND VGND VPWR VPWR _07547_ sky130_fd_sc_hd__a21o_1
XFILLER_0_182_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18167_ _10039_ _10050_ _10150_ VGND VGND VPWR VPWR _10151_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_25_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15379_ net537 _07477_ VGND VGND VPWR VPWR _07478_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17118_ top0.pid_q.curr_int\[0\] top0.pid_q.prev_int\[0\] VGND VGND VPWR VPWR _09137_
+ sky130_fd_sc_hd__xor2_1
X_18098_ _10080_ _10081_ VGND VGND VPWR VPWR _10082_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17049_ _05448_ _08855_ VGND VGND VPWR VPWR _09099_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20060_ _11494_ _11922_ VGND VGND VPWR VPWR _11923_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_22_clk_sys clknet_3_2__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_22_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_116_Left_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23750_ _03106_ _03107_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__nor2_1
X_20962_ _12739_ net1021 _12809_ VGND VGND VPWR VPWR _12810_ sky130_fd_sc_hd__or3_1
XFILLER_0_68_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22701_ _02194_ _02219_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23681_ _02997_ _02999_ _02976_ _02977_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__o22a_1
X_20893_ net732 _12034_ _12037_ _12741_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__a31o_1
X_25420_ _04763_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__inv_2
X_22632_ _02140_ _02165_ _02166_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_165_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25351_ _04691_ _04695_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22563_ _02116_ _02117_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__xor2_1
XFILLER_0_119_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24302_ _03290_ _03287_ _03294_ _03293_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__o211a_1
X_21514_ net114 _01075_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__xnor2_4
X_25282_ _04546_ _04551_ _04627_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_125_Left_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22494_ _02030_ _02034_ _02011_ VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27021_ clknet_leaf_18_clk_sys _00638_ net614 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24233_ _03565_ _03576_ _03577_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__and3_1
X_21445_ _01004_ _01010_ _12815_ _12926_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_160_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24164_ _03513_ _03521_ _03482_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__o21ba_1
X_21376_ _00941_ _00943_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__xnor2_2
X_23115_ _02478_ _02598_ _02609_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__and3_1
X_20327_ _12150_ _12151_ _12166_ _12175_ VGND VGND VPWR VPWR _12176_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24095_ _03451_ _03409_ _03452_ _03415_ _03422_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__o221a_1
X_23046_ net26 top0.svm0.counter\[14\] _02543_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__or3b_1
X_20258_ net305 net290 VGND VGND VPWR VPWR _12107_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_134_Left_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20189_ net245 net237 VGND VGND VPWR VPWR _12038_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26805_ clknet_leaf_70_clk_sys _00422_ net658 VGND VGND VPWR VPWR top0.pid_q.prev_int\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24997_ _04336_ _04346_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__xor2_4
X_14750_ _06926_ _06932_ VGND VGND VPWR VPWR _06952_ sky130_fd_sc_hd__nand2_2
X_26736_ clknet_leaf_101_clk_sys _00353_ net587 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_23948_ _02994_ _02996_ _03076_ _03077_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__o22a_1
XFILLER_0_169_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13701_ net67 _05579_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__nand2_1
X_14681_ _05626_ _06760_ net20 VGND VGND VPWR VPWR _06885_ sky130_fd_sc_hd__a21o_1
X_26667_ clknet_leaf_82_clk_sys _00284_ net647 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_23879_ _03235_ _03236_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__xnor2_4
X_16420_ _08420_ _08425_ _08508_ VGND VGND VPWR VPWR _08509_ sky130_fd_sc_hd__a21o_1
X_13632_ _05564_ _05570_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__xor2_1
X_25618_ net70 top0.matmul0.cos\[12\] VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26598_ clknet_leaf_67_clk_sys _00221_ net661 VGND VGND VPWR VPWR top0.pid_q.curr_int\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_183_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16351_ _08429_ _08440_ VGND VGND VPWR VPWR _08441_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13563_ _05774_ _05775_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__xnor2_1
X_25549_ _04861_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_143_Left_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15302_ net527 net495 net491 net1026 VGND VGND VPWR VPWR _07401_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19070_ _11016_ _11038_ _11040_ VGND VGND VPWR VPWR _11042_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_180_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16282_ _08272_ _08273_ _08372_ VGND VGND VPWR VPWR _08373_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_125_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13494_ _05703_ _05706_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18021_ _10003_ _10005_ VGND VGND VPWR VPWR _10006_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15233_ _07238_ _07331_ VGND VGND VPWR VPWR _07332_ sky130_fd_sc_hd__xnor2_2
X_27219_ clknet_3_1__leaf_clk_mosi _00833_ VGND VGND VPWR VPWR spi0.data_packed\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_151_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15164_ _07255_ _07262_ VGND VGND VPWR VPWR _07263_ sky130_fd_sc_hd__xnor2_1
X_14115_ net24 _05894_ _05497_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19972_ _11431_ _11840_ net177 VGND VGND VPWR VPWR _11841_ sky130_fd_sc_hd__o21ai_1
X_15095_ net540 net457 VGND VGND VPWR VPWR _07194_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14046_ _06085_ _06130_ _06136_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__a21oi_1
X_18923_ _10894_ _10896_ VGND VGND VPWR VPWR _10898_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_152_Left_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18854_ _10828_ _10829_ VGND VGND VPWR VPWR _10830_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17805_ net388 net346 VGND VGND VPWR VPWR _09792_ sky130_fd_sc_hd__nand2_1
X_15997_ _08012_ _08037_ _08026_ VGND VGND VPWR VPWR _08091_ sky130_fd_sc_hd__a21bo_1
X_18785_ net437 _09339_ _10754_ _10761_ VGND VGND VPWR VPWR _10762_ sky130_fd_sc_hd__a31o_1
XFILLER_0_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17736_ _09505_ _09507_ _09719_ _09722_ VGND VGND VPWR VPWR _09723_ sky130_fd_sc_hd__o2bb2a_1
X_14948_ _07095_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__clkbuf_1
X_17667_ _09609_ _09612_ VGND VGND VPWR VPWR _09654_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14879_ _07059_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19406_ top0.pid_d.curr_int\[2\] VGND VGND VPWR VPWR _11309_ sky130_fd_sc_hd__inv_2
XFILLER_0_187_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16618_ _08702_ _08703_ VGND VGND VPWR VPWR _08704_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17598_ net422 net349 VGND VGND VPWR VPWR _09585_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_161_Left_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16549_ _08561_ _08562_ _08635_ VGND VGND VPWR VPWR _08636_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_128_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19337_ _11274_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19268_ net326 _11094_ VGND VGND VPWR VPWR _11213_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18219_ _10114_ _10125_ _10201_ VGND VGND VPWR VPWR _10202_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19199_ top0.matmul0.alpha_pass\[3\] _11141_ VGND VGND VPWR VPWR _11150_ sky130_fd_sc_hd__or2_2
XFILLER_0_170_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21230_ _13066_ _13067_ _13069_ _13073_ VGND VGND VPWR VPWR _13074_ sky130_fd_sc_hd__o31a_1
XFILLER_0_5_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold201 top0.cordic0.slte0.opA\[0\] VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _00124_ VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold223 top0.pid_d.curr_error\[8\] VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__dlygate4sd3_1
X_21161_ _13004_ _13005_ VGND VGND VPWR VPWR _13006_ sky130_fd_sc_hd__or2b_1
Xhold234 top0.currT_r\[3\] VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _05368_ VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_170_Left_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold256 spi0.data_packed\[42\] VGND VGND VPWR VPWR net956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold267 spi0.data_packed\[39\] VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold278 top0.pid_d.curr_int\[12\] VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__dlygate4sd3_1
X_20112_ _11515_ _11968_ _11969_ VGND VGND VPWR VPWR _11970_ sky130_fd_sc_hd__a21o_1
Xhold289 top0.svm0.tA\[9\] VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__dlygate4sd3_1
X_21092_ _12935_ _12937_ VGND VGND VPWR VPWR _12938_ sky130_fd_sc_hd__and2_1
Xfanout703 net117 VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24920_ _03006_ _03826_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20043_ net181 _11906_ VGND VGND VPWR VPWR _11907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24851_ _04199_ _04202_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23802_ _03021_ _03031_ _03159_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__o21a_2
X_24782_ _04039_ _04134_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__nor2_2
X_21994_ _01319_ _01378_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__xnor2_1
X_26521_ clknet_leaf_66_clk_sys _00144_ net660 VGND VGND VPWR VPWR top0.pid_q.out\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_23733_ net567 net558 top0.matmul0.matmul_stage_inst.e\[11\] VGND VGND VPWR VPWR
+ _03091_ sky130_fd_sc_hd__o21a_4
XFILLER_0_200_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20945_ _12792_ _12791_ VGND VGND VPWR VPWR _12793_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26452_ clknet_leaf_55_clk_sys _00093_ net668 VGND VGND VPWR VPWR top0.kiq\[9\] sky130_fd_sc_hd__dfrtp_1
X_23664_ net569 net573 top0.matmul0.matmul_stage_inst.f\[3\] VGND VGND VPWR VPWR _03022_
+ sky130_fd_sc_hd__o21a_1
X_20876_ net235 top0.cordic0.vec\[0\]\[15\] net214 _12236_ VGND VGND VPWR VPWR _12725_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_152_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25403_ _04742_ _04746_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22615_ _02098_ _02119_ _02120_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__a21o_1
X_26383_ clknet_leaf_42_clk_sys _00024_ net684 VGND VGND VPWR VPWR top0.svm0.tC\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23595_ _02964_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25334_ _04676_ _04678_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22546_ _02060_ _02068_ _02099_ _01948_ _02100_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__a221o_2
XFILLER_0_107_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25265_ _04570_ _04574_ _04568_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__a21o_1
X_22477_ _02033_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__inv_2
X_27004_ clknet_leaf_28_clk_sys _00621_ net622 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_24216_ _03571_ _03573_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21428_ _00958_ _00925_ _00991_ _13154_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__and4b_2
X_25196_ _04541_ _04542_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24147_ _03503_ _03504_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__nor2_2
XFILLER_0_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21359_ _00918_ _00923_ _13188_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__a21o_1
X_24078_ _03266_ _03435_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__xnor2_4
X_23029_ _02530_ _02526_ top0.svm0.delta\[15\] VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__mux2_1
X_15920_ net453 net523 VGND VGND VPWR VPWR _08015_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15851_ net536 _07649_ _07838_ _07946_ _07837_ VGND VGND VPWR VPWR _07947_ sky130_fd_sc_hd__o32a_1
X_14802_ _06989_ _06993_ _07001_ _06949_ VGND VGND VPWR VPWR _07002_ sky130_fd_sc_hd__o22a_1
X_18570_ _10541_ _10548_ VGND VGND VPWR VPWR _10549_ sky130_fd_sc_hd__xnor2_2
X_15782_ _07876_ _07878_ VGND VGND VPWR VPWR _07879_ sky130_fd_sc_hd__xor2_1
X_14733_ _06919_ _06933_ VGND VGND VPWR VPWR _06936_ sky130_fd_sc_hd__nor2_1
X_17521_ _09505_ _09507_ _09413_ VGND VGND VPWR VPWR _09508_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26719_ clknet_leaf_81_clk_sys _00336_ net634 VGND VGND VPWR VPWR top0.pid_d.curr_int\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17452_ _09373_ _09375_ VGND VGND VPWR VPWR _09439_ sky130_fd_sc_hd__or2b_1
X_14664_ _06823_ _06826_ VGND VGND VPWR VPWR _06868_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16403_ _08413_ _08463_ _08464_ VGND VGND VPWR VPWR _08492_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13615_ _05815_ _05821_ _05827_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_157_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17383_ net412 net343 VGND VGND VPWR VPWR _09370_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14595_ _06749_ _06791_ VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_184_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16334_ _08422_ _08423_ VGND VGND VPWR VPWR _08424_ sky130_fd_sc_hd__xnor2_1
X_19122_ _05449_ _11092_ VGND VGND VPWR VPWR _11093_ sky130_fd_sc_hd__and2_1
X_13546_ _05757_ _05758_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__xor2_2
XFILLER_0_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19053_ _10996_ _11025_ VGND VGND VPWR VPWR _11026_ sky130_fd_sc_hd__xor2_1
X_16265_ net453 net1029 VGND VGND VPWR VPWR _08356_ sky130_fd_sc_hd__nand2_1
X_13477_ _05687_ _05689_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18004_ _09987_ _09988_ VGND VGND VPWR VPWR _09989_ sky130_fd_sc_hd__xor2_1
X_15216_ net522 net491 VGND VGND VPWR VPWR _07315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16196_ net476 _08287_ VGND VGND VPWR VPWR _08288_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15147_ _07230_ _07225_ _07222_ VGND VGND VPWR VPWR _07246_ sky130_fd_sc_hd__a21o_1
XFILLER_0_168_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19955_ _11824_ net189 net195 net1016 VGND VGND VPWR VPWR _11825_ sky130_fd_sc_hd__and4b_1
X_15078_ net537 net462 VGND VGND VPWR VPWR _07177_ sky130_fd_sc_hd__nand2_1
X_14029_ _06161_ _06240_ _06241_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__a21oi_1
X_18906_ _10790_ net362 _10712_ VGND VGND VPWR VPWR _10881_ sky130_fd_sc_hd__nor3_1
X_19886_ _11714_ _11634_ _11760_ net83 VGND VGND VPWR VPWR _11761_ sky130_fd_sc_hd__a2bb2o_2
X_18837_ net387 _10811_ _10812_ VGND VGND VPWR VPWR _10813_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_93_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18768_ _10662_ _10663_ _10658_ VGND VGND VPWR VPWR _10745_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_89_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17719_ net383 VGND VGND VPWR VPWR _09706_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18699_ _10608_ _10675_ VGND VGND VPWR VPWR _10677_ sky130_fd_sc_hd__and2_1
X_20730_ _12575_ _12578_ VGND VGND VPWR VPWR _12579_ sky130_fd_sc_hd__or2_1
XFILLER_0_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20661_ _12465_ _12509_ VGND VGND VPWR VPWR _12510_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22400_ _01217_ _01917_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20592_ _12059_ _12264_ VGND VGND VPWR VPWR _12441_ sky130_fd_sc_hd__nor2_1
X_23380_ net116 _02820_ _02821_ _02819_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22331_ _01888_ _01889_ _01742_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25050_ _04334_ _04399_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__xor2_1
X_22262_ _01820_ _01821_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24001_ _03353_ _03358_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21213_ _13054_ _13055_ _13056_ VGND VGND VPWR VPWR _13057_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22193_ net126 _01456_ _01752_ _01753_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__a31o_1
XFILLER_0_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21144_ net242 _11739_ VGND VGND VPWR VPWR _12989_ sky130_fd_sc_hd__nand2_1
Xfanout500 net502 VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__buf_4
Xfanout511 net512 VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__clkbuf_4
Xfanout522 net524 VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21075_ _12908_ _12920_ VGND VGND VPWR VPWR _12921_ sky130_fd_sc_hd__xnor2_2
Xfanout533 top0.pid_q.mult0.a\[3\] VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__buf_4
X_25952_ _05163_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__buf_2
Xfanout544 net545 VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__clkbuf_4
Xfanout555 top0.svm0.delta\[0\] VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__buf_2
X_24903_ _04252_ _04253_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__nand2_1
Xfanout566 net567 VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__clkbuf_4
X_20026_ net201 net185 _11574_ _11890_ VGND VGND VPWR VPWR _11891_ sky130_fd_sc_hd__a211o_1
Xfanout577 net606 VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__buf_4
X_25883_ _05088_ _05095_ _05100_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__o21a_1
Xfanout588 net589 VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__clkbuf_4
Xfanout599 net600 VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__clkbuf_4
X_24834_ _04091_ _04092_ _04090_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_197_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24765_ _04111_ _04116_ _04117_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__and3_1
X_21977_ _01537_ _01538_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26504_ clknet_leaf_84_clk_sys net829 net633 VGND VGND VPWR VPWR top0.pid_d.prev_int\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23716_ _03065_ _03072_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__or2_1
X_20928_ net261 net267 VGND VGND VPWR VPWR _12776_ sky130_fd_sc_hd__or2b_1
X_24696_ _03946_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26435_ clknet_leaf_79_clk_sys _00076_ net632 VGND VGND VPWR VPWR top0.kid\[8\] sky130_fd_sc_hd__dfrtp_1
X_23647_ net574 top0.matmul0.matmul_stage_inst.d\[5\] top0.matmul0.matmul_stage_inst.c\[5\]
+ net558 VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__a22o_4
XFILLER_0_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20859_ net251 _12039_ _12707_ _12255_ _12085_ VGND VGND VPWR VPWR _12708_ sky130_fd_sc_hd__a221o_2
XFILLER_0_36_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13400_ net56 _05611_ _05612_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__and3_2
XFILLER_0_138_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14380_ _06517_ _06519_ _06588_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_148_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26366_ spi0.opcode\[1\] spi0.opcode\[2\] net691 VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__mux2_1
X_23578_ top0.b_in_matmul\[12\] top0.matmul0.b\[12\] _02948_ VGND VGND VPWR VPWR _02956_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25317_ _04651_ _04652_ _04650_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__o21a_1
X_13331_ top0.matmul0.beta_pass\[7\] _05434_ _05469_ _05463_ top0.c_out_calc\[7\]
+ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__a32o_1
XFILLER_0_135_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22529_ _02009_ _02044_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__nand2_1
X_26297_ _05380_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16050_ _08055_ _08057_ _08053_ VGND VGND VPWR VPWR _08144_ sky130_fd_sc_hd__a21bo_1
X_25248_ _04586_ _04594_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__xnor2_1
X_13262_ top0.matmul0.alpha_pass\[4\] _05466_ _05474_ VGND VGND VPWR VPWR _05475_
+ sky130_fd_sc_hd__nand3_2
XFILLER_0_122_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15001_ spi0.data_packed\[6\] top0.periodTop\[6\] _07125_ VGND VGND VPWR VPWR _07126_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25179_ _04457_ _04458_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__or2_1
X_13193_ spi0.opcode\[0\] spi0.opcode\[2\] spi0.opcode\[3\] spi0.opcode\[4\] VGND
+ VGND VPWR VPWR _05424_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19740_ _11622_ _11623_ _11586_ _11587_ _11609_ VGND VGND VPWR VPWR _11624_ sky130_fd_sc_hd__a2111o_1
X_16952_ net459 _08861_ VGND VGND VPWR VPWR _09010_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_69_clk_sys clknet_3_5__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_69_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15903_ _07905_ _07996_ _07997_ VGND VGND VPWR VPWR _07998_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19671_ top0.cordic0.gm0.iter\[1\] net200 net187 VGND VGND VPWR VPWR _11558_ sky130_fd_sc_hd__and3_1
X_16883_ _08944_ top0.currT_r\[4\] _08917_ top0.currT_r\[3\] _08931_ VGND VGND VPWR
+ VPWR _08945_ sky130_fd_sc_hd__o221a_1
X_18622_ _10439_ _10504_ _10440_ VGND VGND VPWR VPWR _10600_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_189_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15834_ _07847_ _07859_ _07929_ VGND VGND VPWR VPWR _07930_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18553_ _10530_ _10531_ net364 VGND VGND VPWR VPWR _10532_ sky130_fd_sc_hd__o21a_1
X_15765_ _07749_ _07750_ _07759_ VGND VGND VPWR VPWR _07862_ sky130_fd_sc_hd__a21o_1
X_17504_ _09481_ _09490_ VGND VGND VPWR VPWR _09491_ sky130_fd_sc_hd__xnor2_1
X_14716_ _06896_ _06918_ VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_197_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18484_ _10445_ _10463_ VGND VGND VPWR VPWR _10464_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15696_ _07792_ _07793_ VGND VGND VPWR VPWR _07794_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14647_ _06820_ _06851_ VGND VGND VPWR VPWR _06852_ sky130_fd_sc_hd__xor2_2
X_17435_ net330 net333 net422 net425 VGND VGND VPWR VPWR _09422_ sky130_fd_sc_hd__nand4_1
XFILLER_0_131_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_18 top0.pid_d.state\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14578_ _06773_ _06783_ VGND VGND VPWR VPWR _06784_ sky130_fd_sc_hd__xnor2_2
XANTENNA_29 net513 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17366_ _09352_ VGND VGND VPWR VPWR _09353_ sky130_fd_sc_hd__clkbuf_4
X_19105_ _11074_ _11076_ VGND VGND VPWR VPWR _11077_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_103_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13529_ _05730_ _05741_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_137_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16317_ top0.pid_q.out\[9\] top0.pid_q.curr_int\[9\] VGND VGND VPWR VPWR _08407_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17297_ top0.matmul0.matmul_stage_inst.mult2\[7\] VGND VGND VPWR VPWR _09292_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16248_ _08277_ _08279_ _08338_ VGND VGND VPWR VPWR _08339_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_113_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19036_ net356 net360 net316 _10948_ VGND VGND VPWR VPWR _11009_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16179_ net458 net510 VGND VGND VPWR VPWR _08271_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19938_ _11807_ _11808_ net195 VGND VGND VPWR VPWR _11809_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19869_ net237 _11514_ _11717_ VGND VGND VPWR VPWR _11745_ sky130_fd_sc_hd__mux2_1
X_21900_ _01457_ _01461_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__nor2_1
X_22880_ top0.svm0.tB\[11\] _02398_ _02345_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__o21a_1
X_21831_ _01372_ _01392_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__nand2_2
XFILLER_0_78_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24550_ _03901_ _03904_ VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__xnor2_2
X_21762_ _01320_ _01268_ _01323_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23501_ top0.cordic0.cos\[5\] top0.matmul0.cos\[5\] _02915_ VGND VGND VPWR VPWR _02916_
+ sky130_fd_sc_hd__mux2_1
X_20713_ net285 net273 _12277_ _12552_ _12555_ VGND VGND VPWR VPWR _12562_ sky130_fd_sc_hd__o311a_1
X_24481_ _03694_ _03697_ _03836_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_77_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21693_ _01249_ _01253_ _01250_ _01165_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_18_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26220_ spi0.data_packed\[8\] spi0.data_packed\[9\] net694 VGND VGND VPWR VPWR _05342_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23432_ top0.cordic0.vec\[1\]\[14\] _02858_ _02861_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_19_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20644_ _11550_ _12491_ _12492_ _12347_ VGND VGND VPWR VPWR _12493_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26151_ spi0.data_packed\[3\] _05293_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__xnor2_1
X_23363_ net120 _02804_ _02805_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__a21bo_1
X_20575_ _12251_ _12257_ _12422_ VGND VGND VPWR VPWR _12424_ sky130_fd_sc_hd__nand3_1
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25102_ _04363_ _04375_ _04450_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__a21oi_1
X_22314_ _01807_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26082_ top0.a_in_matmul\[12\] _05263_ _05164_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__mux2_1
X_23294_ net220 _11594_ _02740_ _11425_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__a22o_2
XFILLER_0_14_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25033_ _04262_ _04266_ _04264_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22245_ _01804_ _01805_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__nand2_2
XFILLER_0_131_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22176_ _01732_ _01735_ _01736_ _01729_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_44_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21127_ net251 _12785_ VGND VGND VPWR VPWR _12972_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26984_ clknet_leaf_30_clk_sys _00601_ net621 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult2\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout330 net331 VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_4
Xfanout341 net342 VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_70_clk_sys clknet_3_5__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_70_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
Xfanout352 net354 VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__buf_2
X_25935_ _05145_ _05148_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout363 net367 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_2
X_21058_ net259 _12900_ _12901_ _12903_ VGND VGND VPWR VPWR _12904_ sky130_fd_sc_hd__o2bb2a_1
Xfanout374 net376 VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__buf_4
Xfanout385 net386 VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__buf_2
Xfanout396 net397 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__clkbuf_4
X_20009_ _11512_ _11874_ VGND VGND VPWR VPWR _11875_ sky130_fd_sc_hd__nand2_1
X_13880_ _06090_ _06091_ _06088_ _06089_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__a211o_2
X_25866_ _05082_ _05085_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__nand2_1
X_24817_ _04088_ _04123_ _04089_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_119_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25797_ top0.cordic0.out_valid _05022_ top0.cordic_done VGND VGND VPWR VPWR _05026_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_202_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15550_ net448 net540 VGND VGND VPWR VPWR _07649_ sky130_fd_sc_hd__nand2_1
X_24748_ _04099_ _04100_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_189_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14501_ net36 _05625_ VGND VGND VPWR VPWR _06708_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15481_ _07576_ _07579_ VGND VGND VPWR VPWR _07580_ sky130_fd_sc_hd__xnor2_1
X_24679_ _03924_ _03921_ _03922_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_167_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14432_ _05588_ VGND VGND VPWR VPWR _06640_ sky130_fd_sc_hd__buf_2
X_17220_ _09225_ _09226_ VGND VGND VPWR VPWR _09227_ sky130_fd_sc_hd__xnor2_1
X_26418_ clknet_leaf_60_clk_sys _00059_ net650 VGND VGND VPWR VPWR top0.kpq\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17151_ top0.pid_q.curr_int\[4\] top0.pid_q.prev_int\[4\] VGND VGND VPWR VPWR _09166_
+ sky130_fd_sc_hd__xor2_1
X_14363_ _06568_ _06571_ VGND VGND VPWR VPWR _06572_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26349_ _05406_ VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__clkbuf_1
X_16102_ _08193_ _08194_ VGND VGND VPWR VPWR _08195_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13314_ _05519_ _05526_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__xnor2_4
X_17082_ _09116_ VGND VGND VPWR VPWR _09117_ sky130_fd_sc_hd__buf_2
XFILLER_0_80_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14294_ _06398_ _06502_ _06503_ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_12_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16033_ _08125_ _08126_ VGND VGND VPWR VPWR _08127_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13245_ _05459_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17984_ _09961_ _09969_ VGND VGND VPWR VPWR _09970_ sky130_fd_sc_hd__xor2_1
X_19723_ net175 _11593_ _11606_ _11607_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__a31o_1
XFILLER_0_165_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16935_ net550 _08992_ _08993_ VGND VGND VPWR VPWR _08994_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19654_ _11484_ _11504_ _11509_ _11541_ VGND VGND VPWR VPWR _11542_ sky130_fd_sc_hd__a211o_1
X_16866_ net1019 VGND VGND VPWR VPWR _08930_ sky130_fd_sc_hd__buf_2
X_18605_ _10505_ _10583_ _10581_ VGND VGND VPWR VPWR _10584_ sky130_fd_sc_hd__a21o_1
X_15817_ net469 net515 _07911_ _07912_ VGND VGND VPWR VPWR _07913_ sky130_fd_sc_hd__a31o_1
Xclkbuf_3_2__f_clk_sys clknet_0_clk_sys VGND VGND VPWR VPWR clknet_3_2__leaf_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_19585_ top0.cordic0.slte0.opA\[10\] top0.cordic0.slte0.opB\[10\] VGND VGND VPWR
+ VPWR _11474_ sky130_fd_sc_hd__xor2_1
XFILLER_0_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16797_ top0.kiq\[8\] _08863_ _08866_ VGND VGND VPWR VPWR _08872_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18536_ top0.pid_d.out\[8\] top0.pid_d.curr_int\[8\] VGND VGND VPWR VPWR _10515_
+ sky130_fd_sc_hd__xnor2_1
X_15748_ _07839_ _07841_ VGND VGND VPWR VPWR _07845_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18467_ net385 net364 _10446_ _09494_ _09363_ VGND VGND VPWR VPWR _10447_ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15679_ _07775_ _07776_ VGND VGND VPWR VPWR _07777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17418_ _09393_ _09350_ _09404_ VGND VGND VPWR VPWR _09405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18398_ _10377_ _10378_ VGND VGND VPWR VPWR _10379_ sky130_fd_sc_hd__and2b_1
XFILLER_0_184_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17349_ _09333_ _09336_ VGND VGND VPWR VPWR _09337_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20360_ _12206_ _12208_ VGND VGND VPWR VPWR _12209_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19019_ _10982_ _10990_ _10991_ _10926_ VGND VGND VPWR VPWR _10992_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_114_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20291_ net252 net246 VGND VGND VPWR VPWR _12140_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22030_ _01372_ _01393_ net142 VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23981_ _02998_ _03000_ _03015_ _03016_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__o22a_1
X_25720_ top0.matmul0.sin\[7\] _04977_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__xnor2_1
X_22932_ _02444_ _02445_ _02443_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25651_ net73 _04920_ top0.matmul0.sin\[5\] VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__or3b_1
X_22863_ _02352_ top0.svm0.tB\[1\] top0.svm0.tB\[0\] _02298_ VGND VGND VPWR VPWR _02382_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24602_ _03954_ _03956_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21814_ _01362_ _01375_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__xnor2_1
X_25582_ top0.matmul0.a\[13\] top0.matmul0.matmul_stage_inst.e\[13\] _04878_ VGND
+ VGND VPWR VPWR _04879_ sky130_fd_sc_hd__mux2_1
X_22794_ _02313_ top0.svm0.tA\[15\] VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24533_ _03103_ _03104_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21745_ net154 _01093_ _01136_ net164 VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_leaf_9_clk_sys clknet_3_2__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_9_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_171_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_17_clk_sys clknet_3_2__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_17_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_27252_ clknet_3_2__leaf_clk_mosi _00866_ VGND VGND VPWR VPWR spi0.data_packed\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_24464_ _03701_ _03733_ _03819_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21676_ _01066_ _01113_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__nand2_1
X_26203_ _05333_ VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__clkbuf_1
X_23415_ net103 _11857_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__nor2_1
X_20627_ _12463_ _12475_ VGND VGND VPWR VPWR _12476_ sky130_fd_sc_hd__nand2_1
X_27183_ clknet_leaf_58_clk_sys _00797_ net643 VGND VGND VPWR VPWR top0.currT_r\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_24395_ _03679_ _03750_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__or2_1
XFILLER_0_163_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26134_ spi0.data_packed\[29\] _05281_ _05282_ top0.currT_r\[13\] VGND VGND VPWR
+ VPWR _00810_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23346_ _11512_ _02789_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__nand2_2
X_20558_ _12115_ _12116_ _12171_ _12403_ _12406_ VGND VGND VPWR VPWR _12407_ sky130_fd_sc_hd__o311a_1
XFILLER_0_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26065_ net1024 _05237_ _05250_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23277_ net150 _02721_ _02720_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__a21oi_2
X_20489_ net280 _12057_ _12337_ VGND VGND VPWR VPWR _12338_ sky130_fd_sc_hd__o21a_1
X_25016_ _03254_ _04288_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22228_ _11444_ _01787_ _01788_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__and3_1
X_22159_ _01698_ _01720_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14981_ top0.svm0.state\[1\] top0.svm0.state\[0\] VGND VGND VPWR VPWR _07113_ sky130_fd_sc_hd__nor2_1
X_26967_ clknet_leaf_15_clk_sys _00584_ net613 VGND VGND VPWR VPWR top0.matmul0.b\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout160 net161 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout171 net172 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_4
X_16720_ _08750_ _08802_ _08800_ VGND VGND VPWR VPWR _08804_ sky130_fd_sc_hd__a21oi_1
Xfanout182 net186 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_4
X_13932_ net51 _05639_ _05737_ _05624_ net56 VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__a32o_1
X_25918_ _05030_ _05132_ _05133_ _05028_ net939 VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__a32o_1
Xfanout193 top0.cordic0.gm0.iter\[1\] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26898_ clknet_leaf_107_clk_sys _00515_ net577 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13863_ _05905_ _05906_ _05879_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__mux2_1
X_16651_ _08735_ _08736_ VGND VGND VPWR VPWR _08737_ sky130_fd_sc_hd__nand2_1
X_25849_ top0.matmul0.alpha_pass\[7\] top0.matmul0.beta_pass\[7\] VGND VGND VPWR VPWR
+ _05070_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_201_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15602_ net548 _07700_ VGND VGND VPWR VPWR _07701_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19370_ net872 _11285_ _11288_ top0.pid_d.curr_error\[3\] VGND VGND VPWR VPWR _00313_
+ sky130_fd_sc_hd__a22o_1
X_13794_ _06005_ _06006_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__xnor2_1
X_16582_ _08588_ _08590_ _08587_ VGND VGND VPWR VPWR _08669_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18321_ _10301_ _10302_ VGND VGND VPWR VPWR _10303_ sky130_fd_sc_hd__or2b_1
X_15533_ _07572_ _07573_ _07631_ VGND VGND VPWR VPWR _07632_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_201_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18252_ _10233_ _10234_ VGND VGND VPWR VPWR _10235_ sky130_fd_sc_hd__and2b_1
X_15464_ _07554_ _07562_ VGND VGND VPWR VPWR _07563_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_38_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14415_ net36 _05602_ _05603_ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__and3_2
X_17203_ _09209_ _09210_ VGND VGND VPWR VPWR _09212_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18183_ _10151_ _10152_ _10149_ VGND VGND VPWR VPWR _10166_ sky130_fd_sc_hd__o21a_1
X_15395_ _07182_ net539 _07493_ VGND VGND VPWR VPWR _07494_ sky130_fd_sc_hd__nor3_1
XFILLER_0_80_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14346_ _06487_ _06530_ _06481_ VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__a21o_1
X_17134_ _09149_ _09150_ VGND VGND VPWR VPWR _09151_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17065_ _09106_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__clkbuf_1
X_14277_ _06482_ _06486_ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_52_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16016_ net458 net516 VGND VGND VPWR VPWR _08110_ sky130_fd_sc_hd__nand2_1
X_13228_ net553 _05449_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_29_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17967_ _09851_ _09854_ VGND VGND VPWR VPWR _09953_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19706_ net174 _11571_ _11590_ _11591_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__a31o_1
X_16918_ top0.pid_q.prev_error\[7\] top0.pid_q.curr_error\[7\] VGND VGND VPWR VPWR
+ _08978_ sky130_fd_sc_hd__xnor2_1
X_17898_ _09767_ _09773_ _09884_ VGND VGND VPWR VPWR _09885_ sky130_fd_sc_hd__o21a_2
X_19637_ net297 VGND VGND VPWR VPWR _11525_ sky130_fd_sc_hd__inv_2
X_16849_ net488 _08861_ VGND VGND VPWR VPWR _08914_ sky130_fd_sc_hd__or2_1
XFILLER_0_192_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_178_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19568_ top0.cordic0.slte0.opA\[3\] _11456_ VGND VGND VPWR VPWR _11457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18519_ net405 _10497_ _10498_ VGND VGND VPWR VPWR _10499_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_34_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19499_ top0.pid_d.curr_int\[13\] top0.pid_d.prev_int\[13\] VGND VGND VPWR VPWR _11391_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_186_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21530_ net146 _01090_ _01091_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21461_ _11727_ _12180_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23200_ _02650_ _02651_ _11572_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__mux2_1
X_20412_ _12245_ _12248_ _12260_ VGND VGND VPWR VPWR _12261_ sky130_fd_sc_hd__o21a_1
X_24180_ _03524_ _03535_ _03536_ _03537_ _03454_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21392_ net1021 _00958_ _00926_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__or3b_1
XFILLER_0_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23131_ top0.svm0.delta\[10\] _02619_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__or2_1
X_20343_ _12174_ _12181_ VGND VGND VPWR VPWR _12192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23062_ _02560_ _02561_ _02562_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_105_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20274_ net283 _12100_ _12102_ VGND VGND VPWR VPWR _12123_ sky130_fd_sc_hd__nor3_1
XFILLER_0_101_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_47_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22013_ _01090_ _01312_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26821_ clknet_leaf_36_clk_sys _00438_ net676 VGND VGND VPWR VPWR top0.svm0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_23964_ _03248_ _03217_ VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__nor2_1
X_26752_ clknet_leaf_94_clk_sys _00369_ net591 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_22915_ _02313_ top0.svm0.tC\[15\] _02432_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__o21ai_1
X_25703_ net887 _04964_ _04936_ _04966_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__a22o_1
X_26683_ clknet_leaf_62_clk_sys _00300_ net648 VGND VGND VPWR VPWR top0.pid_d.curr_error\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23895_ _03250_ _03106_ _03251_ _03252_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__or4_2
XFILLER_0_169_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22846_ _02361_ _02333_ _02362_ _02364_ _02365_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__a221o_1
X_25634_ _04912_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25565_ top0.matmul0.a\[5\] top0.matmul0.matmul_stage_inst.e\[5\] _04867_ VGND VGND
+ VPWR VPWR _04870_ sky130_fd_sc_hd__mux2_1
X_22777_ top0.svm0.counter\[9\] net169 top0.svm0.counter\[11\] top0.svm0.counter\[12\]
+ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__or4_1
XFILLER_0_137_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24516_ _03106_ _03198_ _03807_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21728_ net126 _01263_ _01138_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__a21o_1
XFILLER_0_192_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25496_ top0.matmul0.matmul_stage_inst.mult1\[4\] _04062_ _04829_ VGND VGND VPWR
+ VPWR _04834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24447_ _03801_ _03802_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27235_ clknet_3_7__leaf_clk_mosi _00849_ VGND VGND VPWR VPWR spi0.data_packed\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_21659_ net96 net78 VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_192_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14200_ _06409_ _06410_ VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15180_ _07273_ _07278_ VGND VGND VPWR VPWR _07279_ sky130_fd_sc_hd__xnor2_2
X_27166_ clknet_leaf_11_clk_sys _00780_ net601 VGND VGND VPWR VPWR top0.a_in_matmul\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24378_ _03701_ _03734_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_201_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14131_ _06341_ _06342_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__nor2_2
XFILLER_0_22_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26117_ net754 _05279_ _05280_ net1030 VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23329_ _02771_ _02773_ VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_132_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27097_ clknet_leaf_0_clk_sys _00714_ net586 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.a\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14062_ _06178_ _06274_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__xnor2_2
X_26048_ top0.pid_d.out\[4\] _05232_ _05233_ spi0.data_packed\[68\] VGND VGND VPWR
+ VPWR _05238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18870_ _10722_ VGND VGND VPWR VPWR _10845_ sky130_fd_sc_hd__clkbuf_4
X_17821_ _09775_ _09807_ VGND VGND VPWR VPWR _09808_ sky130_fd_sc_hd__xor2_1
XFILLER_0_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold5 _00439_ VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__dlygate4sd3_1
X_17752_ _09726_ _09737_ VGND VGND VPWR VPWR _09739_ sky130_fd_sc_hd__and2_1
X_14964_ spi0.data_packed\[24\] top0.kiq\[8\] _07097_ VGND VGND VPWR VPWR _07104_
+ sky130_fd_sc_hd__mux2_1
X_16703_ _08784_ _08786_ VGND VGND VPWR VPWR _08788_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13915_ _06124_ _06125_ _06126_ _06127_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__o211a_1
X_17683_ net388 net349 VGND VGND VPWR VPWR _09670_ sky130_fd_sc_hd__nand2_1
XFILLER_0_199_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14895_ spi0.data_packed\[55\] top0.kpq\[7\] _07064_ VGND VGND VPWR VPWR _07068_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19422_ top0.pid_d.curr_int\[4\] _11290_ _11293_ _11323_ VGND VGND VPWR VPWR _00330_
+ sky130_fd_sc_hd__a22o_1
X_16634_ _08654_ _08647_ _08719_ net459 VGND VGND VPWR VPWR _08720_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_18_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13846_ _06057_ _06058_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19353_ top0.pid_d.curr_error\[9\] _11275_ _11278_ _11212_ VGND VGND VPWR VPWR _00303_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16565_ _08650_ _08651_ VGND VGND VPWR VPWR _08652_ sky130_fd_sc_hd__and2b_1
X_13777_ _05985_ _05987_ _05989_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18304_ _10275_ _10285_ VGND VGND VPWR VPWR _10286_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15516_ _07527_ _07528_ _07531_ _07614_ VGND VGND VPWR VPWR _07615_ sky130_fd_sc_hd__a31o_1
XFILLER_0_183_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19284_ _11225_ _11216_ _11226_ VGND VGND VPWR VPWR _11227_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16496_ _08515_ _08517_ _08583_ VGND VGND VPWR VPWR _08584_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18235_ _10121_ _10123_ _10217_ VGND VGND VPWR VPWR _10218_ sky130_fd_sc_hd__o21a_1
X_15447_ _07533_ _07534_ _07545_ VGND VGND VPWR VPWR _07546_ sky130_fd_sc_hd__nand3_2
XFILLER_0_142_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18166_ _10040_ _10049_ VGND VGND VPWR VPWR _10150_ sky130_fd_sc_hd__nor2_1
XFILLER_0_167_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15378_ net535 net489 _07456_ VGND VGND VPWR VPWR _07477_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17117_ _09135_ VGND VGND VPWR VPWR _09136_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14329_ _06450_ _06451_ _06537_ VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__and3_1
X_18097_ net411 net315 VGND VGND VPWR VPWR _10081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17048_ _09098_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18999_ _10961_ _10971_ VGND VGND VPWR VPWR _10973_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20961_ _12806_ _12808_ VGND VGND VPWR VPWR _12809_ sky130_fd_sc_hd__xor2_2
XFILLER_0_139_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22700_ _02194_ _02219_ net79 VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23680_ _03036_ _03037_ _02993_ _02995_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__o22a_1
X_20892_ _12739_ _12740_ VGND VGND VPWR VPWR _12741_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22631_ _02182_ _02183_ _02171_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25350_ _04510_ _04694_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22562_ net80 _02067_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24301_ _03652_ _03654_ _03657_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21513_ net123 net118 VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__and2b_2
XFILLER_0_63_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25281_ _04546_ _04551_ _04544_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_119_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22493_ _12742_ _02047_ _02048_ _02049_ VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27020_ clknet_leaf_16_clk_sys _00637_ net612 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.f\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_24232_ _03586_ _03587_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21444_ _01008_ _01009_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__xor2_1
XFILLER_0_185_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24163_ _03509_ _03490_ _03498_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__or3_1
X_21375_ net218 _00942_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23114_ _02483_ _02609_ _02596_ VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20326_ net304 _12121_ _12124_ VGND VGND VPWR VPWR _12175_ sky130_fd_sc_hd__a21oi_2
X_24094_ _03419_ _03409_ _03451_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23045_ _02544_ _02545_ _06217_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__a21o_1
X_20257_ _12098_ _12099_ _12104_ VGND VGND VPWR VPWR _12106_ sky130_fd_sc_hd__nand3_1
X_20188_ _12036_ VGND VGND VPWR VPWR _12037_ sky130_fd_sc_hd__buf_6
XFILLER_0_192_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26804_ clknet_leaf_71_clk_sys _00421_ net658 VGND VGND VPWR VPWR top0.pid_q.prev_int\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_24996_ _04344_ _04345_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__or2_2
X_26735_ clknet_leaf_100_clk_sys _00352_ net587 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
X_23947_ _02985_ _02987_ _02976_ _02977_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__o22a_2
XFILLER_0_25_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13700_ _05910_ _05911_ _05912_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__a21o_1
X_14680_ _06832_ _05640_ net20 VGND VGND VPWR VPWR _06884_ sky130_fd_sc_hd__o21a_1
X_23878_ _03038_ _03039_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__xnor2_2
X_26666_ clknet_leaf_82_clk_sys _00283_ net647 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13631_ _05838_ _05842_ _05843_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__o21ai_2
X_22829_ _02347_ top0.svm0.tA\[2\] VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__nor2_1
X_25617_ net752 _04896_ _04891_ _04900_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__o22a_1
X_26597_ clknet_leaf_68_clk_sys _00220_ net662 VGND VGND VPWR VPWR top0.pid_q.curr_int\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13562_ _05573_ _05542_ _05544_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__or3_1
X_16350_ _08434_ _08439_ VGND VGND VPWR VPWR _08440_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25548_ top0.matmul0.b\[13\] top0.matmul0.matmul_stage_inst.f\[13\] _04856_ VGND
+ VGND VPWR VPWR _04861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_181_Right_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15301_ _07351_ _07352_ _07399_ VGND VGND VPWR VPWR _07400_ sky130_fd_sc_hd__a21o_1
X_16281_ _08272_ _08273_ _08271_ VGND VGND VPWR VPWR _08372_ sky130_fd_sc_hd__o21ba_1
X_25479_ _04762_ _04664_ _04821_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__a21o_1
X_13493_ _05535_ _05704_ _05705_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18020_ _09941_ _09946_ _10004_ VGND VGND VPWR VPWR _10005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15232_ _07186_ _07236_ VGND VGND VPWR VPWR _07331_ sky130_fd_sc_hd__xor2_1
X_27218_ clknet_3_1__leaf_clk_mosi _00832_ VGND VGND VPWR VPWR spi0.data_packed\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15163_ _07258_ _07261_ VGND VGND VPWR VPWR _07262_ sky130_fd_sc_hd__xnor2_1
X_27149_ clknet_leaf_31_clk_sys _00763_ net620 VGND VGND VPWR VPWR top0.b_in_matmul\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14114_ _06107_ _06322_ _06324_ _06047_ _06325_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19971_ _11836_ _11839_ VGND VGND VPWR VPWR _11840_ sky130_fd_sc_hd__xor2_1
X_15094_ _07177_ _07178_ _07192_ VGND VGND VPWR VPWR _07193_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14045_ _06085_ _06130_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__nor2_1
X_18922_ _10894_ _10896_ VGND VGND VPWR VPWR _10897_ sky130_fd_sc_hd__nor2_1
X_18853_ _10743_ _10747_ _10748_ VGND VGND VPWR VPWR _10829_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_24_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17804_ net384 net350 VGND VGND VPWR VPWR _09791_ sky130_fd_sc_hd__nand2_1
X_18784_ top0.pid_d.out\[10\] _07137_ _10760_ net432 VGND VGND VPWR VPWR _10761_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15996_ _08000_ _08061_ _08089_ VGND VGND VPWR VPWR _08090_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_173_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17735_ net357 _09720_ _09721_ _09495_ VGND VGND VPWR VPWR _09722_ sky130_fd_sc_hd__a22o_1
X_14947_ spi0.data_packed\[16\] top0.kiq\[0\] _07086_ VGND VGND VPWR VPWR _07095_
+ sky130_fd_sc_hd__mux2_1
X_17666_ _09609_ _09612_ VGND VGND VPWR VPWR _09653_ sky130_fd_sc_hd__nor2_1
X_14878_ spi0.data_packed\[79\] top0.kpd\[15\] _07053_ VGND VGND VPWR VPWR _07059_
+ sky130_fd_sc_hd__mux2_1
X_19405_ _11301_ _11302_ _11307_ VGND VGND VPWR VPWR _11308_ sky130_fd_sc_hd__a21o_1
X_16617_ net447 net504 VGND VGND VPWR VPWR _08703_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13829_ _05999_ _06008_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17597_ net423 net354 _09583_ _09525_ net359 VGND VGND VPWR VPWR _09584_ sky130_fd_sc_hd__a32o_1
XFILLER_0_175_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19336_ _11271_ top0.pid_d.curr_error\[0\] _11273_ VGND VGND VPWR VPWR _11274_ sky130_fd_sc_hd__mux2_1
X_16548_ _08561_ _08562_ _08563_ VGND VGND VPWR VPWR _08635_ sky130_fd_sc_hd__o21a_1
XFILLER_0_174_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19267_ _11120_ _11210_ _11211_ VGND VGND VPWR VPWR _11212_ sky130_fd_sc_hd__and3_1
XFILLER_0_169_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16479_ _08558_ _08566_ VGND VGND VPWR VPWR _08567_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18218_ _10114_ _10125_ _10112_ VGND VGND VPWR VPWR _10201_ sky130_fd_sc_hd__a21o_1
XFILLER_0_170_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19198_ net439 _11147_ _11148_ VGND VGND VPWR VPWR _11149_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18149_ _10009_ _10037_ _10132_ VGND VGND VPWR VPWR _10133_ sky130_fd_sc_hd__o21a_1
Xhold202 top0.svm0.calc_ready VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold213 top0.cordic0.slte0.opA\[10\] VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 top0.pid_q.curr_int\[8\] VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 top0.currT_r\[11\] VGND VGND VPWR VPWR net935 sky130_fd_sc_hd__dlygate4sd3_1
X_21160_ _13000_ _13003_ VGND VGND VPWR VPWR _13005_ sky130_fd_sc_hd__or2_1
Xhold246 spi0.data_packed\[40\] VGND VGND VPWR VPWR net946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 _05375_ VGND VGND VPWR VPWR net957 sky130_fd_sc_hd__dlygate4sd3_1
X_20111_ _11730_ _11519_ _11810_ VGND VGND VPWR VPWR _11969_ sky130_fd_sc_hd__and3_1
Xhold268 top0.pid_d.prev_int\[0\] VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_180_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold279 top0.a_in_matmul\[2\] VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__dlygate4sd3_1
X_21091_ _12865_ _12873_ _12936_ VGND VGND VPWR VPWR _12937_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20042_ _11410_ _11901_ _11902_ _11903_ _11905_ VGND VGND VPWR VPWR _11906_ sky130_fd_sc_hd__o311a_1
X_24850_ _04200_ _04201_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__xnor2_1
X_23801_ _03157_ _03158_ _03031_ _03026_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__a31o_1
X_24781_ _03549_ _04133_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__xnor2_1
X_21993_ _01549_ _01554_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23732_ net570 net574 top0.matmul0.matmul_stage_inst.f\[11\] VGND VGND VPWR VPWR
+ _03090_ sky130_fd_sc_hd__o21a_4
X_26520_ clknet_leaf_66_clk_sys _00143_ net660 VGND VGND VPWR VPWR top0.pid_q.out\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_20944_ _11758_ _12683_ VGND VGND VPWR VPWR _12792_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23663_ _03017_ net1017 VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__nor2_1
X_26451_ clknet_leaf_55_clk_sys _00092_ net668 VGND VGND VPWR VPWR top0.kiq\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20875_ _12238_ _12236_ VGND VGND VPWR VPWR _12724_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25402_ _04572_ _04745_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22614_ _02140_ _02167_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__xnor2_2
X_26382_ clknet_leaf_42_clk_sys _00023_ net684 VGND VGND VPWR VPWR top0.svm0.tC\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23594_ top0.matmul0.alpha_pass\[4\] _09272_ net559 VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25333_ _03829_ _04677_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22545_ net79 _02064_ _02067_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25264_ _04586_ _04590_ _04609_ _04406_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__o22a_1
XFILLER_0_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22476_ net80 _02031_ _02032_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__mux2_1
X_24215_ _03047_ _03195_ _03217_ _03572_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__o211a_1
X_27003_ clknet_leaf_28_clk_sys _00620_ net622 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21427_ net785 _12813_ _00993_ _12963_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__a22o_1
X_25195_ _04190_ _04288_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24146_ _02978_ _03252_ _03120_ _03355_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21358_ _13154_ _00925_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__nand2_1
X_20309_ _12103_ _12157_ VGND VGND VPWR VPWR _12158_ sky130_fd_sc_hd__xnor2_1
X_24077_ _03231_ _03269_ VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__xnor2_2
X_21289_ _13130_ _13131_ VGND VGND VPWR VPWR _13132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23028_ net168 top0.svm0.delta\[14\] VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__nor2_1
XFILLER_0_200_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15850_ _07839_ _07843_ _07945_ _07182_ _07845_ VGND VGND VPWR VPWR _07946_ sky130_fd_sc_hd__o221a_1
X_14801_ _06989_ _06990_ VGND VGND VPWR VPWR _07001_ sky130_fd_sc_hd__and2_1
X_15781_ net508 net481 _07877_ VGND VGND VPWR VPWR _07878_ sky130_fd_sc_hd__and3_1
X_24979_ _04329_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17520_ _09418_ _09421_ _09506_ VGND VGND VPWR VPWR _09507_ sky130_fd_sc_hd__o21ai_1
X_14732_ _06934_ VGND VGND VPWR VPWR _06935_ sky130_fd_sc_hd__buf_6
XFILLER_0_54_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26718_ clknet_leaf_82_clk_sys _00335_ net638 VGND VGND VPWR VPWR top0.pid_d.curr_int\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_99_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17451_ _09379_ _09384_ VGND VGND VPWR VPWR _09438_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14663_ _06268_ VGND VGND VPWR VPWR _06867_ sky130_fd_sc_hd__buf_6
X_26649_ clknet_leaf_75_clk_sys _00266_ net639 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16402_ _08393_ _08410_ _08489_ _08490_ VGND VGND VPWR VPWR _08491_ sky130_fd_sc_hd__a31o_1
X_13614_ _05815_ _05821_ _05826_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__a21o_1
X_17382_ net417 net340 VGND VGND VPWR VPWR _09369_ sky130_fd_sc_hd__nand2_1
X_14594_ net810 _06280_ _06799_ _06381_ VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19121_ net433 top0.pid_d.out_valid _11091_ VGND VGND VPWR VPWR _11092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16333_ net453 net510 VGND VGND VPWR VPWR _08423_ sky130_fd_sc_hd__nand2_1
X_13545_ _05500_ _05493_ _05494_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_65_clk_sys clknet_3_5__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_65_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_153_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_106_clk_sys clknet_3_0__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_106_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_19052_ _10999_ _11024_ VGND VGND VPWR VPWR _11025_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_164_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13476_ _05688_ _05493_ _05494_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__nor3_1
X_16264_ _08351_ _08354_ VGND VGND VPWR VPWR _08355_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18003_ net355 net370 VGND VGND VPWR VPWR _09988_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15215_ net525 net487 VGND VGND VPWR VPWR _07314_ sky130_fd_sc_hd__nand2_1
X_16195_ net504 VGND VGND VPWR VPWR _08287_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15146_ _07241_ _07244_ VGND VGND VPWR VPWR _07245_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19954_ _11410_ net185 VGND VGND VPWR VPWR _11824_ sky130_fd_sc_hd__nor2_1
X_15077_ _07161_ _07175_ VGND VGND VPWR VPWR _07176_ sky130_fd_sc_hd__xor2_1
X_14028_ _06124_ _06125_ _06119_ _06120_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__o22a_1
X_18905_ net320 _10877_ _10879_ VGND VGND VPWR VPWR _10880_ sky130_fd_sc_hd__a21o_1
X_19885_ _11730_ _11629_ VGND VGND VPWR VPWR _11760_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18836_ net308 _10697_ _10810_ _09688_ VGND VGND VPWR VPWR _10812_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18767_ _10655_ _10668_ _10666_ VGND VGND VPWR VPWR _10744_ sky130_fd_sc_hd__o21ai_1
X_15979_ _08072_ _08073_ VGND VGND VPWR VPWR _08074_ sky130_fd_sc_hd__or2b_1
X_17718_ _09699_ _09701_ _09704_ VGND VGND VPWR VPWR _09705_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18698_ _10608_ _10675_ VGND VGND VPWR VPWR _10676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17649_ net426 net319 VGND VGND VPWR VPWR _09636_ sky130_fd_sc_hd__nand2_2
XFILLER_0_77_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20660_ net294 _12505_ _12507_ _12508_ VGND VGND VPWR VPWR _12509_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19319_ _11254_ _11255_ _11258_ VGND VGND VPWR VPWR _11259_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20591_ _12435_ _12439_ VGND VGND VPWR VPWR _12440_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22330_ _01745_ _01867_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22261_ _01166_ net89 VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__nor2_2
X_24000_ _03305_ _03217_ _03060_ _03354_ _03357_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_143_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21212_ _12660_ _12575_ VGND VGND VPWR VPWR _13056_ sky130_fd_sc_hd__nand2_1
X_22192_ net127 _01144_ _01456_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__nor3_1
X_21143_ net257 net251 VGND VGND VPWR VPWR _12988_ sky130_fd_sc_hd__nand2_1
Xfanout501 net502 VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout512 net1029 VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__clkbuf_4
X_21074_ _12914_ _12919_ VGND VGND VPWR VPWR _12920_ sky130_fd_sc_hd__xor2_1
X_25951_ _12025_ _12010_ _12014_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__and3_1
Xfanout523 net524 VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout534 net535 VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout545 top0.pid_q.state\[4\] VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__clkbuf_4
Xfanout556 net557 VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__clkbuf_4
X_24902_ _03355_ _03765_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__xnor2_1
X_20025_ net201 net185 net195 VGND VGND VPWR VPWR _11890_ sky130_fd_sc_hd__o21a_1
Xfanout567 top0.matmul0.matmul_stage_inst.state\[4\] VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__clkbuf_4
X_25882_ _05088_ _05093_ top0.matmul0.beta_pass\[8\] VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__a21o_1
Xfanout578 net579 VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__clkbuf_4
Xfanout589 net606 VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__clkbuf_4
X_24833_ _04180_ _04184_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_38_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24764_ _04114_ _04115_ _04112_ _04113_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__o211ai_1
X_21976_ net156 net137 _01488_ _01486_ _01483_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__a311o_1
XFILLER_0_197_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26503_ clknet_leaf_82_clk_sys _00126_ net637 VGND VGND VPWR VPWR top0.pid_d.prev_int\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_23715_ _03056_ _03060_ _03065_ _03072_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__a22o_1
X_20927_ _12768_ _12774_ VGND VGND VPWR VPWR _12775_ sky130_fd_sc_hd__xnor2_2
X_24695_ _04032_ _04048_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26434_ clknet_leaf_98_clk_sys _00075_ net589 VGND VGND VPWR VPWR top0.kid\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23646_ net570 top0.matmul0.matmul_stage_inst.b\[5\] top0.matmul0.matmul_stage_inst.a\[5\]
+ net566 VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__a22o_4
X_20858_ net250 net259 VGND VGND VPWR VPWR _12707_ sky130_fd_sc_hd__or2b_1
XFILLER_0_7_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23577_ _02955_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26365_ _05414_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__clkbuf_1
X_20789_ _12622_ _12626_ _12628_ _12637_ VGND VGND VPWR VPWR _12638_ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13330_ _05542_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__buf_6
X_25316_ _04607_ _04656_ _04655_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__o21a_2
X_22528_ _02009_ _02044_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__nor2_2
X_26296_ net969 spi0.data_packed\[47\] net693 VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__mux2_1
X_13261_ _05467_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__buf_6
X_25247_ _04406_ _04590_ _04591_ _04593_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22459_ _01292_ _01770_ _02015_ net109 VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__a211o_1
X_15000_ _07041_ VGND VGND VPWR VPWR _07125_ sky130_fd_sc_hd__clkbuf_4
X_25178_ _04457_ _04458_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13192_ spi0.cs_sync\[2\] spi0.opcode\[6\] spi0.opcode\[7\] spi0.cs_sync\[1\] VGND
+ VGND VPWR VPWR _05423_ sky130_fd_sc_hd__and4b_1
XFILLER_0_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24129_ _03476_ _03456_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__xor2_2
XFILLER_0_130_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16951_ net550 _09007_ _09008_ VGND VGND VPWR VPWR _09009_ sky130_fd_sc_hd__and3_1
XFILLER_0_198_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15902_ _07987_ _07989_ VGND VGND VPWR VPWR _07997_ sky130_fd_sc_hd__or2_1
X_19670_ _11553_ _11554_ _11555_ _11556_ _11419_ net193 VGND VGND VPWR VPWR _11557_
+ sky130_fd_sc_hd__mux4_1
X_16882_ top0.matmul0.beta_pass\[4\] VGND VGND VPWR VPWR _08944_ sky130_fd_sc_hd__inv_2
X_18621_ _10596_ _10597_ VGND VGND VPWR VPWR _10599_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15833_ _07847_ _07859_ _07848_ VGND VGND VPWR VPWR _07929_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18552_ _10456_ _10483_ VGND VGND VPWR VPWR _10531_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15764_ _07847_ _07860_ VGND VGND VPWR VPWR _07861_ sky130_fd_sc_hd__xnor2_1
X_17503_ _09486_ _09489_ VGND VGND VPWR VPWR _09490_ sky130_fd_sc_hd__xnor2_1
X_14715_ _06916_ _06917_ VGND VGND VPWR VPWR _06918_ sky130_fd_sc_hd__xor2_1
X_18483_ _10461_ _10462_ VGND VGND VPWR VPWR _10463_ sky130_fd_sc_hd__and2b_1
X_15695_ _07716_ _07791_ VGND VGND VPWR VPWR _07793_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17434_ _09369_ _09419_ _09420_ VGND VGND VPWR VPWR _09421_ sky130_fd_sc_hd__a21bo_2
X_14646_ _06849_ _06850_ VGND VGND VPWR VPWR _06851_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17365_ net400 VGND VGND VPWR VPWR _09352_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_19 top0.svm0.out_valid VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14577_ _06775_ _06782_ VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19104_ _10996_ _11025_ _11075_ VGND VGND VPWR VPWR _11076_ sky130_fd_sc_hd__o21a_1
X_16316_ _08404_ _08326_ _08405_ VGND VGND VPWR VPWR _08406_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13528_ _05734_ _05740_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__xnor2_1
X_17296_ _09291_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19035_ _09966_ _10384_ _11005_ _11006_ _11007_ VGND VGND VPWR VPWR _11008_ sky130_fd_sc_hd__o41a_2
X_16247_ _08277_ _08279_ _08275_ VGND VGND VPWR VPWR _08338_ sky130_fd_sc_hd__a21bo_1
X_13459_ _05670_ _05671_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__nand2_2
XFILLER_0_88_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16178_ _08191_ _08196_ _08269_ VGND VGND VPWR VPWR _08270_ sky130_fd_sc_hd__o21a_1
X_15129_ net489 net484 VGND VGND VPWR VPWR _07228_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_10_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_195_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19937_ net201 _11510_ VGND VGND VPWR VPWR _11808_ sky130_fd_sc_hd__nor2_2
X_19868_ net241 _11721_ VGND VGND VPWR VPWR _11744_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18819_ net323 net327 VGND VGND VPWR VPWR _10795_ sky130_fd_sc_hd__or2b_1
X_19799_ _11679_ VGND VGND VPWR VPWR _11680_ sky130_fd_sc_hd__inv_2
X_21830_ net158 net153 VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_37_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21761_ _01321_ _01322_ _01266_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20712_ _12550_ _12557_ _12559_ _12560_ VGND VGND VPWR VPWR _12561_ sky130_fd_sc_hd__a211o_1
X_23500_ _05460_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_175_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24480_ _03694_ _03697_ _03695_ _03696_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21692_ _01165_ _01253_ _01250_ _01249_ _01160_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__o221ai_1
X_23431_ _02865_ _02867_ VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20643_ _12065_ _12491_ net298 VGND VGND VPWR VPWR _12492_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26150_ net18 _05292_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23362_ net120 _11783_ _02803_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__or3_1
X_20574_ _12251_ _12257_ _12340_ _12422_ VGND VGND VPWR VPWR _12423_ sky130_fd_sc_hd__or4_1
XFILLER_0_116_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25101_ _04363_ _04375_ _04361_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_117_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22313_ _01867_ _01872_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__xnor2_2
X_26081_ top0.matmul0.alpha_pass\[12\] _05237_ _05262_ VGND VGND VPWR VPWR _05263_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23293_ _02663_ _02665_ _02739_ _02664_ _11576_ net188 VGND VGND VPWR VPWR _02740_
+ sky130_fd_sc_hd__mux4_1
X_25032_ _04177_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__buf_4
XFILLER_0_131_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22244_ _01742_ _01803_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22175_ _01729_ _01732_ _01735_ _01736_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__or4_2
XFILLER_0_30_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21126_ _11788_ _12910_ _12969_ _12180_ _12970_ VGND VGND VPWR VPWR _12971_ sky130_fd_sc_hd__a221o_1
X_26983_ clknet_leaf_25_clk_sys _00600_ net628 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[15\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_13_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_13_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
Xfanout320 net1023 VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_5_clk_sys clknet_3_0__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_5_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout331 net332 VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkbuf_8
Xfanout342 top0.pid_d.mult0.b\[4\] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__buf_4
X_25934_ _05146_ _05147_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__xnor2_1
Xfanout353 net354 VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__clkbuf_2
X_21057_ _12844_ _12847_ _12902_ VGND VGND VPWR VPWR _12903_ sky130_fd_sc_hd__and3_1
Xfanout364 net367 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_4
Xfanout375 net376 VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__buf_2
Xfanout386 net387 VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkbuf_2
X_20008_ net201 _11411_ _11873_ net194 _11823_ VGND VGND VPWR VPWR _11874_ sky130_fd_sc_hd__o221a_1
Xfanout397 top0.pid_d.mult0.a\[7\] VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkbuf_2
X_25865_ _05083_ _05084_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__xor2_1
XFILLER_0_198_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24816_ _04125_ _04139_ _04167_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__o21a_1
X_25796_ _05025_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24747_ _02979_ _02980_ _03093_ _03094_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__o22a_1
XFILLER_0_68_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21959_ _01515_ _01520_ _01516_ net137 VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__o211a_1
XFILLER_0_179_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14500_ net33 _05605_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__nand2_2
XFILLER_0_56_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15480_ _07577_ _07578_ VGND VGND VPWR VPWR _07579_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24678_ _03993_ _04031_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_182_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14431_ _06583_ _06585_ VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__or2b_1
XFILLER_0_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26417_ clknet_leaf_59_clk_sys _00058_ net650 VGND VGND VPWR VPWR top0.kpq\[6\] sky130_fd_sc_hd__dfrtp_1
X_23629_ _02986_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17150_ _09163_ _09157_ _09164_ VGND VGND VPWR VPWR _09165_ sky130_fd_sc_hd__o21ai_2
X_14362_ _06569_ _06570_ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__xor2_1
X_26348_ spi0.data_packed\[72\] spi0.data_packed\[73\] net692 VGND VGND VPWR VPWR
+ _05406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16101_ net453 net1028 VGND VGND VPWR VPWR _08194_ sky130_fd_sc_hd__nand2_1
XFILLER_0_181_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13313_ _05522_ _05525_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__xor2_2
X_14293_ _06401_ _06406_ VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__or2_1
X_17081_ _00008_ _08855_ VGND VGND VPWR VPWR _09116_ sky130_fd_sc_hd__nor2_2
X_26279_ _05371_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16032_ net468 net507 VGND VGND VPWR VPWR _08126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13244_ top0.pid_d.state\[5\] net1019 VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17983_ _09964_ _09968_ VGND VGND VPWR VPWR _09969_ sky130_fd_sc_hd__xnor2_2
X_19722_ net1013 _11605_ _11593_ VGND VGND VPWR VPWR _11607_ sky130_fd_sc_hd__a21oi_1
X_16934_ _08990_ _08991_ VGND VGND VPWR VPWR _08993_ sky130_fd_sc_hd__or2_1
X_19653_ _11424_ _11528_ VGND VGND VPWR VPWR _11541_ sky130_fd_sc_hd__nor2_1
X_16865_ net546 _08920_ _08928_ net550 _08881_ VGND VGND VPWR VPWR _08929_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18604_ _10438_ _10582_ _10580_ VGND VGND VPWR VPWR _10583_ sky130_fd_sc_hd__a21o_1
X_15816_ _07813_ _07815_ VGND VGND VPWR VPWR _07912_ sky130_fd_sc_hd__nor2_1
X_19584_ _11469_ _11470_ _11471_ _11472_ VGND VGND VPWR VPWR _11473_ sky130_fd_sc_hd__or4_1
X_16796_ top0.pid_q.mult0.a\[7\] _08856_ _08859_ net775 _08871_ VGND VGND VPWR VPWR
+ _00156_ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18535_ _10512_ _10429_ _10513_ VGND VGND VPWR VPWR _10514_ sky130_fd_sc_hd__a21o_1
X_15747_ net541 net536 _07841_ _07843_ net448 VGND VGND VPWR VPWR _07844_ sky130_fd_sc_hd__o32a_1
XFILLER_0_88_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18466_ net392 _10203_ _09362_ VGND VGND VPWR VPWR _10446_ sky130_fd_sc_hd__o21ai_1
X_15678_ _07763_ _07774_ VGND VGND VPWR VPWR _07776_ sky130_fd_sc_hd__and2_1
X_17417_ net353 _09398_ _09400_ _09401_ _09403_ VGND VGND VPWR VPWR _09404_ sky130_fd_sc_hd__a221o_1
X_14629_ _06106_ _05629_ _05640_ net20 VGND VGND VPWR VPWR _06834_ sky130_fd_sc_hd__o211a_1
XFILLER_0_200_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18397_ _10371_ _10376_ VGND VGND VPWR VPWR _10378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17348_ _09329_ _09334_ _09335_ VGND VGND VPWR VPWR _09336_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17279_ top0.matmul0.matmul_stage_inst.mult1\[5\] top0.matmul0.matmul_stage_inst.mult2\[5\]
+ VGND VGND VPWR VPWR _09277_ sky130_fd_sc_hd__xor2_1
XFILLER_0_130_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19018_ _10982_ _10990_ _10903_ VGND VGND VPWR VPWR _10991_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20290_ net245 _12096_ _12138_ VGND VGND VPWR VPWR _12139_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23980_ _02989_ _02991_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__or2_1
XFILLER_0_199_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22931_ _02443_ _02444_ _02445_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25650_ top0.matmul0.sin\[4\] top0.matmul0.sin\[5\] _04914_ VGND VGND VPWR VPWR _04926_
+ sky130_fd_sc_hd__or3_2
X_22862_ top0.svm0.tB\[10\] VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24601_ _03842_ _03844_ _03955_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__o21ai_2
X_21813_ _01374_ _01350_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__xnor2_1
X_22793_ top0.svm0.counter\[15\] VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__inv_2
X_25581_ _05456_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24532_ _03883_ _03886_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__xnor2_2
X_21744_ net159 net141 VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27251_ clknet_3_2__leaf_clk_mosi _00865_ VGND VGND VPWR VPWR spi0.data_packed\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24463_ _03702_ _03733_ _03817_ _03700_ _03818_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__o221a_1
X_21675_ _01066_ _01113_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26202_ net3 spi0.data_packed\[0\] net694 VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__mux2_1
X_20626_ _12464_ _12471_ _12474_ VGND VGND VPWR VPWR _12475_ sky130_fd_sc_hd__o21a_1
X_23414_ _11439_ _02852_ net176 VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__o21ai_1
X_24394_ _03679_ _03750_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__nand2_2
X_27182_ clknet_leaf_88_clk_sys _00796_ net642 VGND VGND VPWR VPWR top0.periodTop_r\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26133_ spi0.data_packed\[28\] _05281_ _05282_ net922 VGND VGND VPWR VPWR _00809_
+ sky130_fd_sc_hd__a22o_1
X_23345_ _02771_ _02772_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__nand2_1
X_20557_ _12113_ _12114_ _12084_ _12404_ _12405_ VGND VGND VPWR VPWR _12406_ sky130_fd_sc_hd__o41a_1
XFILLER_0_104_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26064_ top0.pid_d.out\[8\] _05232_ _05233_ spi0.data_packed\[72\] VGND VGND VPWR
+ VPWR _05250_ sky130_fd_sc_hd__a22o_1
X_23276_ net150 _02723_ _02724_ _02722_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__a22o_1
X_20488_ net294 net280 VGND VGND VPWR VPWR _12337_ sky130_fd_sc_hd__nand2_2
XFILLER_0_104_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25015_ _03112_ _03900_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__nor2_1
X_22227_ _01777_ _01785_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__nand2_1
X_22158_ _01706_ _01719_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21109_ _12953_ _12954_ _12675_ VGND VGND VPWR VPWR _12955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26966_ clknet_leaf_30_clk_sys _00583_ net621 VGND VGND VPWR VPWR top0.matmul0.b\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14980_ _07112_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__clkbuf_1
X_22089_ _01618_ _01641_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__xnor2_1
Xfanout150 net151 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__buf_4
Xfanout161 top0.cordic0.vec\[1\]\[1\] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__buf_2
Xfanout172 net173 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_2
X_13931_ _05737_ _05738_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__or2b_1
X_25917_ _05128_ _05131_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__or2_1
Xfanout183 net184 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__buf_2
Xfanout194 net196 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__buf_2
X_26897_ clknet_leaf_107_clk_sys _00514_ net577 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_16650_ _08732_ _08734_ VGND VGND VPWR VPWR _08736_ sky130_fd_sc_hd__or2_1
X_13862_ _05950_ _05952_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__xnor2_1
X_25848_ _05031_ _05068_ _05069_ _05028_ net867 VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__a32o_1
XFILLER_0_69_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15601_ _07699_ VGND VGND VPWR VPWR _07700_ sky130_fd_sc_hd__clkbuf_4
X_16581_ _08660_ _08667_ VGND VGND VPWR VPWR _08668_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13793_ top0.periodTop_r\[2\] _05523_ _05524_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__and3_1
X_25779_ net205 _02282_ _12019_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__a21o_1
XFILLER_0_201_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18320_ _10299_ _10300_ VGND VGND VPWR VPWR _10302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15532_ _07572_ _07573_ _07569_ VGND VGND VPWR VPWR _07631_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_56_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18251_ _10224_ _10232_ VGND VGND VPWR VPWR _10234_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15463_ _07556_ _07561_ VGND VGND VPWR VPWR _07562_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17202_ _09209_ _09210_ VGND VGND VPWR VPWR _09211_ sky130_fd_sc_hd__nand2_1
X_14414_ net41 _05625_ _06620_ _06621_ VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__a31o_1
XFILLER_0_154_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18182_ _10064_ _10163_ _10164_ VGND VGND VPWR VPWR _10165_ sky130_fd_sc_hd__a21oi_2
X_15394_ net472 net478 VGND VGND VPWR VPWR _07493_ sky130_fd_sc_hd__or2b_2
XFILLER_0_182_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17133_ top0.pid_q.curr_int\[2\] top0.pid_q.prev_int\[2\] VGND VGND VPWR VPWR _09150_
+ sky130_fd_sc_hd__xnor2_1
X_14345_ _06553_ VGND VGND VPWR VPWR _06554_ sky130_fd_sc_hd__inv_1
XFILLER_0_135_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17064_ net1018 _09105_ VGND VGND VPWR VPWR _09106_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14276_ _06484_ _06485_ VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16015_ net461 net1029 VGND VGND VPWR VPWR _08109_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13227_ _05443_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17966_ _09851_ _09854_ VGND VGND VPWR VPWR _09952_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16917_ top0.pid_q.prev_error\[6\] _08975_ _08976_ VGND VGND VPWR VPWR _08977_ sky130_fd_sc_hd__a21oi_2
X_19705_ net1013 _11589_ _11571_ VGND VGND VPWR VPWR _11591_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17897_ _09767_ _09773_ _09770_ VGND VGND VPWR VPWR _09884_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16848_ _08911_ _08912_ net550 VGND VGND VPWR VPWR _08913_ sky130_fd_sc_hd__o21a_1
X_19636_ _11438_ _11523_ _11524_ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_195_Right_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19567_ top0.cordic0.slte0.opA\[2\] top0.cordic0.slte0.opB\[2\] VGND VGND VPWR VPWR
+ _11456_ sky130_fd_sc_hd__or2b_1
XFILLER_0_88_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16779_ top0.kiq\[0\] _08860_ _08861_ VGND VGND VPWR VPWR _08862_ sky130_fd_sc_hd__and3_1
XFILLER_0_137_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18518_ net310 _10355_ _10496_ _09401_ VGND VGND VPWR VPWR _10498_ sky130_fd_sc_hd__a211o_1
XFILLER_0_158_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19498_ top0.pid_d.curr_int\[14\] top0.pid_d.prev_int\[14\] VGND VGND VPWR VPWR _11390_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18449_ _10427_ _10339_ _10428_ VGND VGND VPWR VPWR _10429_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21460_ _01022_ _01024_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20411_ _12245_ _12248_ _12259_ VGND VGND VPWR VPWR _12260_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21391_ _12883_ _00926_ _00958_ VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_160_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23130_ _07117_ _02621_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20342_ _12163_ _12187_ _12188_ _12189_ _12190_ VGND VGND VPWR VPWR _12191_ sky130_fd_sc_hd__o311a_1
XFILLER_0_3_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23061_ _05541_ top0.svm0.counter\[5\] _02557_ _02561_ VGND VGND VPWR VPWR _02562_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20273_ net289 _12102_ VGND VGND VPWR VPWR _12122_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22012_ net142 _01269_ _01569_ _01572_ _01573_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__a32o_1
X_26820_ clknet_leaf_48_clk_sys _00437_ net676 VGND VGND VPWR VPWR top0.svm0.state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_26751_ clknet_leaf_94_clk_sys _00368_ net591 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_23963_ _03308_ _03311_ _03320_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_166_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25702_ top0.matmul0.sin\[1\] _04965_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__xnor2_1
X_22914_ _02313_ top0.svm0.tC\[15\] _02430_ _02431_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__a22o_1
X_26682_ clknet_leaf_62_clk_sys _00299_ net648 VGND VGND VPWR VPWR top0.pid_d.curr_error\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_23894_ _03063_ _03064_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__nor2_4
XFILLER_0_98_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_162_Right_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25633_ _04886_ _05456_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__nor2_1
X_22845_ _02326_ _02328_ _02329_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_155_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_184_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25564_ _04869_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__clkbuf_1
X_22776_ top0.svm0.counter\[5\] top0.svm0.counter\[6\] top0.svm0.counter\[8\] top0.svm0.rising
+ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24515_ _03195_ _03825_ _03808_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__and3_1
XFILLER_0_186_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21727_ _01286_ _01288_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__xor2_2
XFILLER_0_66_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25495_ _04833_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27234_ clknet_3_6__leaf_clk_mosi _00848_ VGND VGND VPWR VPWR spi0.data_packed\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_24446_ _03004_ _03005_ _03093_ _03094_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__o22a_1
X_21658_ _01215_ _01219_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_201_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27165_ clknet_leaf_11_clk_sys _00779_ net601 VGND VGND VPWR VPWR top0.a_in_matmul\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_20609_ _12446_ _12455_ _12457_ VGND VGND VPWR VPWR _12458_ sky130_fd_sc_hd__a21o_1
X_24377_ _03702_ _03733_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21589_ _01071_ _01139_ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_90_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14130_ _06304_ _06305_ _06340_ VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__and3_1
X_26116_ net886 _05279_ _05280_ net32 VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__a22o_1
X_23328_ net1016 _02772_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__nor2_1
X_27096_ clknet_leaf_17_clk_sys _00713_ net611 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.a\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14061_ _06257_ _06273_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__xor2_1
X_26047_ _05168_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__buf_2
X_23259_ _02692_ _02693_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__and2b_1
XFILLER_0_123_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17820_ _09788_ _09806_ VGND VGND VPWR VPWR _09807_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17751_ _09726_ _09737_ VGND VGND VPWR VPWR _09738_ sky130_fd_sc_hd__or2_1
Xhold6 net6 VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__dlygate4sd3_1
X_14963_ _07103_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__clkbuf_1
X_26949_ clknet_leaf_9_clk_sys _00566_ net596 VGND VGND VPWR VPWR top0.matmul0.a\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16702_ _08784_ _08786_ VGND VGND VPWR VPWR _08787_ sky130_fd_sc_hd__and2_1
X_13914_ _06118_ _06102_ _06103_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__nand3_1
X_17682_ _09608_ _09663_ _09664_ _09668_ VGND VGND VPWR VPWR _09669_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14894_ _07067_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19421_ net431 _10243_ _11322_ VGND VGND VPWR VPWR _11323_ sky130_fd_sc_hd__a21o_1
X_16633_ _08718_ _08647_ VGND VGND VPWR VPWR _08719_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13845_ _06031_ _06030_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19352_ net923 _11275_ _11281_ _11201_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__a22o_1
X_16564_ _08645_ _08649_ VGND VGND VPWR VPWR _08651_ sky130_fd_sc_hd__nand2_1
X_13776_ _05988_ _05981_ _05984_ _05968_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18303_ _10283_ _10284_ VGND VGND VPWR VPWR _10285_ sky130_fd_sc_hd__or2b_1
XFILLER_0_174_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15515_ _07596_ _07613_ VGND VGND VPWR VPWR _07614_ sky130_fd_sc_hd__xnor2_1
X_19283_ _11225_ _11216_ top0.pid_d.prev_error\[10\] VGND VGND VPWR VPWR _11226_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_167_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16495_ _08515_ _08517_ _08513_ VGND VGND VPWR VPWR _08583_ sky130_fd_sc_hd__a21bo_1
X_18234_ _10121_ _10123_ _10119_ VGND VGND VPWR VPWR _10217_ sky130_fd_sc_hd__a21bo_1
X_15446_ _07543_ _07544_ VGND VGND VPWR VPWR _07545_ sky130_fd_sc_hd__xor2_1
XFILLER_0_167_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18165_ _10131_ _10148_ VGND VGND VPWR VPWR _10149_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15377_ _07182_ _07233_ _07475_ VGND VGND VPWR VPWR _07476_ sky130_fd_sc_hd__or3b_1
XFILLER_0_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17116_ net549 _07698_ _09134_ _05442_ VGND VGND VPWR VPWR _09135_ sky130_fd_sc_hd__o211a_2
XFILLER_0_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14328_ _06450_ _06451_ _06537_ VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18096_ net416 net313 VGND VGND VPWR VPWR _10080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17047_ net1018 _09097_ VGND VGND VPWR VPWR _09098_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14259_ _06389_ _06390_ _06469_ VGND VGND VPWR VPWR _06470_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18998_ _10961_ _10971_ VGND VGND VPWR VPWR _10972_ sky130_fd_sc_hd__nand2_1
X_17949_ net361 net370 VGND VGND VPWR VPWR _09935_ sky130_fd_sc_hd__nand2_1
X_20960_ _12675_ _12736_ _12807_ VGND VGND VPWR VPWR _12808_ sky130_fd_sc_hd__o21a_2
XFILLER_0_139_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19619_ top0.cordic0.slte0.opA\[2\] _11505_ _11462_ _11506_ _11507_ VGND VGND VPWR
+ VPWR _11508_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_177_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20891_ _12035_ VGND VGND VPWR VPWR _12740_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22630_ _02125_ _02173_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__and2_1
XFILLER_0_192_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22561_ _02108_ _02115_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24300_ _03653_ _03655_ _03656_ _03301_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__a31o_2
X_21512_ net111 net94 VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__xnor2_4
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25280_ _04617_ _04625_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__xnor2_4
X_22492_ top0.cordic0.sin\[5\] _12004_ _12035_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24231_ _03586_ _03587_ _03588_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__mux2_1
X_21443_ _00979_ _00980_ _00975_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24162_ _03518_ _03519_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21374_ net241 net223 VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23113_ top0.svm0.delta\[4\] top0.svm0.delta\[5\] _02604_ VGND VGND VPWR VPWR _02609_
+ sky130_fd_sc_hd__or3_1
X_20325_ _12163_ VGND VGND VPWR VPWR _12174_ sky130_fd_sc_hd__inv_2
X_24093_ _03384_ _03402_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__or2b_1
X_23044_ net168 _02543_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__or2_1
X_20256_ _12098_ _12099_ _12104_ VGND VGND VPWR VPWR _12105_ sky130_fd_sc_hd__a21o_1
XFILLER_0_177_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20187_ _12035_ VGND VGND VPWR VPWR _12036_ sky130_fd_sc_hd__buf_6
XFILLER_0_110_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26803_ clknet_leaf_65_clk_sys _00420_ net657 VGND VGND VPWR VPWR top0.pid_q.prev_int\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_24995_ _04341_ _04343_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__and2_1
X_26734_ clknet_leaf_100_clk_sys _00351_ net587 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_23946_ _03207_ _03208_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__or2_1
XFILLER_0_192_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26665_ clknet_leaf_75_clk_sys _00282_ net637 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_23877_ _03006_ _03234_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__nor2_2
XFILLER_0_169_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13630_ _05834_ _05835_ _05837_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__a21o_1
X_25616_ net70 top0.matmul0.cos\[11\] VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22828_ _02347_ top0.svm0.tA\[2\] VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26596_ clknet_leaf_68_clk_sys _00219_ net659 VGND VGND VPWR VPWR top0.pid_q.curr_int\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13561_ _05530_ _05538_ _05539_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__nor3_1
X_25547_ _04860_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22759_ net977 _02292_ _02295_ top0.pid_q.curr_int\[3\] VGND VGND VPWR VPWR _00422_
+ sky130_fd_sc_hd__a22o_1
X_15300_ _07377_ _07397_ _07398_ VGND VGND VPWR VPWR _07399_ sky130_fd_sc_hd__a21o_1
XFILLER_0_183_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16280_ _08262_ _08264_ _08370_ VGND VGND VPWR VPWR _08371_ sky130_fd_sc_hd__a21oi_2
X_25478_ _04754_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__inv_2
X_13492_ net52 net49 _05585_ _05587_ _05540_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__a41o_1
XFILLER_0_152_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15231_ net481 _07327_ _07329_ VGND VGND VPWR VPWR _07330_ sky130_fd_sc_hd__a21oi_2
X_27217_ clknet_3_1__leaf_clk_mosi _00831_ VGND VGND VPWR VPWR spi0.data_packed\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_24429_ _03726_ _03727_ _03060_ _03123_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27148_ clknet_leaf_30_clk_sys _00762_ net619 VGND VGND VPWR VPWR top0.b_in_matmul\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_15162_ _07233_ _07260_ VGND VGND VPWR VPWR _07261_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14113_ _05683_ _05894_ _05567_ _06320_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__and4_1
XFILLER_0_120_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27079_ clknet_leaf_22_clk_sys _00696_ net607 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_19970_ _11837_ _11838_ VGND VGND VPWR VPWR _11839_ sky130_fd_sc_hd__nor2_1
X_15093_ _07177_ _07178_ _07179_ VGND VGND VPWR VPWR _07192_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14044_ _06255_ _06256_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__nand2_1
X_18921_ _10808_ _10895_ _10819_ VGND VGND VPWR VPWR _10896_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18852_ _10766_ _10827_ VGND VGND VPWR VPWR _10828_ sky130_fd_sc_hd__xnor2_4
Xclkbuf_leaf_61_clk_sys clknet_3_4__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_61_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_102_clk_sys clknet_3_0__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_102_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_17803_ _09652_ _09660_ _09655_ VGND VGND VPWR VPWR _09790_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18783_ top0.pid_d.out\[10\] _10755_ _10759_ VGND VGND VPWR VPWR _10760_ sky130_fd_sc_hd__mux2_1
X_15995_ _08000_ _08061_ _08010_ VGND VGND VPWR VPWR _08089_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_66_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17734_ net392 net353 VGND VGND VPWR VPWR _09721_ sky130_fd_sc_hd__nand2_1
X_14946_ _07094_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17665_ _09648_ _09651_ VGND VGND VPWR VPWR _09652_ sky130_fd_sc_hd__xnor2_2
X_14877_ _07058_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__clkbuf_1
X_16616_ net507 net445 VGND VGND VPWR VPWR _08702_ sky130_fd_sc_hd__nand2_1
X_19404_ top0.pid_d.prev_int\[2\] VGND VGND VPWR VPWR _11307_ sky130_fd_sc_hd__inv_2
X_13828_ _06024_ _06026_ _06035_ _06040_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__a31o_1
XFILLER_0_134_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17596_ _09567_ net359 net349 VGND VGND VPWR VPWR _09583_ sky130_fd_sc_hd__a21o_1
X_16547_ _08630_ _08633_ VGND VGND VPWR VPWR _08634_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19335_ _11272_ VGND VGND VPWR VPWR _11273_ sky130_fd_sc_hd__buf_2
X_13759_ _05932_ _05933_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__xor2_1
XFILLER_0_57_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19266_ net1024 _11190_ top0.matmul0.alpha_pass\[9\] VGND VGND VPWR VPWR _11211_
+ sky130_fd_sc_hd__o21ai_1
X_16478_ _08560_ _08565_ VGND VGND VPWR VPWR _08566_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_75_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_183_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18217_ _10183_ _10199_ VGND VGND VPWR VPWR _10200_ sky130_fd_sc_hd__xnor2_2
X_15429_ _07351_ _07352_ _07302_ VGND VGND VPWR VPWR _07528_ sky130_fd_sc_hd__a21o_1
XFILLER_0_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19197_ _11145_ _11146_ VGND VGND VPWR VPWR _11148_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18148_ _10009_ _10037_ _10007_ VGND VGND VPWR VPWR _10132_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_14_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold203 top0.pid_d.prev_error\[12\] VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold214 top0.pid_q.prev_int\[11\] VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18079_ _10059_ _10061_ _10062_ _10058_ VGND VGND VPWR VPWR _10064_ sky130_fd_sc_hd__a31o_1
Xhold225 spi0.data_packed\[44\] VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 top0.c_out_calc\[13\] VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold247 _05374_ VGND VGND VPWR VPWR net947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 spi0.data_packed\[33\] VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__dlygate4sd3_1
X_20110_ _11426_ _11775_ VGND VGND VPWR VPWR _11968_ sky130_fd_sc_hd__and2_1
Xhold269 spi0.data_packed\[46\] VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__dlygate4sd3_1
X_21090_ _12865_ _12873_ _12868_ VGND VGND VPWR VPWR _12936_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20041_ _11807_ _11904_ _11901_ VGND VGND VPWR VPWR _11905_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23800_ _03018_ _03019_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__or2_2
X_24780_ _03017_ _03185_ _04132_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__a21oi_1
X_21992_ _01552_ _01553_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__xor2_1
XFILLER_0_197_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23731_ net569 net556 top0.matmul0.matmul_stage_inst.b\[0\] VGND VGND VPWR VPWR _03089_
+ sky130_fd_sc_hd__o21a_2
X_20943_ _12790_ _12708_ _12706_ VGND VGND VPWR VPWR _12791_ sky130_fd_sc_hd__nor3b_1
X_26450_ clknet_leaf_55_clk_sys _00091_ net667 VGND VGND VPWR VPWR top0.kiq\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23662_ _03018_ _03019_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__nor2_1
X_20874_ _12720_ _12721_ _12686_ _12687_ VGND VGND VPWR VPWR _12723_ sky130_fd_sc_hd__o211ai_1
X_25401_ _04743_ _04744_ _04518_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22613_ _02165_ _02166_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__xnor2_1
X_26381_ clknet_leaf_42_clk_sys _00022_ net684 VGND VGND VPWR VPWR top0.svm0.tC\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23593_ _02963_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_93_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25332_ _03123_ _03200_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__xnor2_1
X_22544_ _02064_ _02067_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25263_ _04475_ _04608_ _04588_ _04586_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22475_ _01230_ _01967_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__nor2_1
X_27002_ clknet_leaf_27_clk_sys _00619_ net615 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24214_ _03337_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__buf_2
X_21426_ _00991_ _00992_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__xnor2_2
X_25194_ _03900_ _04097_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24145_ _03234_ _03195_ _03121_ _03502_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__o211a_1
X_21357_ _00917_ _00924_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20308_ net304 _12156_ _12107_ net280 VGND VGND VPWR VPWR _12157_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24076_ _03345_ _03428_ _03433_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21288_ net214 _13129_ VGND VGND VPWR VPWR _13131_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23027_ net168 top0.svm0.delta\[14\] _02297_ _02522_ _02527_ VGND VGND VPWR VPWR
+ _02529_ sky130_fd_sc_hd__o2111ai_1
X_20239_ _12087_ _12038_ _11653_ VGND VGND VPWR VPWR _12088_ sky130_fd_sc_hd__o21ai_1
X_14800_ net868 _06279_ _07000_ _05465_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__a22o_1
X_15780_ _07767_ VGND VGND VPWR VPWR _07877_ sky130_fd_sc_hd__inv_2
X_24978_ top0.matmul0.matmul_stage_inst.mult2\[7\] _04328_ _03642_ VGND VGND VPWR
+ VPWR _04329_ sky130_fd_sc_hd__mux2_1
X_14731_ _06919_ _06933_ VGND VGND VPWR VPWR _06934_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26717_ clknet_leaf_75_clk_sys _00334_ net636 VGND VGND VPWR VPWR top0.pid_d.curr_int\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23929_ _03276_ _03286_ VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_118_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17450_ _09353_ _09430_ _09435_ net355 _09436_ VGND VGND VPWR VPWR _09437_ sky130_fd_sc_hd__a221o_2
XFILLER_0_54_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14662_ _06820_ _06849_ _06850_ VGND VGND VPWR VPWR _06866_ sky130_fd_sc_hd__o21ai_1
X_26648_ clknet_leaf_75_clk_sys _00265_ net639 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16401_ _08474_ _08477_ VGND VGND VPWR VPWR _08490_ sky130_fd_sc_hd__nor2_1
X_13613_ _05590_ _05825_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__xnor2_2
X_17381_ _09350_ _09361_ _09367_ VGND VGND VPWR VPWR _09368_ sky130_fd_sc_hd__o21ai_2
X_14593_ _06796_ _06798_ VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_138_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26579_ clknet_leaf_50_clk_sys _00202_ net672 VGND VGND VPWR VPWR top0.pid_q.prev_error\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19120_ top0.pid_d.state\[3\] net438 _07136_ VGND VGND VPWR VPWR _11091_ sky130_fd_sc_hd__or3_1
X_16332_ net456 net507 VGND VGND VPWR VPWR _08422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13544_ net32 _05488_ _05490_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__and3_2
XFILLER_0_109_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19051_ _11014_ _11023_ VGND VGND VPWR VPWR _11024_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16263_ _08352_ _08353_ VGND VGND VPWR VPWR _08354_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13475_ net38 VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__inv_1
XFILLER_0_109_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18002_ net351 net372 VGND VGND VPWR VPWR _09987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15214_ net520 net493 VGND VGND VPWR VPWR _07313_ sky130_fd_sc_hd__nand2_2
X_16194_ _08049_ VGND VGND VPWR VPWR _08286_ sky130_fd_sc_hd__inv_2
X_15145_ _07243_ VGND VGND VPWR VPWR _07244_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19953_ net195 net183 VGND VGND VPWR VPWR _11823_ sky130_fd_sc_hd__nand2_1
X_15076_ _07166_ _07168_ _07174_ VGND VGND VPWR VPWR _07175_ sky130_fd_sc_hd__a21bo_1
X_14027_ _06124_ _06125_ _06119_ _06120_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__or4_1
X_18904_ net363 _10878_ VGND VGND VPWR VPWR _10879_ sky130_fd_sc_hd__nand2_1
X_19884_ _11758_ VGND VGND VPWR VPWR _11759_ sky130_fd_sc_hd__clkbuf_4
X_18835_ _10494_ _10810_ VGND VGND VPWR VPWR _10811_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18766_ _10731_ _10742_ VGND VGND VPWR VPWR _10743_ sky130_fd_sc_hd__xnor2_2
X_15978_ _08068_ _08071_ VGND VGND VPWR VPWR _08073_ sky130_fd_sc_hd__nand2_1
XFILLER_0_175_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17717_ _09481_ _09480_ _09703_ VGND VGND VPWR VPWR _09704_ sky130_fd_sc_hd__a21o_1
X_14929_ _07085_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__clkbuf_1
X_18697_ _10670_ _10674_ VGND VGND VPWR VPWR _10675_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17648_ _09619_ _09632_ _09634_ VGND VGND VPWR VPWR _09635_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17579_ _09555_ _09562_ _09556_ _09565_ VGND VGND VPWR VPWR _09566_ sky130_fd_sc_hd__a31o_1
XFILLER_0_175_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19318_ _11249_ _11256_ _11257_ VGND VGND VPWR VPWR _11258_ sky130_fd_sc_hd__o21ai_1
X_20590_ _12436_ _12438_ VGND VGND VPWR VPWR _12439_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19249_ _11194_ _11185_ top0.pid_d.prev_error\[7\] VGND VGND VPWR VPWR _11195_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_182_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22260_ net91 net87 VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__and2b_1
XFILLER_0_115_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21211_ _12515_ _12531_ _12532_ VGND VGND VPWR VPWR _13055_ sky130_fd_sc_hd__nand3_1
XFILLER_0_5_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22191_ net132 _01144_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_182_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21142_ _12982_ _12986_ VGND VGND VPWR VPWR _12987_ sky130_fd_sc_hd__xnor2_2
Xfanout502 top0.pid_q.mult0.a\[14\] VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__clkbuf_4
Xfanout513 top0.pid_q.mult0.a\[10\] VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__buf_2
XFILLER_0_1_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21073_ _12916_ _12918_ VGND VGND VPWR VPWR _12919_ sky130_fd_sc_hd__xnor2_2
X_25950_ net207 _05015_ _12016_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__o21ai_1
Xfanout524 top0.pid_q.mult0.a\[6\] VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__clkbuf_4
Xfanout535 net536 VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__clkbuf_4
X_24901_ _03011_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__buf_2
X_20024_ top0.cordic0.slte0.opA\[6\] _11888_ _11889_ VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__a21bo_1
Xfanout546 net547 VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__clkbuf_4
Xfanout557 net558 VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__clkbuf_4
X_25881_ top0.c_out_calc\[9\] _05029_ _05099_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__a21bo_1
Xfanout568 net569 VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__clkbuf_4
Xfanout579 net586 VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__clkbuf_4
X_24832_ _04181_ _04183_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__xor2_1
X_24763_ _04112_ _04113_ _04114_ _04115_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__a211o_1
XFILLER_0_197_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21975_ net130 _01488_ _01486_ _01483_ _01489_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_179_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26502_ clknet_leaf_81_clk_sys _00125_ net636 VGND VGND VPWR VPWR top0.pid_d.prev_int\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_23714_ _03066_ _03067_ _03069_ _03071_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__o22a_1
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20926_ _12771_ _12773_ VGND VGND VPWR VPWR _12774_ sky130_fd_sc_hd__xnor2_1
X_24694_ _04035_ _04047_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26433_ clknet_leaf_99_clk_sys _00074_ net631 VGND VGND VPWR VPWR top0.kid\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_193_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23645_ _02983_ _03002_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__xnor2_4
X_20857_ _12206_ _12705_ net246 VGND VGND VPWR VPWR _12706_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_1_clk_sys clknet_3_2__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_1_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26364_ spi0.opcode\[0\] spi0.opcode\[1\] net691 VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__mux2_1
X_23576_ net980 top0.matmul0.b\[11\] _02948_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__mux2_1
X_20788_ _12308_ _12629_ _12632_ _12636_ VGND VGND VPWR VPWR _12637_ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25315_ _04660_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22527_ _02080_ _02082_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26295_ net950 VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25246_ _04406_ _04592_ _04475_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__o21ai_1
X_13260_ net47 _05472_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__nand2_2
XFILLER_0_122_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22458_ _01292_ _01770_ _01287_ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_33_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21409_ _12832_ _12833_ net241 VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__mux2_1
X_25177_ _04475_ _04524_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__xnor2_2
X_13191_ top0.ready VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22389_ _12742_ _01946_ _01947_ _12812_ net712 VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__a32o_1
X_24128_ _03485_ _03484_ _03481_ _03480_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24059_ _03409_ _03410_ _03412_ _03415_ _03416_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__o221a_1
X_16950_ _09005_ _09006_ VGND VGND VPWR VPWR _09008_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15901_ _07995_ VGND VGND VPWR VPWR _07996_ sky130_fd_sc_hd__inv_2
X_16881_ net476 _08890_ _08943_ _08930_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__o211a_1
XFILLER_0_159_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18620_ _10596_ _10597_ VGND VGND VPWR VPWR _10598_ sky130_fd_sc_hd__nand2_1
X_15832_ _07919_ _07927_ VGND VGND VPWR VPWR _07928_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_21_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18551_ _10483_ _10458_ net341 VGND VGND VPWR VPWR _10530_ sky130_fd_sc_hd__o21a_1
X_15763_ _07848_ _07859_ VGND VGND VPWR VPWR _07860_ sky130_fd_sc_hd__xor2_1
X_14714_ net37 _06268_ VGND VGND VPWR VPWR _06917_ sky130_fd_sc_hd__nand2_1
X_17502_ _09487_ _09488_ VGND VGND VPWR VPWR _09489_ sky130_fd_sc_hd__xor2_1
X_18482_ _10455_ _10460_ VGND VGND VPWR VPWR _10462_ sky130_fd_sc_hd__nand2_1
X_15694_ _07716_ _07791_ VGND VGND VPWR VPWR _07792_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17433_ net413 net343 net347 net407 VGND VGND VPWR VPWR _09420_ sky130_fd_sc_hd__a22o_1
X_14645_ _06829_ _06848_ VGND VGND VPWR VPWR _06850_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_170_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17364_ net396 VGND VGND VPWR VPWR _09351_ sky130_fd_sc_hd__inv_2
X_14576_ _05579_ _06776_ _06212_ _06645_ _06781_ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__o32a_1
XFILLER_0_131_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16315_ _08404_ _08326_ top0.pid_q.out\[8\] VGND VGND VPWR VPWR _08405_ sky130_fd_sc_hd__o21ba_1
X_19103_ _10996_ _11025_ _10994_ VGND VGND VPWR VPWR _11075_ sky130_fd_sc_hd__a21o_1
X_13527_ _05736_ _05739_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__xnor2_2
X_17295_ top0.matmul0.beta_pass\[7\] _09290_ net563 VGND VGND VPWR VPWR _09291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19034_ _11005_ _11006_ net311 net370 VGND VGND VPWR VPWR _11007_ sky130_fd_sc_hd__a2bb2o_1
X_16246_ _08286_ _08295_ _08336_ net468 VGND VGND VPWR VPWR _08337_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_179_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13458_ net60 _05604_ _05613_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_149_Left_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16177_ _08191_ _08196_ _08189_ VGND VGND VPWR VPWR _08269_ sky130_fd_sc_hd__a21bo_1
X_13389_ _05599_ _05600_ net173 _05601_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__a211o_2
XFILLER_0_11_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15128_ net489 net484 VGND VGND VPWR VPWR _07227_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19936_ _11410_ net1016 VGND VGND VPWR VPWR _11807_ sky130_fd_sc_hd__nor2_2
X_15059_ _07156_ _07157_ VGND VGND VPWR VPWR _07158_ sky130_fd_sc_hd__xnor2_1
X_19867_ _11727_ _11733_ VGND VGND VPWR VPWR _11743_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18818_ net323 net368 VGND VGND VPWR VPWR _10794_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_158_Left_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19798_ _11676_ _11678_ VGND VGND VPWR VPWR _11679_ sky130_fd_sc_hd__xor2_1
XFILLER_0_179_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18749_ _10631_ _10646_ _10647_ VGND VGND VPWR VPWR _10726_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21760_ _01177_ _01269_ net162 VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20711_ _12552_ _12555_ _11571_ _11608_ VGND VGND VPWR VPWR _12560_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_187_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21691_ _01130_ _01162_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23430_ _11515_ _02866_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20642_ net285 net273 VGND VGND VPWR VPWR _12491_ sky130_fd_sc_hd__xor2_4
XFILLER_0_190_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20573_ net304 _12329_ _12249_ VGND VGND VPWR VPWR _12422_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23361_ _11650_ _02803_ net1020 VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_167_Left_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25100_ _04434_ _04448_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22312_ _01868_ _01871_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26080_ top0.pid_d.out\[12\] _05232_ _05233_ spi0.data_packed\[76\] VGND VGND VPWR
+ VPWR _05262_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23292_ _11788_ _11427_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25031_ _04347_ _04380_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_147_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22243_ _01742_ _01803_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22174_ _01247_ _01253_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21125_ _11759_ _12910_ _12911_ VGND VGND VPWR VPWR _12970_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_111_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26982_ clknet_leaf_25_clk_sys _00599_ net627 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[14\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout310 top0.pid_d.mult0.b\[14\] VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__buf_4
Xfanout321 net322 VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__buf_1
Xfanout332 top0.pid_d.mult0.b\[7\] VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__buf_4
X_25933_ top0.matmul0.alpha_pass\[14\] net428 VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__xor2_1
Xfanout343 net344 VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__buf_2
X_21056_ net262 _12208_ VGND VGND VPWR VPWR _12902_ sky130_fd_sc_hd__or2_1
Xfanout354 net355 VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__clkbuf_4
Xfanout365 net367 VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_4
Xfanout376 top0.pid_d.mult0.a\[12\] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__buf_4
X_20007_ net189 _11824_ VGND VGND VPWR VPWR _11873_ sky130_fd_sc_hd__nor2_1
XFILLER_0_185_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout387 net389 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__buf_2
X_25864_ net1024 top0.matmul0.beta_pass\[8\] VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__xor2_1
Xfanout398 top0.pid_d.mult0.a\[7\] VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_198_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24815_ _04125_ _04139_ _04128_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__a21o_1
X_25795_ _05023_ _05024_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__and2_1
XFILLER_0_201_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24746_ _02989_ _02991_ _03090_ _03091_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__o22a_1
X_21958_ net161 _01102_ _01356_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20909_ net271 _12095_ VGND VGND VPWR VPWR _12757_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_189_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24677_ _03995_ _04030_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_167_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21889_ _01428_ _01447_ _01450_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14430_ net23 net1015 _06637_ VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__nand3_2
XFILLER_0_166_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26416_ clknet_leaf_61_clk_sys _00057_ net650 VGND VGND VPWR VPWR top0.kpq\[5\] sky130_fd_sc_hd__dfrtp_1
X_23628_ net565 net557 top0.matmul0.matmul_stage_inst.e\[5\] VGND VGND VPWR VPWR _02986_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14361_ net36 _05639_ VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26347_ _05405_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__clkbuf_1
X_23559_ top0.b_in_matmul\[3\] top0.matmul0.b\[3\] _02937_ VGND VGND VPWR VPWR _02946_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16100_ net450 net521 VGND VGND VPWR VPWR _08193_ sky130_fd_sc_hd__nand2_1
X_13312_ net43 _05523_ _05524_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17080_ _09114_ VGND VGND VPWR VPWR _09115_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14292_ _06401_ _06406_ VGND VGND VPWR VPWR _06502_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26278_ net973 spi0.data_packed\[38\] net688 VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16031_ net474 net503 VGND VGND VPWR VPWR _08125_ sky130_fd_sc_hd__nand2_1
X_25229_ _04568_ _04575_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13243_ _05458_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_176_Right_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17982_ net424 net426 _09967_ VGND VGND VPWR VPWR _09968_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19721_ _11430_ _11605_ VGND VGND VPWR VPWR _11606_ sky130_fd_sc_hd__or2_1
XFILLER_0_202_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16933_ _08990_ _08991_ VGND VGND VPWR VPWR _08992_ sky130_fd_sc_hd__nand2_1
X_19652_ net84 _11539_ _11422_ VGND VGND VPWR VPWR _11540_ sky130_fd_sc_hd__mux2_2
XFILLER_0_189_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16864_ _08927_ VGND VGND VPWR VPWR _08928_ sky130_fd_sc_hd__inv_2
X_18603_ _10421_ _10433_ _10436_ VGND VGND VPWR VPWR _10582_ sky130_fd_sc_hd__a21o_1
X_15815_ _07813_ _07815_ VGND VGND VPWR VPWR _07911_ sky130_fd_sc_hd__nand2_1
X_19583_ top0.cordic0.slte0.opA\[15\] top0.cordic0.slte0.opB\[15\] VGND VGND VPWR
+ VPWR _11472_ sky130_fd_sc_hd__and2b_1
X_16795_ top0.kiq\[7\] _08863_ _08866_ VGND VGND VPWR VPWR _08871_ sky130_fd_sc_hd__and3_1
XFILLER_0_172_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_189_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18534_ _10512_ _10429_ top0.pid_d.out\[7\] VGND VGND VPWR VPWR _10513_ sky130_fd_sc_hd__o21ba_1
X_15746_ net443 _07842_ _07838_ VGND VGND VPWR VPWR _07843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18465_ _10352_ _10357_ _10444_ _10255_ VGND VGND VPWR VPWR _10445_ sky130_fd_sc_hd__a2bb2o_1
X_15677_ _07763_ _07774_ VGND VGND VPWR VPWR _07775_ sky130_fd_sc_hd__nor2_1
XFILLER_0_200_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14628_ net25 _06832_ VGND VGND VPWR VPWR _06833_ sky130_fd_sc_hd__nand2_2
XFILLER_0_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17416_ _09360_ _09402_ VGND VGND VPWR VPWR _09403_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18396_ _10371_ _10376_ VGND VGND VPWR VPWR _10377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17347_ top0.matmul0.matmul_stage_inst.mult1\[14\] top0.matmul0.matmul_stage_inst.mult2\[14\]
+ VGND VGND VPWR VPWR _09335_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14559_ _06707_ _06709_ _06708_ VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17278_ _09274_ _09270_ _09275_ VGND VGND VPWR VPWR _09276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19017_ _10983_ VGND VGND VPWR VPWR _10990_ sky130_fd_sc_hd__inv_2
X_16229_ net545 _08247_ _08248_ net548 _08320_ VGND VGND VPWR VPWR _08321_ sky130_fd_sc_hd__a32o_1
XFILLER_0_67_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19919_ net224 _11779_ _11780_ VGND VGND VPWR VPWR _11792_ sky130_fd_sc_hd__o21ba_1
X_22930_ top0.svm0.counter\[1\] top0.svm0.delta\[1\] net555 top0.svm0.counter\[0\]
+ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_155_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22861_ top0.svm0.calc_ready _02297_ _02380_ net704 _02309_ VGND VGND VPWR VPWR _00439_
+ sky130_fd_sc_hd__a32o_1
X_24600_ _03842_ _03844_ _03840_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_39_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21812_ _01367_ _01371_ _01373_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__a21oi_1
X_25580_ _04877_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22792_ net168 top0.svm0.tA\[14\] VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24531_ _03884_ _03885_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__xnor2_1
X_21743_ _01303_ _01304_ net164 VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27250_ clknet_3_2__leaf_clk_mosi _00864_ VGND VGND VPWR VPWR spi0.data_packed\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_24462_ _03206_ _03223_ _03694_ _03698_ _03699_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__a2111o_1
X_21674_ net99 _01113_ net77 VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__o21a_1
XFILLER_0_163_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26201_ top0.ready _05331_ _05332_ net207 VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23413_ _02849_ _02851_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20625_ _12464_ _12471_ _12473_ VGND VGND VPWR VPWR _12474_ sky130_fd_sc_hd__a21bo_1
X_27181_ clknet_leaf_88_clk_sys _00795_ net643 VGND VGND VPWR VPWR top0.periodTop_r\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_191_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24393_ _03735_ _03749_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26132_ spi0.data_packed\[27\] _05281_ _05282_ net935 VGND VGND VPWR VPWR _00808_
+ sky130_fd_sc_hd__a22o_1
X_23344_ _11560_ _02652_ _02787_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__a21o_2
XFILLER_0_190_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20556_ _12083_ _12070_ _12071_ _12171_ VGND VGND VPWR VPWR _12405_ sky130_fd_sc_hd__nand4_1
XFILLER_0_22_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26063_ _05249_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__clkbuf_1
X_23275_ net150 _11857_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__nor2_1
X_20487_ net304 net281 _12287_ VGND VGND VPWR VPWR _12336_ sky130_fd_sc_hd__or3_1
XFILLER_0_132_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25014_ _03325_ _03743_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__nor2_1
X_22226_ _01777_ _01785_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22157_ _01711_ _01718_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21108_ _12738_ VGND VGND VPWR VPWR _12954_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26965_ clknet_leaf_31_clk_sys _00582_ net621 VGND VGND VPWR VPWR top0.matmul0.b\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_22088_ _01557_ _01558_ _01649_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__a21oi_1
Xfanout140 top0.cordic0.vec\[1\]\[5\] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout151 top0.cordic0.vec\[1\]\[3\] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout162 net167 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_4
X_13930_ _06139_ _06142_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__xnor2_4
Xfanout173 top0.svm0.state\[2\] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_4
X_25916_ _05128_ _05131_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__nand2_1
X_21039_ _12883_ _12885_ VGND VGND VPWR VPWR _12886_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26896_ clknet_leaf_106_clk_sys _00513_ net577 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout184 net185 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_195_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout195 net196 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__buf_2
X_13861_ _05959_ _05990_ _06073_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__a21o_1
X_25847_ _05067_ _05065_ net12 VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__or3_1
XFILLER_0_199_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15600_ top0.pid_q.state\[0\] net546 _07698_ VGND VGND VPWR VPWR _07699_ sky130_fd_sc_hd__nor3_1
XFILLER_0_199_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16580_ _08662_ _08666_ VGND VGND VPWR VPWR _08667_ sky130_fd_sc_hd__xor2_1
XFILLER_0_201_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13792_ top0.periodTop_r\[1\] _05520_ _05521_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25778_ net207 net209 _05010_ VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15531_ _07621_ _07629_ VGND VGND VPWR VPWR _07630_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24729_ _03883_ _03884_ _03885_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18250_ _10224_ _10232_ VGND VGND VPWR VPWR _10233_ sky130_fd_sc_hd__and2_1
X_15462_ _07557_ _07560_ VGND VGND VPWR VPWR _07561_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_195_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17201_ top0.pid_q.curr_int\[10\] top0.pid_q.prev_int\[10\] VGND VGND VPWR VPWR _09210_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_194_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14413_ _06568_ _06570_ VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18181_ _10073_ _10162_ VGND VGND VPWR VPWR _10164_ sky130_fd_sc_hd__nor2_1
X_15393_ net475 net472 net542 VGND VGND VPWR VPWR _07492_ sky130_fd_sc_hd__and3b_1
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17132_ _09147_ _09148_ VGND VGND VPWR VPWR _09149_ sky130_fd_sc_hd__nand2_1
X_14344_ _06484_ _06485_ _06552_ VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_92_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17063_ _09002_ top0.pid_q.curr_error\[9\] _09096_ VGND VGND VPWR VPWR _09105_ sky130_fd_sc_hd__mux2_1
X_14275_ net55 _06135_ VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__and2_2
X_16014_ _08019_ _08024_ _08107_ VGND VGND VPWR VPWR _08108_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13226_ _05448_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17965_ _09866_ _09949_ _09950_ VGND VGND VPWR VPWR _09951_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19704_ _11526_ _11589_ VGND VGND VPWR VPWR _11590_ sky130_fd_sc_hd__or2_1
X_16916_ top0.pid_q.curr_error\[6\] _08963_ _08964_ VGND VGND VPWR VPWR _08976_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17896_ _09858_ _09882_ VGND VGND VPWR VPWR _09883_ sky130_fd_sc_hd__xnor2_2
X_19635_ net300 _11435_ _11522_ VGND VGND VPWR VPWR _11524_ sky130_fd_sc_hd__and3_1
X_16847_ _08908_ _08909_ _08910_ VGND VGND VPWR VPWR _08912_ sky130_fd_sc_hd__a21oi_1
X_19566_ top0.cordic0.slte0.opA\[5\] _11453_ _11454_ VGND VGND VPWR VPWR _11455_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16778_ _08854_ VGND VGND VPWR VPWR _08861_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18517_ _10494_ _10496_ VGND VGND VPWR VPWR _10497_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15729_ _07817_ _07825_ VGND VGND VPWR VPWR _07826_ sky130_fd_sc_hd__xnor2_2
X_19497_ top0.pid_d.curr_int\[13\] _11289_ _11341_ _10985_ _11389_ VGND VGND VPWR
+ VPWR _00339_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18448_ _10427_ _10339_ top0.pid_d.out\[6\] VGND VGND VPWR VPWR _10428_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_185_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_56_clk_sys clknet_3_6__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_56_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18379_ _10293_ _10295_ _10359_ VGND VGND VPWR VPWR _10360_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20410_ _12252_ _12258_ VGND VGND VPWR VPWR _12259_ sky130_fd_sc_hd__nor2_1
X_21390_ _00928_ _00957_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20341_ _12161_ VGND VGND VPWR VPWR _12190_ sky130_fd_sc_hd__inv_2
XFILLER_0_183_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23060_ net49 top0.svm0.counter\[6\] VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__xnor2_1
X_20272_ _12100_ _12119_ _12120_ VGND VGND VPWR VPWR _12121_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22011_ _01155_ _01338_ net153 VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26750_ clknet_leaf_92_clk_sys _00367_ net599 VGND VGND VPWR VPWR top0.cordic0.slte0.opA\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_23962_ _03316_ _03319_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__xnor2_4
X_25701_ net72 top0.matmul0.sin\[0\] VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__nand2_1
X_22913_ _02405_ top0.svm0.tC\[14\] VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26681_ clknet_leaf_63_clk_sys _00298_ net647 VGND VGND VPWR VPWR top0.pid_d.curr_error\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_169_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23893_ _03068_ _03070_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25632_ top0.matmul0.sin\[2\] _04910_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__xnor2_1
X_22844_ _02341_ _02348_ _02363_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__or3b_1
XFILLER_0_168_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25563_ top0.matmul0.a\[4\] top0.matmul0.matmul_stage_inst.e\[4\] _04867_ VGND VGND
+ VPWR VPWR _04869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22775_ _02298_ top0.svm0.counter\[1\] top0.svm0.counter\[2\] top0.svm0.counter\[3\]
+ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__or4_1
XFILLER_0_52_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24514_ _03252_ _03719_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__nor2_1
X_21726_ net113 _01287_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25494_ top0.matmul0.matmul_stage_inst.mult1\[3\] _03960_ _04829_ VGND VGND VPWR
+ VPWR _04833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27233_ clknet_3_6__leaf_clk_mosi _00847_ VGND VGND VPWR VPWR spi0.data_packed\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24445_ _03207_ _03208_ _03090_ _03091_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__o22a_1
X_21657_ net118 _01100_ _01216_ _01218_ _01072_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__a221o_2
XFILLER_0_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27164_ clknet_leaf_11_clk_sys _00778_ net602 VGND VGND VPWR VPWR top0.a_in_matmul\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_20608_ _12436_ _12438_ _12456_ VGND VGND VPWR VPWR _12457_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_35_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24376_ _03716_ _03732_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__xor2_2
X_21588_ net149 _01149_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26115_ net895 _05279_ _05280_ net35 VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23327_ _02741_ _02742_ _02753_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__nor3_1
X_27095_ clknet_leaf_22_clk_sys _00712_ net608 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.a\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_20539_ _12361_ _12387_ _12372_ VGND VGND VPWR VPWR _12388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_201_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14060_ _06266_ _06272_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__or2_1
X_26046_ _05236_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23258_ _02686_ _02695_ _02701_ _02705_ _02706_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__o221a_1
XFILLER_0_162_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22209_ _01166_ _01769_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__xnor2_4
X_23189_ _02646_ _06799_ _02649_ net776 VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14962_ spi0.data_packed\[23\] top0.kiq\[7\] _07097_ VGND VGND VPWR VPWR _07103_
+ sky130_fd_sc_hd__mux2_1
X_17750_ _09733_ _09736_ VGND VGND VPWR VPWR _09737_ sky130_fd_sc_hd__or2_1
Xhold7 _00441_ VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__dlygate4sd3_1
X_26948_ clknet_leaf_9_clk_sys _00565_ net595 VGND VGND VPWR VPWR top0.matmul0.a\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16701_ _08730_ _08728_ _08785_ VGND VGND VPWR VPWR _08786_ sky130_fd_sc_hd__o21a_1
X_13913_ _06102_ _06103_ _06118_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__a21o_1
X_17681_ _09665_ _09666_ _09667_ VGND VGND VPWR VPWR _09668_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14893_ spi0.data_packed\[54\] top0.kpq\[6\] _07064_ VGND VGND VPWR VPWR _07067_
+ sky130_fd_sc_hd__mux2_1
X_26879_ clknet_leaf_42_clk_sys _00496_ net685 VGND VGND VPWR VPWR top0.svm0.tB\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19420_ net442 _11320_ _11321_ net436 _11159_ VGND VGND VPWR VPWR _11322_ sky130_fd_sc_hd__a32o_1
XFILLER_0_159_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16632_ net461 net466 VGND VGND VPWR VPWR _08718_ sky130_fd_sc_hd__nand2_1
X_13844_ net58 _05683_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19351_ net927 _11275_ _11281_ _11192_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__a22o_1
X_16563_ _08645_ _08649_ VGND VGND VPWR VPWR _08650_ sky130_fd_sc_hd__nor2_1
X_13775_ _05969_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18302_ _10277_ _10282_ VGND VGND VPWR VPWR _10284_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15514_ _07220_ _07605_ _07609_ _07612_ VGND VGND VPWR VPWR _07613_ sky130_fd_sc_hd__a211o_1
XFILLER_0_155_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16494_ _08509_ _08580_ _08581_ VGND VGND VPWR VPWR _08582_ sky130_fd_sc_hd__a21oi_2
X_19282_ top0.pid_d.curr_error\[10\] VGND VGND VPWR VPWR _11225_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18233_ _10077_ _10085_ _10086_ VGND VGND VPWR VPWR _10216_ sky130_fd_sc_hd__o21ai_1
X_15445_ net518 net480 _07258_ VGND VGND VPWR VPWR _07544_ sky130_fd_sc_hd__and3_1
XFILLER_0_154_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18164_ _10133_ _10147_ VGND VGND VPWR VPWR _10148_ sky130_fd_sc_hd__xor2_1
X_15376_ net541 net484 _07473_ _07474_ VGND VGND VPWR VPWR _07475_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14327_ _06453_ _06457_ VGND VGND VPWR VPWR _06537_ sky130_fd_sc_hd__xnor2_1
X_17115_ net546 _08853_ VGND VGND VPWR VPWR _09134_ sky130_fd_sc_hd__nor2_2
XFILLER_0_151_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18095_ _09986_ _09988_ _10078_ VGND VGND VPWR VPWR _10079_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_150_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17046_ _08885_ top0.pid_q.curr_error\[0\] _09096_ VGND VGND VPWR VPWR _09097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14258_ _06393_ _06468_ VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13209_ _05434_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14189_ net44 _05639_ _06289_ _05625_ net48 VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__a32o_1
XFILLER_0_96_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18997_ _10963_ _10970_ VGND VGND VPWR VPWR _10971_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17948_ _09840_ _09932_ _09933_ VGND VGND VPWR VPWR _09934_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17879_ _09862_ _09865_ VGND VGND VPWR VPWR _09866_ sky130_fd_sc_hd__xnor2_2
X_19618_ top0.cordic0.slte0.opA\[1\] top0.cordic0.slte0.opA\[0\] _11456_ VGND VGND
+ VPWR VPWR _11507_ sky130_fd_sc_hd__or3b_1
XFILLER_0_36_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20890_ _12675_ _12738_ VGND VGND VPWR VPWR _12739_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_75_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19549_ _11437_ VGND VGND VPWR VPWR _11438_ sky130_fd_sc_hd__buf_4
XFILLER_0_165_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22560_ _02111_ _02114_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__xor2_1
XFILLER_0_158_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21511_ net118 _01069_ _01070_ _01071_ _01072_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__a221o_2
XFILLER_0_63_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22491_ _01877_ _02003_ _02046_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__or3_1
XFILLER_0_185_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24230_ _03559_ _03568_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__xor2_2
XFILLER_0_145_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21442_ _00973_ _01007_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__xor2_2
XFILLER_0_44_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24161_ _03471_ _03517_ _03487_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21373_ _12761_ _12981_ net248 VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__mux2_1
X_23112_ _07117_ _02608_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__nor2_1
X_20324_ _12170_ _12171_ VGND VGND VPWR VPWR _12173_ sky130_fd_sc_hd__and2_1
X_24092_ _03423_ _03449_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__and2_1
X_23043_ net168 _02543_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__nand2_1
X_20255_ _12103_ VGND VGND VPWR VPWR _12104_ sky130_fd_sc_hd__inv_2
X_20186_ net176 _11429_ VGND VGND VPWR VPWR _12035_ sky130_fd_sc_hd__nand2_2
XFILLER_0_122_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26802_ clknet_leaf_64_clk_sys _00419_ net658 VGND VGND VPWR VPWR top0.pid_q.prev_int\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_24994_ _04341_ _04343_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__nor2_1
XFILLER_0_192_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23945_ _03207_ _03208_ _02976_ _02977_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__o22a_1
X_26733_ clknet_leaf_100_clk_sys _00350_ net587 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_98_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26664_ clknet_leaf_63_clk_sys _00281_ net656 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_103_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23876_ _02984_ _02986_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__nor2_2
XFILLER_0_196_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25615_ net753 _04896_ _04887_ _04899_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__o22a_1
X_22827_ top0.svm0.counter\[2\] VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__inv_2
X_26595_ clknet_leaf_68_clk_sys _00218_ net662 VGND VGND VPWR VPWR top0.pid_q.curr_int\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13560_ net44 _05586_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__nand2_1
X_25546_ top0.matmul0.b\[12\] top0.matmul0.matmul_stage_inst.f\[12\] _04856_ VGND
+ VGND VPWR VPWR _04860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22758_ net995 _02292_ _02295_ top0.pid_q.curr_int\[2\] VGND VGND VPWR VPWR _00421_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21709_ net141 _01270_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25477_ _04807_ _04819_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__xnor2_2
X_13491_ net52 _05587_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22689_ _02208_ _02239_ _02223_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_109_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15230_ _07241_ _07233_ _07328_ _07243_ VGND VGND VPWR VPWR _07329_ sky130_fd_sc_hd__o211a_1
XFILLER_0_191_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24428_ _03726_ _03727_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__and2_1
X_27216_ clknet_3_1__leaf_clk_mosi _00830_ VGND VGND VPWR VPWR spi0.data_packed\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27147_ clknet_leaf_31_clk_sys _00761_ net619 VGND VGND VPWR VPWR top0.b_in_matmul\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_15161_ net517 _07259_ VGND VGND VPWR VPWR _07260_ sky130_fd_sc_hd__xnor2_1
X_24359_ _03714_ _03715_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_112_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14112_ net32 _05496_ _06323_ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__and3_1
X_27078_ clknet_leaf_110_clk_sys _00695_ net579 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15092_ _07187_ _07190_ VGND VGND VPWR VPWR _07191_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14043_ _06179_ _06254_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__nand2_2
X_18920_ _10818_ VGND VGND VPWR VPWR _10895_ sky130_fd_sc_hd__inv_2
X_26029_ top0.matmul0.alpha_pass\[0\] _05203_ _05222_ VGND VGND VPWR VPWR _05223_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18851_ _10825_ _10826_ VGND VGND VPWR VPWR _10827_ sky130_fd_sc_hd__nor2_2
XFILLER_0_158_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17802_ _09652_ _09660_ VGND VGND VPWR VPWR _09789_ sky130_fd_sc_hd__or2_1
X_18782_ top0.pid_d.curr_int\[10\] _10758_ VGND VGND VPWR VPWR _10759_ sky130_fd_sc_hd__xnor2_1
X_15994_ _08073_ _08087_ _08072_ VGND VGND VPWR VPWR _08088_ sky130_fd_sc_hd__a21o_1
X_17733_ _09459_ _09708_ net395 _09688_ VGND VGND VPWR VPWR _09720_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_121_Left_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14945_ spi0.data_packed\[47\] top0.kid\[15\] _07086_ VGND VGND VPWR VPWR _07094_
+ sky130_fd_sc_hd__mux2_1
X_17664_ _09649_ _09650_ VGND VGND VPWR VPWR _09651_ sky130_fd_sc_hd__xnor2_1
X_14876_ spi0.data_packed\[78\] top0.kpd\[14\] _07053_ VGND VGND VPWR VPWR _07058_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19403_ top0.pid_d.curr_int\[2\] _11290_ _11293_ _11306_ VGND VGND VPWR VPWR _00328_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16615_ net510 net444 VGND VGND VPWR VPWR _08701_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_15_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13827_ net68 _06025_ _06039_ _06029_ _06034_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__a311oi_1
X_17595_ net423 _09531_ _09552_ _09581_ VGND VGND VPWR VPWR _09582_ sky130_fd_sc_hd__o31a_1
XFILLER_0_187_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19334_ _00006_ _11095_ VGND VGND VPWR VPWR _11272_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16546_ _08631_ _08632_ VGND VGND VPWR VPWR _08633_ sky130_fd_sc_hd__xnor2_1
X_13758_ net54 _05495_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19265_ net1024 top0.matmul0.alpha_pass\[9\] _11190_ VGND VGND VPWR VPWR _11210_
+ sky130_fd_sc_hd__or3_1
X_16477_ _08561_ _08564_ VGND VGND VPWR VPWR _08565_ sky130_fd_sc_hd__xnor2_2
X_13689_ _05886_ _05899_ _05901_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_143_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18216_ _10197_ _10198_ VGND VGND VPWR VPWR _10199_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15428_ _07302_ _07350_ _07400_ _07518_ _07526_ VGND VGND VPWR VPWR _07527_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_130_Left_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19196_ _11145_ _11146_ VGND VGND VPWR VPWR _11147_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18147_ _10095_ _10130_ VGND VGND VPWR VPWR _10131_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_81_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15359_ net486 _07456_ _07457_ VGND VGND VPWR VPWR _07458_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_198_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold204 _00322_ VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 top0.cordic0.out_valid VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__dlygate4sd3_1
X_18078_ _10058_ _10059_ _10061_ _10062_ VGND VGND VPWR VPWR _10063_ sky130_fd_sc_hd__and4_1
Xhold226 _05378_ VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold237 top0.kpq\[15\] VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 top0.currT_r\[8\] VGND VGND VPWR VPWR net948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 top0.svm0.delta\[11\] VGND VGND VPWR VPWR net959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17029_ net428 VGND VGND VPWR VPWR _09081_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20040_ net202 _11902_ VGND VGND VPWR VPWR _11904_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21991_ _01069_ _01101_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23730_ net574 top0.matmul0.matmul_stage_inst.d\[0\] top0.matmul0.matmul_stage_inst.a\[0\]
+ net566 VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__a22o_2
X_20942_ net235 _12702_ _12703_ VGND VGND VPWR VPWR _12790_ sky130_fd_sc_hd__a21o_1
XFILLER_0_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23661_ net569 top0.matmul0.matmul_stage_inst.b\[10\] top0.matmul0.matmul_stage_inst.a\[10\]
+ net564 VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__a22o_2
X_20873_ _12686_ _12687_ _12720_ _12721_ VGND VGND VPWR VPWR _12722_ sky130_fd_sc_hd__a211o_1
X_25400_ _04561_ _04687_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__nand2_1
X_22612_ _01948_ _02067_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__or2_1
X_26380_ clknet_leaf_42_clk_sys _00021_ net684 VGND VGND VPWR VPWR top0.svm0.tC\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23592_ top0.matmul0.alpha_pass\[3\] _09267_ net559 VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25331_ _04097_ _04131_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22543_ _02026_ _02096_ _02097_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_10_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25262_ _04586_ _04592_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22474_ net79 _01166_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27001_ clknet_leaf_27_clk_sys _00618_ net615 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_24213_ _03185_ _03106_ _03323_ _03315_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21425_ _00958_ _00926_ _12883_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__o21a_1
X_25193_ _03200_ _04131_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24144_ _03501_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21356_ _00918_ _00923_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20307_ net289 net282 VGND VGND VPWR VPWR _12156_ sky130_fd_sc_hd__nand2b_2
X_24075_ _03345_ _03428_ _03349_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__a21bo_1
X_21287_ net213 _13129_ VGND VGND VPWR VPWR _13130_ sky130_fd_sc_hd__nand2_2
X_23026_ _02439_ _02526_ _02527_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__or3_1
X_20238_ net253 net249 VGND VGND VPWR VPWR _12087_ sky130_fd_sc_hd__and2_1
XFILLER_0_200_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20169_ top0.clarke_done top0.cordic0.out_valid _05437_ VGND VGND VPWR VPWR _12021_
+ sky130_fd_sc_hd__a21o_1
X_24977_ _04251_ _04327_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__xnor2_1
X_14730_ _06926_ _06932_ VGND VGND VPWR VPWR _06933_ sky130_fd_sc_hd__xor2_1
X_26716_ clknet_leaf_74_clk_sys _00333_ net638 VGND VGND VPWR VPWR top0.pid_d.curr_int\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_157_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23928_ _03284_ _03285_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14661_ _06852_ _06856_ _06864_ VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_200_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23859_ _03216_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__clkbuf_4
X_26647_ clknet_leaf_76_clk_sys _00264_ net639 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_197_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13612_ _05823_ _05824_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16400_ _08474_ _08477_ VGND VGND VPWR VPWR _08489_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14592_ _06697_ _06746_ _06797_ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17380_ _09350_ _09361_ _09366_ _09353_ VGND VGND VPWR VPWR _09367_ sky130_fd_sc_hd__a22o_1
X_26578_ clknet_leaf_50_clk_sys _00201_ net671 VGND VGND VPWR VPWR top0.pid_q.prev_error\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16331_ net449 net1029 VGND VGND VPWR VPWR _08421_ sky130_fd_sc_hd__nand2_1
X_13543_ net1030 _05484_ _05486_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__and3_2
XFILLER_0_109_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25529_ top0.matmul0.b\[4\] top0.matmul0.matmul_stage_inst.f\[4\] _04846_ VGND VGND
+ VPWR VPWR _04851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16262_ net521 net446 VGND VGND VPWR VPWR _08353_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19050_ _11016_ _11022_ VGND VGND VPWR VPWR _11023_ sky130_fd_sc_hd__xnor2_1
X_13474_ net35 _05488_ _05490_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18001_ net361 net366 VGND VGND VPWR VPWR _09986_ sky130_fd_sc_hd__nand2_2
X_15213_ _07310_ _07311_ VGND VGND VPWR VPWR _07312_ sky130_fd_sc_hd__xnor2_4
X_16193_ _08200_ _08211_ _08284_ VGND VGND VPWR VPWR _08285_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15144_ _07163_ _07164_ _07242_ VGND VGND VPWR VPWR _07243_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_65_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19952_ top0.cordic0.slte0.opA\[1\] _11802_ _11820_ _11821_ _11426_ VGND VGND VPWR
+ VPWR _11822_ sky130_fd_sc_hd__o221ai_4
X_15075_ _07166_ _07168_ _07173_ VGND VGND VPWR VPWR _07174_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_121_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14026_ _06204_ _06238_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__xnor2_4
X_18903_ net320 net324 net327 VGND VGND VPWR VPWR _10878_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19883_ _11757_ VGND VGND VPWR VPWR _11758_ sky130_fd_sc_hd__buf_4
X_18834_ net383 net379 _10495_ VGND VGND VPWR VPWR _10810_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18765_ _10732_ _10741_ VGND VGND VPWR VPWR _10742_ sky130_fd_sc_hd__xor2_1
XFILLER_0_175_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15977_ _08068_ _08071_ VGND VGND VPWR VPWR _08072_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17716_ _09481_ _09480_ _09490_ VGND VGND VPWR VPWR _09703_ sky130_fd_sc_hd__o21a_1
XFILLER_0_188_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14928_ spi0.data_packed\[39\] top0.kid\[7\] _07075_ VGND VGND VPWR VPWR _07085_
+ sky130_fd_sc_hd__mux2_1
X_18696_ _10671_ _10673_ VGND VGND VPWR VPWR _10674_ sky130_fd_sc_hd__xor2_1
X_17647_ _09619_ _09632_ _09633_ VGND VGND VPWR VPWR _09634_ sky130_fd_sc_hd__o21a_1
X_14859_ spi0.data_packed\[70\] top0.kpd\[6\] _07042_ VGND VGND VPWR VPWR _07049_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17578_ _09537_ _09564_ VGND VGND VPWR VPWR _09565_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19317_ top0.pid_d.prev_error\[13\] top0.pid_d.curr_error\[13\] VGND VGND VPWR VPWR
+ _11257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16529_ top0.pid_q.out\[11\] _07705_ _08616_ net544 VGND VGND VPWR VPWR _08617_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19248_ top0.pid_d.curr_error\[7\] VGND VGND VPWR VPWR _11194_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19179_ _09356_ _11125_ VGND VGND VPWR VPWR _11132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21210_ _12531_ _12532_ _12515_ VGND VGND VPWR VPWR _13054_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22190_ _01456_ _01749_ _01750_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_112_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21141_ _12984_ _12985_ VGND VGND VPWR VPWR _12986_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout503 net504 VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__clkbuf_4
X_21072_ _12785_ _12917_ VGND VGND VPWR VPWR _12918_ sky130_fd_sc_hd__xor2_1
Xfanout514 net515 VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout525 net526 VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__clkbuf_4
Xfanout536 top0.pid_q.mult0.a\[2\] VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__buf_2
X_24900_ _03863_ _04153_ _04246_ _04250_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__a31o_1
X_20023_ top0.cordic0.slte0.opA\[6\] _11784_ _11887_ VGND VGND VPWR VPWR _11889_ sky130_fd_sc_hd__or3_1
Xfanout547 top0.pid_q.state\[3\] VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__clkbuf_4
X_25880_ _05082_ _05092_ _05098_ _05439_ _12014_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__a221o_1
Xfanout558 net561 VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__clkbuf_4
Xfanout569 top0.matmul0.matmul_stage_inst.state\[2\] VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__clkbuf_4
X_24831_ _03006_ _04182_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__nor2_1
XFILLER_0_198_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24762_ _03996_ _03998_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__nor2_1
X_21974_ _01534_ _01535_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23713_ _03070_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__clkbuf_4
X_26501_ clknet_leaf_82_clk_sys net912 net636 VGND VGND VPWR VPWR top0.pid_d.prev_int\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20925_ net244 _12094_ _12772_ _12293_ _12138_ VGND VGND VPWR VPWR _12773_ sky130_fd_sc_hd__a221o_2
X_24693_ _04038_ _04046_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23644_ _02992_ _03001_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__xor2_2
X_26432_ clknet_leaf_77_clk_sys _00073_ net631 VGND VGND VPWR VPWR top0.kid\[5\] sky130_fd_sc_hd__dfrtp_1
X_20856_ net238 net234 VGND VGND VPWR VPWR _12705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_187_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26363_ _05413_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__clkbuf_1
X_23575_ _02954_ VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20787_ net299 net288 _12623_ _12635_ _11408_ VGND VGND VPWR VPWR _12636_ sky130_fd_sc_hd__o311a_1
XFILLER_0_147_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25314_ top0.matmul0.matmul_stage_inst.mult2\[12\] _04659_ _03146_ VGND VGND VPWR
+ VPWR _04660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22526_ _02081_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26294_ net949 spi0.data_packed\[46\] net693 VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25245_ _04517_ _04587_ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22457_ _01135_ _01292_ _02012_ _02013_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__a211o_1
XFILLER_0_84_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21408_ net248 _00971_ _00972_ _00974_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__a211o_1
X_25176_ _04515_ _04523_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__xnor2_1
X_13190_ top0.matmul0.matmul_stage_inst.state\[0\] _05421_ top0.matmul0.done_pass
+ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22388_ net210 _01885_ _01945_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__nand3_1
XFILLER_0_33_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24127_ _03468_ _03470_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21339_ _13179_ _13180_ VGND VGND VPWR VPWR _13181_ sky130_fd_sc_hd__and2b_1
X_24058_ _03401_ _03410_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__nand2_1
X_23009_ _02374_ _02297_ _02511_ _02513_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15900_ _07987_ _07989_ VGND VGND VPWR VPWR _07995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16880_ net546 _08935_ _08942_ net550 _08881_ VGND VGND VPWR VPWR _08943_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15831_ _07924_ _07926_ VGND VGND VPWR VPWR _07927_ sky130_fd_sc_hd__nand2_2
XFILLER_0_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18550_ _10523_ _10528_ VGND VGND VPWR VPWR _10529_ sky130_fd_sc_hd__xor2_1
X_15762_ _07853_ _07858_ VGND VGND VPWR VPWR _07859_ sky130_fd_sc_hd__xnor2_1
X_17501_ net329 net422 VGND VGND VPWR VPWR _09488_ sky130_fd_sc_hd__nand2_1
X_14713_ net36 _06824_ _06914_ _06915_ VGND VGND VPWR VPWR _06916_ sky130_fd_sc_hd__a31o_1
X_18481_ _10455_ _10460_ VGND VGND VPWR VPWR _10461_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15693_ _07778_ _07790_ VGND VGND VPWR VPWR _07791_ sky130_fd_sc_hd__xnor2_1
X_17432_ net413 net407 net343 net347 VGND VGND VPWR VPWR _09419_ sky130_fd_sc_hd__nand4_1
X_14644_ _06829_ _06848_ VGND VGND VPWR VPWR _06849_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14575_ _06780_ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__inv_2
X_17363_ _09344_ _09349_ VGND VGND VPWR VPWR _09350_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19102_ _11046_ _11073_ VGND VGND VPWR VPWR _11074_ sky130_fd_sc_hd__xnor2_4
X_16314_ top0.pid_q.curr_int\[8\] VGND VGND VPWR VPWR _08404_ sky130_fd_sc_hd__inv_2
X_13526_ _05737_ _05738_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17294_ _09288_ _09289_ VGND VGND VPWR VPWR _09290_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19033_ net371 net308 _11004_ VGND VGND VPWR VPWR _11006_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13457_ net60 _05604_ _05613_ _05624_ net64 VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__a32o_1
X_16245_ _08287_ net497 _08170_ _08335_ _08168_ VGND VGND VPWR VPWR _08336_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_126_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16176_ _08259_ _08267_ VGND VGND VPWR VPWR _08268_ sky130_fd_sc_hd__xnor2_4
X_13388_ top0.matmul0.done_pass top0.matmul0.state\[1\] VGND VGND VPWR VPWR _05601_
+ sky130_fd_sc_hd__nand2_4
X_15127_ _07225_ VGND VGND VPWR VPWR _07226_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19935_ _11510_ _11803_ _11805_ _11797_ VGND VGND VPWR VPWR _11806_ sky130_fd_sc_hd__o22a_1
X_15058_ net526 net475 VGND VGND VPWR VPWR _07157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_195_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14009_ _05504_ _05531_ _05532_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__or3_2
X_19866_ _11740_ _11741_ VGND VGND VPWR VPWR _11742_ sky130_fd_sc_hd__xnor2_2
X_18817_ net327 _10790_ VGND VGND VPWR VPWR _10793_ sky130_fd_sc_hd__and2_1
X_19797_ _11513_ _11677_ VGND VGND VPWR VPWR _11678_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18748_ _10716_ _10724_ VGND VGND VPWR VPWR _10725_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18679_ _10555_ _10557_ _10656_ VGND VGND VPWR VPWR _10657_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20710_ _12558_ VGND VGND VPWR VPWR _12559_ sky130_fd_sc_hd__buf_6
XFILLER_0_188_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21690_ _01249_ _01250_ _01251_ _01165_ _01160_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20641_ net280 _12287_ VGND VGND VPWR VPWR _12490_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23360_ _02799_ _02802_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20572_ _12340_ VGND VGND VPWR VPWR _12421_ sky130_fd_sc_hd__inv_2
XFILLER_0_190_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22311_ _01745_ _01870_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23291_ _02738_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25030_ _04377_ _04379_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__xor2_1
X_22242_ _01745_ _01802_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__xor2_2
X_22173_ _01247_ _01253_ _01734_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_112_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21124_ net227 _12910_ _12968_ VGND VGND VPWR VPWR _12969_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26981_ clknet_leaf_31_clk_sys _00598_ net619 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[13\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout300 net301 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__clkbuf_4
Xfanout311 net312 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_4
Xfanout322 top0.pid_d.mult0.b\[10\] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_4
X_25932_ top0.matmul0.alpha_pass\[13\] top0.matmul0.beta_pass\[13\] VGND VGND VPWR
+ VPWR _05146_ sky130_fd_sc_hd__nor2_2
X_21055_ _12039_ _12847_ VGND VGND VPWR VPWR _12901_ sky130_fd_sc_hd__nor2_1
Xfanout333 net335 VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__clkbuf_4
Xfanout344 net345 VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__clkbuf_4
Xfanout355 net356 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkbuf_4
Xfanout366 net367 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__clkbuf_2
X_20006_ top0.cordic0.slte0.opA\[5\] _11871_ _11872_ _11870_ VGND VGND VPWR VPWR _00365_
+ sky130_fd_sc_hd__a22o_1
Xfanout377 net379 VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__buf_2
X_25863_ top0.matmul0.alpha_pass\[7\] top0.matmul0.beta_pass\[7\] VGND VGND VPWR VPWR
+ _05083_ sky130_fd_sc_hd__nor2_2
Xfanout388 net389 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__clkbuf_4
Xfanout399 top0.pid_d.mult0.a\[7\] VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__clkbuf_2
X_24814_ _04161_ _04162_ _04164_ _04165_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__a211o_1
XFILLER_0_158_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25794_ _12024_ _05022_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24745_ _03496_ _04097_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__nor2_1
X_21957_ _01516_ _01518_ _01311_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20908_ _12715_ _12753_ _12755_ VGND VGND VPWR VPWR _12756_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24676_ _04028_ _04029_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21888_ _01448_ _01449_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23627_ _02984_ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__clkbuf_4
X_26415_ clknet_leaf_61_clk_sys _00056_ net650 VGND VGND VPWR VPWR top0.kpq\[4\] sky130_fd_sc_hd__dfrtp_1
X_20839_ net277 _12040_ _12212_ VGND VGND VPWR VPWR _12688_ sky130_fd_sc_hd__o21a_1
XFILLER_0_193_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14360_ net41 _05625_ VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__nand2_1
X_23558_ _02945_ VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__clkbuf_1
X_26346_ spi0.data_packed\[71\] spi0.data_packed\[72\] net689 VGND VGND VPWR VPWR
+ _05405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13311_ _05479_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__buf_2
XFILLER_0_108_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22509_ _01230_ _01775_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__nor2_1
X_14291_ _06492_ _06500_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__xnor2_4
X_26277_ net974 VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23489_ _02909_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16030_ net476 net502 VGND VGND VPWR VPWR _08124_ sky130_fd_sc_hd__nand2_1
X_13242_ _05457_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__clkbuf_4
X_25228_ _04570_ _04574_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25159_ _04436_ _04447_ _04434_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17981_ _09965_ _09966_ VGND VGND VPWR VPWR _09967_ sky130_fd_sc_hd__nor2_4
X_19720_ _11602_ _11604_ VGND VGND VPWR VPWR _11605_ sky130_fd_sc_hd__xnor2_1
X_16932_ top0.pid_q.prev_error\[8\] top0.pid_q.curr_error\[8\] VGND VGND VPWR VPWR
+ _08991_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19651_ _11535_ _11536_ _11537_ _11538_ _11419_ _11420_ VGND VGND VPWR VPWR _11539_
+ sky130_fd_sc_hd__mux4_1
X_16863_ _08925_ _08926_ VGND VGND VPWR VPWR _08927_ sky130_fd_sc_hd__xnor2_1
X_18602_ _10438_ _10580_ VGND VGND VPWR VPWR _10581_ sky130_fd_sc_hd__and2_1
XFILLER_0_172_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15814_ _07906_ _07909_ VGND VGND VPWR VPWR _07910_ sky130_fd_sc_hd__xnor2_4
X_19582_ top0.cordic0.slte0.opB\[15\] top0.cordic0.slte0.opA\[15\] VGND VGND VPWR
+ VPWR _11471_ sky130_fd_sc_hd__and2b_1
X_16794_ net524 _08856_ _08859_ net719 _08870_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18533_ top0.pid_d.curr_int\[7\] VGND VGND VPWR VPWR _10512_ sky130_fd_sc_hd__inv_2
X_15745_ _07182_ net443 VGND VGND VPWR VPWR _07842_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18464_ net390 _09518_ _09429_ _10074_ VGND VGND VPWR VPWR _10444_ sky130_fd_sc_hd__a22o_1
X_15676_ _07765_ _07773_ VGND VGND VPWR VPWR _07774_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17415_ net410 _09401_ net352 VGND VGND VPWR VPWR _09402_ sky130_fd_sc_hd__o21a_1
X_14627_ _05605_ VGND VGND VPWR VPWR _06832_ sky130_fd_sc_hd__buf_2
XFILLER_0_68_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18395_ _10372_ _10375_ VGND VGND VPWR VPWR _10376_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17346_ top0.matmul0.matmul_stage_inst.mult1\[14\] top0.matmul0.matmul_stage_inst.mult2\[14\]
+ VGND VGND VPWR VPWR _09334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14558_ _06760_ _06763_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13509_ top0.periodTop_r\[0\] _05721_ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__nand2_1
X_17277_ _09274_ _09270_ top0.matmul0.matmul_stage_inst.mult1\[4\] VGND VGND VPWR
+ VPWR _09275_ sky130_fd_sc_hd__o21ba_1
X_14489_ _06661_ _06662_ _06663_ _06695_ VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_3_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19016_ top0.pid_d.out\[13\] _09339_ _10989_ _10067_ VGND VGND VPWR VPWR _00258_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16228_ _08250_ _08319_ VGND VGND VPWR VPWR _08320_ sky130_fd_sc_hd__xor2_1
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16159_ _08227_ _08225_ _08228_ VGND VGND VPWR VPWR _08251_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19918_ net82 _11790_ VGND VGND VPWR VPWR _11791_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_52_clk_sys clknet_3_6__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_52_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_19849_ net234 VGND VGND VPWR VPWR _11726_ sky130_fd_sc_hd__inv_2
X_22860_ _02321_ _02359_ _02379_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_39_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21811_ net147 _01372_ _01332_ _01331_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22791_ top0.svm0.counter\[12\] top0.svm0.tA\[12\] VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__xor2_1
XFILLER_0_195_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24530_ _02989_ _02991_ _03061_ _03062_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21742_ net159 _01294_ _01093_ net157 VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__o22a_1
XFILLER_0_175_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24461_ _03206_ _03223_ _03694_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_171_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21673_ _01114_ _01233_ _01234_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__a21o_1
XFILLER_0_188_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23412_ _02838_ _02842_ _02850_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__a21o_1
X_26200_ net208 _12017_ top0.ready VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__o21a_1
X_20624_ net245 _12472_ VGND VGND VPWR VPWR _12473_ sky130_fd_sc_hd__xor2_1
X_27180_ clknet_leaf_88_clk_sys _00794_ net643 VGND VGND VPWR VPWR top0.periodTop_r\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_24392_ _03736_ _03748_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26131_ spi0.data_packed\[26\] _05281_ _05282_ top0.currT_r\[10\] VGND VGND VPWR
+ VPWR _00807_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23343_ net182 _02786_ _02668_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20555_ _12077_ _12082_ _12076_ VGND VGND VPWR VPWR _12404_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26062_ top0.a_in_matmul\[7\] _05248_ _05230_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23274_ net1014 _02722_ net176 VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20486_ _12333_ _12334_ net280 VGND VGND VPWR VPWR _12335_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25013_ _04278_ _04283_ _04362_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__o21a_1
X_22225_ _01784_ _01785_ net77 VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__o21a_1
X_22156_ _01714_ _01717_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_160_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21107_ _12736_ VGND VGND VPWR VPWR _12953_ sky130_fd_sc_hd__inv_2
X_26964_ clknet_leaf_31_clk_sys _00581_ net617 VGND VGND VPWR VPWR top0.matmul0.b\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout130 top0.cordic0.vec\[1\]\[6\] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_4
X_22087_ _01557_ _01558_ _01555_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_100_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout141 net143 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__buf_2
XFILLER_0_195_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout152 net154 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_4
X_25915_ _05129_ _05130_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21038_ _12807_ _12881_ _12884_ _12675_ VGND VGND VPWR VPWR _12885_ sky130_fd_sc_hd__a22o_1
Xfanout163 net167 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
Xfanout174 net175 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_4
X_26895_ clknet_leaf_106_clk_sys _00512_ net577 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout185 net186 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_191_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout196 top0.cordic0.gm0.iter\[1\] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13860_ _05959_ _05990_ _06071_ _06072_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__o22a_1
X_25846_ _05065_ _05066_ _05067_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_198_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22989_ top0.svm0.counter\[9\] _02495_ _02496_ _02494_ VGND VGND VPWR VPWR _00451_
+ sky130_fd_sc_hd__a22o_1
X_13791_ net68 _05517_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25777_ _02282_ _05009_ _05427_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__o21a_1
X_15530_ _07623_ _07628_ VGND VGND VPWR VPWR _07629_ sky130_fd_sc_hd__xnor2_1
X_24728_ _03980_ _04079_ _04080_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_96_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15461_ _07558_ _07559_ VGND VGND VPWR VPWR _07560_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24659_ _03106_ _03826_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17200_ _09207_ _09203_ _09208_ VGND VGND VPWR VPWR _09209_ sky130_fd_sc_hd__o21a_1
X_14412_ _06568_ _06570_ VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18180_ _10073_ _10162_ VGND VGND VPWR VPWR _10163_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15392_ net541 _07407_ VGND VGND VPWR VPWR _07491_ sky130_fd_sc_hd__nor2_1
X_17131_ top0.pid_q.curr_int\[1\] top0.pid_q.prev_int\[1\] top0.pid_q.prev_int\[0\]
+ top0.pid_q.curr_int\[0\] VGND VGND VPWR VPWR _09148_ sky130_fd_sc_hd__o211ai_2
X_14343_ _06484_ _06485_ _06482_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__a21o_1
X_26329_ _05396_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14274_ _06403_ _06404_ _06483_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__o21a_2
X_17062_ top0.pid_q.curr_error\[8\] _09100_ _09102_ _08987_ VGND VGND VPWR VPWR _00189_
+ sky130_fd_sc_hd__a22o_1
X_16013_ _08019_ _08024_ _08017_ VGND VGND VPWR VPWR _08107_ sky130_fd_sc_hd__a21bo_1
X_13225_ _05447_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__buf_2
XFILLER_0_111_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_186_Left_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17964_ _09869_ _09872_ VGND VGND VPWR VPWR _09950_ sky130_fd_sc_hd__nor2_1
X_19703_ _11585_ _11588_ VGND VGND VPWR VPWR _11589_ sky130_fd_sc_hd__xnor2_1
X_16915_ _08963_ _08964_ top0.pid_q.curr_error\[6\] VGND VGND VPWR VPWR _08975_ sky130_fd_sc_hd__a21o_1
X_17895_ _09880_ _09881_ VGND VGND VPWR VPWR _09882_ sky130_fd_sc_hd__and2b_1
X_19634_ net1014 _11522_ net174 VGND VGND VPWR VPWR _11523_ sky130_fd_sc_hd__o21ai_1
X_16846_ _08908_ _08909_ _08910_ VGND VGND VPWR VPWR _08911_ sky130_fd_sc_hd__and3_1
XFILLER_0_137_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19565_ top0.cordic0.slte0.opA\[5\] _11453_ top0.cordic0.slte0.opB\[5\] VGND VGND
+ VPWR VPWR _11454_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_177_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16777_ _05448_ VGND VGND VPWR VPWR _08860_ sky130_fd_sc_hd__buf_2
XFILLER_0_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13989_ _06200_ _06201_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_195_Left_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18516_ net401 net396 _10495_ VGND VGND VPWR VPWR _10496_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15728_ _07819_ _07824_ VGND VGND VPWR VPWR _07825_ sky130_fd_sc_hd__xnor2_1
X_19496_ _11252_ _11387_ _11388_ VGND VGND VPWR VPWR _11389_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18447_ top0.pid_d.curr_int\[6\] VGND VGND VPWR VPWR _10427_ sky130_fd_sc_hd__inv_2
XFILLER_0_185_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15659_ _07755_ _07756_ VGND VGND VPWR VPWR _07757_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18378_ _10293_ _10295_ _10291_ VGND VGND VPWR VPWR _10359_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17329_ _09318_ _09319_ VGND VGND VPWR VPWR _09320_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_160_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20340_ _12176_ _12178_ _12164_ VGND VGND VPWR VPWR _12189_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20271_ _12108_ _12100_ _12102_ _12118_ VGND VGND VPWR VPWR _12120_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_113_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22010_ _01570_ _01571_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23961_ _03317_ _03318_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__xnor2_2
X_25700_ _04890_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__clkbuf_4
X_22912_ _02405_ top0.svm0.tC\[14\] top0.svm0.tC\[13\] _02317_ _02429_ VGND VGND VPWR
+ VPWR _02430_ sky130_fd_sc_hd__a221o_1
X_23892_ _03054_ _03055_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__nor2_2
X_26680_ clknet_leaf_64_clk_sys _00297_ net656 VGND VGND VPWR VPWR top0.pid_d.curr_error\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_22843_ _02356_ _02355_ _02353_ _02349_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__a211o_1
X_25631_ net72 _04905_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__or2_1
XFILLER_0_196_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22774_ top0.svm0.counter\[0\] VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__inv_2
X_25562_ _04868_ VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27301_ clknet_3_1__leaf_clk_mosi _00915_ VGND VGND VPWR VPWR spi0.opcode\[7\] sky130_fd_sc_hd__dfxtp_1
X_24513_ _03864_ _03867_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__xnor2_4
X_21725_ net129 net1031 VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__nand2_2
XFILLER_0_66_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25493_ _04832_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27232_ clknet_3_4__leaf_clk_mosi _00846_ VGND VGND VPWR VPWR spi0.data_packed\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_24444_ _03114_ _03799_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__nor2_1
X_21656_ net126 _01217_ VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20607_ _12436_ _12438_ _12435_ VGND VGND VPWR VPWR _12456_ sky130_fd_sc_hd__a21o_1
X_24375_ _03730_ _03731_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__xor2_2
XFILLER_0_46_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27163_ clknet_leaf_10_clk_sys _00777_ net602 VGND VGND VPWR VPWR top0.a_in_matmul\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_21587_ _01147_ _01148_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23326_ net216 _11631_ _02770_ _11426_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__a22oi_4
X_26114_ net832 _05279_ _05280_ net38 VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__a22o_1
XFILLER_0_201_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20538_ _12280_ _12360_ _12361_ VGND VGND VPWR VPWR _12387_ sky130_fd_sc_hd__a21oi_1
X_27094_ clknet_leaf_22_clk_sys _00711_ net608 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.a\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_1__f_clk_sys clknet_0_clk_sys VGND VGND VPWR VPWR clknet_3_1__leaf_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_162_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23257_ net155 _02695_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__or2_1
X_26045_ top0.a_in_matmul\[3\] _05235_ _05230_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__mux2_1
X_20469_ _11739_ _12317_ VGND VGND VPWR VPWR _12318_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22208_ net100 net95 VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__nor2b_4
X_23188_ _02646_ _06748_ _02649_ net834 VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__a22o_1
X_22139_ _01076_ _01206_ _01699_ _01700_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_100_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14961_ _07102_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__clkbuf_1
X_26947_ clknet_leaf_13_clk_sys _00564_ net595 VGND VGND VPWR VPWR top0.matmul0.a\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold8 net5 VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__dlygate4sd3_1
X_16700_ _08730_ _08728_ _08664_ VGND VGND VPWR VPWR _08785_ sky130_fd_sc_hd__a21bo_1
X_13912_ _05772_ _05783_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__nor2_1
X_17680_ net326 net329 net424 net427 VGND VGND VPWR VPWR _09667_ sky130_fd_sc_hd__and4_1
X_26878_ clknet_leaf_42_clk_sys _00495_ net684 VGND VGND VPWR VPWR top0.svm0.tB\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_14892_ _07066_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16631_ _08643_ _08651_ _08650_ VGND VGND VPWR VPWR _08717_ sky130_fd_sc_hd__a21o_1
XFILLER_0_202_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25829_ top0.matmul0.alpha_pass\[3\] top0.matmul0.beta_pass\[3\] VGND VGND VPWR VPWR
+ _05053_ sky130_fd_sc_hd__nor2_1
X_13843_ _06054_ _06055_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__and2_1
XFILLER_0_187_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19350_ _11280_ VGND VGND VPWR VPWR _11281_ sky130_fd_sc_hd__clkbuf_2
X_16562_ _08647_ _08648_ VGND VGND VPWR VPWR _08649_ sky130_fd_sc_hd__xnor2_1
X_13774_ _05945_ _05986_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18301_ _10277_ _10282_ VGND VGND VPWR VPWR _10283_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15513_ _07610_ _07611_ _07298_ VGND VGND VPWR VPWR _07612_ sky130_fd_sc_hd__mux2_1
X_19281_ net322 _11117_ _11220_ _11224_ _08889_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__o221a_1
XFILLER_0_195_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16493_ _08509_ _08580_ _08507_ VGND VGND VPWR VPWR _08581_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_84_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18232_ _10209_ _10214_ VGND VGND VPWR VPWR _10215_ sky130_fd_sc_hd__xor2_4
XFILLER_0_26_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15444_ net511 _07535_ _07536_ _07538_ _07542_ VGND VGND VPWR VPWR _07543_ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18163_ _10135_ _10146_ VGND VGND VPWR VPWR _10147_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15375_ net537 net534 net493 net489 VGND VGND VPWR VPWR _07474_ sky130_fd_sc_hd__and4_1
XFILLER_0_142_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17114_ net758 _09114_ _09133_ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__a21o_1
X_14326_ _06535_ VGND VGND VPWR VPWR _06536_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_4_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18094_ _09986_ _09988_ _09987_ VGND VGND VPWR VPWR _10078_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17045_ net551 _08881_ VGND VGND VPWR VPWR _09096_ sky130_fd_sc_hd__or2_4
XFILLER_0_1_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14257_ _06464_ _06467_ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13208_ _05433_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__buf_6
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14188_ _05565_ _05731_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__nor2_1
X_18996_ _10968_ _10969_ VGND VGND VPWR VPWR _10970_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17947_ _09841_ _09842_ _09856_ VGND VGND VPWR VPWR _09933_ sky130_fd_sc_hd__and3_1
XFILLER_0_178_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17878_ _09863_ _09864_ VGND VGND VPWR VPWR _09865_ sky130_fd_sc_hd__xnor2_1
X_16829_ top0.pid_q.prev_error\[0\] top0.pid_q.curr_error\[0\] VGND VGND VPWR VPWR
+ _08895_ sky130_fd_sc_hd__nand2_1
X_19617_ top0.cordic0.slte0.opB\[3\] top0.cordic0.slte0.opA\[3\] VGND VGND VPWR VPWR
+ _11506_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19548_ net299 VGND VGND VPWR VPWR _11437_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19479_ top0.pid_d.curr_int\[11\] _11290_ _11293_ _11372_ _11373_ VGND VGND VPWR
+ VPWR _00337_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21510_ net124 net118 VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22490_ _01877_ _02003_ _02046_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21441_ net241 _01005_ _01006_ net223 VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24160_ _03471_ _03517_ _03487_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21372_ net231 _13171_ _00934_ _00935_ _00939_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__o221a_1
XFILLER_0_114_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23111_ top0.svm0.delta\[5\] _02607_ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__xnor2_1
X_20323_ _12084_ _12117_ _12170_ _12171_ VGND VGND VPWR VPWR _12172_ sky130_fd_sc_hd__o22a_1
X_24091_ _03432_ _03448_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23042_ net36 net34 net32 _02542_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__or4_2
X_20254_ _12100_ _12102_ VGND VGND VPWR VPWR _12103_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20185_ _12004_ VGND VGND VPWR VPWR _12034_ sky130_fd_sc_hd__buf_6
XFILLER_0_122_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26801_ clknet_leaf_6_clk_sys _00418_ net591 VGND VGND VPWR VPWR top0.cordic0.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_24993_ _04295_ _04297_ _04342_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__o21a_1
X_26732_ clknet_leaf_103_clk_sys _00349_ net576 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_23944_ _03234_ _03114_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__nor2_2
XFILLER_0_99_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26663_ clknet_leaf_63_clk_sys _00280_ net656 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_23875_ _03044_ _03232_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_169_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25614_ net71 top0.matmul0.cos\[10\] VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__and2_1
X_22826_ _02345_ top0.svm0.tA\[11\] VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__nor2_1
X_26594_ clknet_leaf_68_clk_sys _00217_ net662 VGND VGND VPWR VPWR top0.pid_q.curr_int\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_67_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25545_ _04859_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22757_ top0.pid_q.prev_int\[1\] _02292_ _02295_ top0.pid_q.curr_int\[1\] VGND VGND
+ VPWR VPWR _00420_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13490_ _05701_ _05473_ _05702_ VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__o21ai_2
X_21708_ _01268_ _01269_ net162 VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__mux2_1
X_25476_ _04717_ _04810_ _04813_ _04712_ _04818_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__o221a_1
X_22688_ _02172_ _02238_ _02231_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__a21o_1
X_27215_ clknet_3_1__leaf_clk_mosi _00829_ VGND VGND VPWR VPWR spi0.data_packed\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_24427_ _03716_ _03732_ _03782_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__a21o_1
X_21639_ _01103_ _01200_ _01108_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27146_ clknet_leaf_14_clk_sys _00760_ net617 VGND VGND VPWR VPWR top0.b_in_matmul\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_15160_ _07230_ _07226_ VGND VGND VPWR VPWR _07259_ sky130_fd_sc_hd__nor2_1
X_24358_ _03713_ _03707_ _03708_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14111_ _06217_ net22 VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__and2_2
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23309_ _02753_ _02754_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__xor2_2
X_15091_ _07188_ _07189_ VGND VGND VPWR VPWR _07190_ sky130_fd_sc_hd__xor2_1
XFILLER_0_105_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24289_ _03644_ _03645_ _03623_ _03631_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__o211ai_1
X_27077_ clknet_leaf_22_clk_sys _00694_ net607 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14042_ _06179_ _06254_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__or2_1
X_26028_ top0.pid_d.out\[0\] _05198_ _05199_ spi0.data_packed\[64\] VGND VGND VPWR
+ VPWR _05222_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18850_ _10822_ _10823_ _10821_ VGND VGND VPWR VPWR _10826_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_30_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17801_ _09780_ _09787_ VGND VGND VPWR VPWR _09788_ sky130_fd_sc_hd__xnor2_1
X_18781_ _10756_ _10596_ _10757_ VGND VGND VPWR VPWR _10758_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15993_ _07905_ _07997_ _07995_ VGND VGND VPWR VPWR _08087_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_98_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17732_ _09353_ _09351_ net392 _09363_ VGND VGND VPWR VPWR _09719_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_99_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_99_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_14944_ _07093_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_173_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_199_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17663_ net326 net420 VGND VGND VPWR VPWR _09650_ sky130_fd_sc_hd__nand2_1
X_14875_ _07057_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19402_ net431 _10065_ _11305_ net442 _11139_ VGND VGND VPWR VPWR _11306_ sky130_fd_sc_hd__a221o_1
X_16614_ _08630_ _08631_ _08699_ VGND VGND VPWR VPWR _08700_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13826_ net62 _05523_ _05524_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__and3_1
XFILLER_0_187_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17594_ _09531_ _09580_ VGND VGND VPWR VPWR _09581_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19333_ top0.matmul0.alpha_pass\[0\] _05443_ _11120_ VGND VGND VPWR VPWR _11271_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16545_ net447 net507 VGND VGND VPWR VPWR _08632_ sky130_fd_sc_hd__nand2_1
X_13757_ _05968_ _05969_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19264_ net439 _11207_ _11208_ VGND VGND VPWR VPWR _11209_ sky130_fd_sc_hd__and3_1
X_16476_ _08562_ _08563_ VGND VGND VPWR VPWR _08564_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13688_ _05865_ _05900_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18215_ _10185_ _10196_ VGND VGND VPWR VPWR _10198_ sky130_fd_sc_hd__and2_1
X_15427_ _07520_ _07399_ _07524_ _07525_ VGND VGND VPWR VPWR _07526_ sky130_fd_sc_hd__o211a_1
XFILLER_0_182_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19195_ top0.pid_d.prev_error\[3\] top0.pid_d.curr_error\[3\] VGND VGND VPWR VPWR
+ _11146_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18146_ _10128_ _10129_ VGND VGND VPWR VPWR _10130_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15358_ net534 net491 VGND VGND VPWR VPWR _07457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14309_ net33 _05588_ VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__nand2_2
Xhold205 top0.currT_r\[5\] VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18077_ _09972_ _09974_ VGND VGND VPWR VPWR _10062_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold216 top0.c_out_calc\[14\] VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ _07233_ _07387_ VGND VGND VPWR VPWR _07388_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold227 top0.pid_d.curr_error\[7\] VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold238 top0.pid_d.prev_int\[6\] VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ _05662_ top0.currT_r\[14\] _08899_ VGND VGND VPWR VPWR _09080_ sky130_fd_sc_hd__or3_1
Xhold249 spi0.data_packed\[45\] VGND VGND VPWR VPWR net949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18979_ _10848_ _10952_ VGND VGND VPWR VPWR _10953_ sky130_fd_sc_hd__xnor2_1
X_21990_ net124 _01312_ _01551_ _01105_ _01125_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__a221o_1
X_20941_ _12786_ _12787_ net225 VGND VGND VPWR VPWR _12789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23660_ net572 top0.matmul0.matmul_stage_inst.d\[10\] top0.matmul0.matmul_stage_inst.c\[10\]
+ net557 VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__a22o_2
X_20872_ _12718_ _12719_ _12695_ VGND VGND VPWR VPWR _12721_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22611_ _02143_ _02164_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__xnor2_2
X_23591_ _02962_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25330_ _04621_ _04622_ _04674_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__a21oi_1
X_22542_ _02095_ _02069_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25261_ _04534_ _04538_ _04602_ _04606_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__a31o_1
XFILLER_0_173_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22473_ _02017_ _02029_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__xnor2_2
X_27000_ clknet_leaf_27_clk_sys _00617_ net615 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.mult1\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24212_ _03559_ _03566_ _03569_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__o21a_1
X_21424_ _00964_ _00990_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__xnor2_2
X_25192_ _04534_ _04537_ _04538_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24143_ _02976_ _02977_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__or2_1
X_21355_ _13141_ _13146_ _13110_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20306_ _12062_ _12068_ _12063_ VGND VGND VPWR VPWR _12155_ sky130_fd_sc_hd__or3b_1
X_24074_ _03425_ _03427_ _03431_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__nor3_1
X_21286_ _12911_ _13128_ _12761_ net222 _12826_ VGND VGND VPWR VPWR _13129_ sky130_fd_sc_hd__a221o_1
XFILLER_0_188_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23025_ top0.svm0.counter\[15\] top0.svm0.delta\[15\] VGND VGND VPWR VPWR _02527_
+ sky130_fd_sc_hd__xnor2_1
X_20237_ net249 _12038_ _12085_ VGND VGND VPWR VPWR _12086_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_200_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20168_ net205 _05437_ _12019_ VGND VGND VPWR VPWR _12020_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24976_ _04325_ _04326_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__nand2_1
X_20099_ top0.cordic0.slte0.opA\[12\] _11949_ VGND VGND VPWR VPWR _11958_ sky130_fd_sc_hd__nor2_1
XFILLER_0_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26715_ clknet_leaf_74_clk_sys _00332_ net638 VGND VGND VPWR VPWR top0.pid_d.curr_int\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_23927_ _03282_ _03283_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14660_ _06852_ _06856_ _06854_ VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__a21bo_1
X_26646_ clknet_leaf_75_clk_sys _00263_ net637 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_23858_ _03076_ _03077_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13611_ net57 _05588_ _05822_ _05536_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__a211o_1
X_22809_ top0.svm0.tA\[7\] net170 VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__and2b_1
X_14591_ _06697_ _06746_ _06691_ VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__o21ba_1
X_26577_ clknet_leaf_50_clk_sys _00200_ net671 VGND VGND VPWR VPWR top0.pid_q.prev_error\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23789_ net567 net560 VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__or2_1
XFILLER_0_200_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16330_ _08416_ _08419_ VGND VGND VPWR VPWR _08420_ sky130_fd_sc_hd__xnor2_2
X_13542_ _05752_ _05753_ _05751_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__a21bo_1
X_25528_ _04850_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16261_ net447 net1028 VGND VGND VPWR VPWR _08352_ sky130_fd_sc_hd__nand2_1
X_25459_ _04742_ _04739_ _04771_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__and3_1
X_13473_ net32 _05683_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18000_ _09983_ _09984_ VGND VGND VPWR VPWR _09985_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15212_ _07169_ _07170_ VGND VGND VPWR VPWR _07311_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_180_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16192_ _08200_ _08211_ _08198_ VGND VGND VPWR VPWR _08284_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27129_ clknet_leaf_33_clk_sys _00743_ net664 VGND VGND VPWR VPWR top0.c_out_calc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_15143_ _07163_ _07164_ _07162_ VGND VGND VPWR VPWR _07242_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19951_ top0.cordic0.slte0.opA\[1\] _11802_ _11814_ net189 _11806_ VGND VGND VPWR
+ VPWR _11821_ sky130_fd_sc_hd__a221o_1
X_15074_ net539 net470 _07171_ _07172_ VGND VGND VPWR VPWR _07173_ sky130_fd_sc_hd__a31o_1
X_14025_ _06221_ _06237_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__xnor2_4
X_18902_ net323 net327 _10876_ VGND VGND VPWR VPWR _10877_ sky130_fd_sc_hd__a21o_1
X_19882_ net225 VGND VGND VPWR VPWR _11757_ sky130_fd_sc_hd__inv_2
X_18833_ _10688_ _10705_ _10704_ VGND VGND VPWR VPWR _10809_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18764_ _10733_ _10740_ VGND VGND VPWR VPWR _10741_ sky130_fd_sc_hd__xnor2_2
X_15976_ _07979_ _08069_ _08070_ VGND VGND VPWR VPWR _08071_ sky130_fd_sc_hd__a21oi_1
X_17715_ _09699_ _09701_ VGND VGND VPWR VPWR _09702_ sky130_fd_sc_hd__or2_1
X_14927_ _07084_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__clkbuf_1
X_18695_ _10566_ _10567_ _10672_ VGND VGND VPWR VPWR _10673_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17646_ _09486_ _09489_ VGND VGND VPWR VPWR _09633_ sky130_fd_sc_hd__or2b_1
XFILLER_0_72_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14858_ _07048_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13809_ _06017_ _06019_ _06021_ _06012_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__o2bb2a_1
X_17577_ _09539_ _09542_ VGND VGND VPWR VPWR _09564_ sky130_fd_sc_hd__xnor2_1
X_14789_ _06951_ _06967_ VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19316_ top0.pid_d.prev_error\[13\] top0.pid_d.curr_error\[13\] VGND VGND VPWR VPWR
+ _11256_ sky130_fd_sc_hd__nor2_1
X_16528_ top0.pid_q.out\[11\] _08611_ _08615_ VGND VGND VPWR VPWR _08616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19247_ net332 _11117_ _11189_ _11193_ _08889_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__o221a_1
X_16459_ _08543_ _08546_ VGND VGND VPWR VPWR _08548_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19178_ _11120_ _11130_ VGND VGND VPWR VPWR _11131_ sky130_fd_sc_hd__and2_1
XFILLER_0_182_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18129_ _10015_ _10020_ _10013_ VGND VGND VPWR VPWR _10113_ sky130_fd_sc_hd__o21ba_1
X_21140_ net262 net238 VGND VGND VPWR VPWR _12985_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21071_ net265 net244 VGND VGND VPWR VPWR _12917_ sky130_fd_sc_hd__xnor2_2
Xfanout504 net505 VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__clkbuf_2
Xfanout515 net516 VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__buf_2
XFILLER_0_10_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20022_ _11650_ _11887_ net1020 VGND VGND VPWR VPWR _11888_ sky130_fd_sc_hd__a21o_1
Xfanout526 net527 VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__buf_4
Xfanout537 net538 VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__clkbuf_4
Xfanout548 net549 VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__clkbuf_4
Xfanout559 net561 VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24830_ _03719_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_198_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24761_ _03996_ _03998_ _03997_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__a21oi_2
X_21973_ _01471_ _01472_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__xnor2_1
X_26500_ clknet_leaf_74_clk_sys _00123_ net637 VGND VGND VPWR VPWR top0.pid_d.prev_int\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23712_ net567 net558 top0.matmul0.matmul_stage_inst.e\[8\] VGND VGND VPWR VPWR _03070_
+ sky130_fd_sc_hd__o21a_1
X_20924_ net244 net254 VGND VGND VPWR VPWR _12772_ sky130_fd_sc_hd__or2b_1
XFILLER_0_83_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24692_ _03942_ _04045_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26431_ clknet_leaf_99_clk_sys _00072_ net631 VGND VGND VPWR VPWR top0.kid\[4\] sky130_fd_sc_hd__dfrtp_1
X_23643_ _02994_ _02996_ _02998_ _03000_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__o22a_1
X_20855_ net235 _12702_ _12703_ VGND VGND VPWR VPWR _12704_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26362_ spi0.data_packed\[79\] spi0.opcode\[0\] net690 VGND VGND VPWR VPWR _05413_
+ sky130_fd_sc_hd__mux2_1
X_23574_ top0.b_in_matmul\[10\] top0.matmul0.b\[10\] _02948_ VGND VGND VPWR VPWR _02954_
+ sky130_fd_sc_hd__mux2_1
X_20786_ _12611_ _12633_ _12634_ net285 VGND VGND VPWR VPWR _12635_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25313_ _04607_ _04658_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22525_ _02077_ _02079_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_47_clk_sys clknet_3_7__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_47_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_162_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26293_ net926 VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25244_ _04475_ _04588_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22456_ _01770_ _01065_ _01135_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__and3b_1
XFILLER_0_150_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21407_ net228 _00942_ _00973_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__and3_1
X_25175_ _04517_ _04522_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22387_ net210 _01885_ _01945_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24126_ _03468_ _03470_ _03483_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__o21ba_1
X_21338_ _13176_ _13178_ VGND VGND VPWR VPWR _13180_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24057_ _03413_ _03414_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_8_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21269_ _13027_ _13033_ _13111_ VGND VGND VPWR VPWR _13112_ sky130_fd_sc_hd__a21o_2
XFILLER_0_25_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23008_ _02374_ _02512_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__nor2_1
XFILLER_0_194_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15830_ _07925_ VGND VGND VPWR VPWR _07926_ sky130_fd_sc_hd__inv_2
XFILLER_0_189_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15761_ _07855_ _07857_ VGND VGND VPWR VPWR _07858_ sky130_fd_sc_hd__xnor2_1
X_24959_ _04226_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__inv_2
XFILLER_0_188_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17500_ net325 net427 VGND VGND VPWR VPWR _09487_ sky130_fd_sc_hd__nand2_1
X_14712_ _06889_ _06890_ VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__nor2_1
X_18480_ net364 _10459_ VGND VGND VPWR VPWR _10460_ sky130_fd_sc_hd__nand2_1
X_15692_ _07786_ _07789_ VGND VGND VPWR VPWR _07790_ sky130_fd_sc_hd__xor2_1
X_17431_ _09414_ _09417_ VGND VGND VPWR VPWR _09418_ sky130_fd_sc_hd__xnor2_4
X_14643_ _06831_ _06847_ VGND VGND VPWR VPWR _06848_ sky130_fd_sc_hd__xnor2_1
X_26629_ clknet_leaf_64_clk_sys _00246_ net656 VGND VGND VPWR VPWR top0.pid_d.out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_196_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17362_ _09345_ _09348_ VGND VGND VPWR VPWR _09349_ sky130_fd_sc_hd__xnor2_2
X_14574_ _06776_ _06777_ _06779_ net28 VGND VGND VPWR VPWR _06780_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_131_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19101_ _11050_ _11072_ VGND VGND VPWR VPWR _11073_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16313_ _05443_ VGND VGND VPWR VPWR _08403_ sky130_fd_sc_hd__clkbuf_2
X_13525_ _05541_ _05637_ _05638_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__or3_1
XFILLER_0_153_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17293_ top0.matmul0.matmul_stage_inst.mult1\[7\] top0.matmul0.matmul_stage_inst.mult2\[7\]
+ VGND VGND VPWR VPWR _09289_ sky130_fd_sc_hd__xor2_1
XFILLER_0_166_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19032_ net371 net308 _11004_ VGND VGND VPWR VPWR _11005_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16244_ net503 _08290_ _08170_ VGND VGND VPWR VPWR _08335_ sky130_fd_sc_hd__a21boi_1
X_13456_ _05667_ _05668_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16175_ _08261_ _08266_ VGND VGND VPWR VPWR _08267_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_51_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13387_ top0.svm0.state\[0\] net430 top0.svm0.state\[1\] VGND VGND VPWR VPWR _05600_
+ sky130_fd_sc_hd__nand3b_1
XFILLER_0_112_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15126_ _07145_ _07223_ _07224_ VGND VGND VPWR VPWR _07225_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_195_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19934_ _11632_ _11804_ VGND VGND VPWR VPWR _11805_ sky130_fd_sc_hd__nor2_1
X_15057_ net528 net471 VGND VGND VPWR VPWR _07156_ sky130_fd_sc_hd__nand2_1
X_14008_ _06209_ _06220_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_128_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19865_ _11728_ _11732_ _11514_ VGND VGND VPWR VPWR _11741_ sky130_fd_sc_hd__o21ai_1
X_18816_ net368 _10711_ _10791_ VGND VGND VPWR VPWR _10792_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19796_ _11662_ _11661_ VGND VGND VPWR VPWR _11677_ sky130_fd_sc_hd__nand2b_1
X_15959_ _07954_ _07956_ _07952_ VGND VGND VPWR VPWR _08054_ sky130_fd_sc_hd__a21bo_1
X_18747_ _10718_ _10723_ VGND VGND VPWR VPWR _10724_ sky130_fd_sc_hd__xnor2_1
X_18678_ _10555_ _10557_ _10536_ VGND VGND VPWR VPWR _10656_ sky130_fd_sc_hd__o21a_1
XFILLER_0_194_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17629_ net427 VGND VGND VPWR VPWR _09616_ sky130_fd_sc_hd__inv_2
X_20640_ _12460_ _12461_ _12488_ VGND VGND VPWR VPWR _12489_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_190_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20571_ _12385_ _12409_ _12415_ _12419_ VGND VGND VPWR VPWR _12420_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22310_ _01869_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__inv_2
X_23290_ _02736_ _02737_ _01102_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22241_ _01796_ _01801_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__xor2_2
XFILLER_0_103_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22172_ _01160_ _01733_ _01168_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_169_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21123_ _11788_ _12765_ VGND VGND VPWR VPWR _12968_ sky130_fd_sc_hd__or2_2
XFILLER_0_2_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26980_ clknet_leaf_25_clk_sys _00597_ net628 VGND VGND VPWR VPWR top0.matmul0.alpha_pass\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout301 top0.cordic0.vec\[0\]\[1\] VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__clkbuf_4
Xfanout312 net313 VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__buf_2
X_25931_ _05139_ _05143_ _05144_ _05138_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__o2bb2a_1
Xfanout323 net324 VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_4
X_21054_ net255 _12208_ VGND VGND VPWR VPWR _12900_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout334 net336 VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__buf_4
Xfanout345 net346 VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__clkbuf_4
Xfanout356 top0.pid_d.mult0.b\[1\] VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__buf_4
X_20005_ top0.cordic0.slte0.opA\[5\] _11785_ VGND VGND VPWR VPWR _11872_ sky130_fd_sc_hd__nor2_1
Xfanout367 top0.pid_d.mult0.a\[15\] VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__buf_2
X_25862_ _05081_ _05073_ _05074_ net11 _05601_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__a221o_2
Xfanout378 net379 VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__clkbuf_4
Xfanout389 top0.pid_d.mult0.a\[9\] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24813_ _04141_ _04159_ _04142_ _03942_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__o211a_1
X_25793_ _05439_ _05022_ top0.clarke_done VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__a21o_1
XFILLER_0_198_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24744_ _03799_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_190_Right_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21956_ _01442_ _01517_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20907_ _11608_ net265 _12095_ _12754_ VGND VGND VPWR VPWR _12755_ sky130_fd_sc_hd__o31a_1
XFILLER_0_167_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24675_ _04027_ _04011_ _04012_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__and3b_1
X_21887_ _01376_ _01389_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26414_ clknet_leaf_62_clk_sys _00055_ net650 VGND VGND VPWR VPWR top0.kpq\[3\] sky130_fd_sc_hd__dfrtp_1
X_23626_ net569 net572 top0.matmul0.matmul_stage_inst.f\[5\] VGND VGND VPWR VPWR _02984_
+ sky130_fd_sc_hd__o21a_1
X_20838_ _12678_ _12679_ _12685_ VGND VGND VPWR VPWR _12687_ sky130_fd_sc_hd__nand3_2
XFILLER_0_194_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26345_ _05404_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__clkbuf_1
X_23557_ top0.b_in_matmul\[2\] top0.matmul0.b\[2\] _02937_ VGND VGND VPWR VPWR _02945_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20769_ _12609_ _12610_ _12617_ VGND VGND VPWR VPWR _12618_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13310_ _05478_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__buf_2
XFILLER_0_92_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22508_ _02061_ _02063_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__xnor2_4
X_14290_ _06494_ _06499_ VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__xnor2_2
X_26276_ spi0.data_packed\[36\] net973 net688 VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__mux2_1
X_23488_ net1007 top0.matmul0.sin\[13\] _02904_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__mux2_1
X_25227_ _04572_ _04573_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_165_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13241_ _05456_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__inv_2
X_22439_ _12036_ _01996_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25158_ _04490_ _04505_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_202_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24109_ _03305_ _03120_ _03324_ _03461_ VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__a31o_1
X_17980_ net311 VGND VGND VPWR VPWR _09966_ sky130_fd_sc_hd__inv_2
X_25089_ _03112_ _04288_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__nor2_1
X_16931_ _08988_ _08977_ _08989_ VGND VGND VPWR VPWR _08990_ sky130_fd_sc_hd__a21o_1
X_16862_ top0.pid_q.prev_error\[3\] top0.pid_q.curr_error\[3\] VGND VGND VPWR VPWR
+ _08926_ sky130_fd_sc_hd__xnor2_1
X_19650_ net157 net150 net144 net140 net198 net191 VGND VGND VPWR VPWR _11538_ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15813_ _07907_ _07908_ VGND VGND VPWR VPWR _07909_ sky130_fd_sc_hd__xnor2_2
X_18601_ _10421_ _10433_ _10436_ VGND VGND VPWR VPWR _10580_ sky130_fd_sc_hd__and3_1
X_19581_ top0.cordic0.slte0.opA\[14\] top0.cordic0.slte0.opB\[14\] VGND VGND VPWR
+ VPWR _11470_ sky130_fd_sc_hd__and2b_1
X_16793_ top0.kiq\[6\] _08863_ _08866_ VGND VGND VPWR VPWR _08870_ sky130_fd_sc_hd__and3_1
X_18532_ _10511_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15744_ net443 _07838_ VGND VGND VPWR VPWR _07841_ sky130_fd_sc_hd__xor2_1
XFILLER_0_172_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18463_ _10416_ _10442_ VGND VGND VPWR VPWR _10443_ sky130_fd_sc_hd__and2_2
XFILLER_0_197_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15675_ _07767_ _07772_ VGND VGND VPWR VPWR _07773_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17414_ net407 VGND VGND VPWR VPWR _09401_ sky130_fd_sc_hd__inv_2
X_14626_ _06766_ _06771_ _06830_ VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18394_ _10373_ _10374_ VGND VGND VPWR VPWR _10375_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17345_ top0.matmul0.matmul_stage_inst.mult1\[15\] top0.matmul0.matmul_stage_inst.mult2\[15\]
+ VGND VGND VPWR VPWR _09333_ sky130_fd_sc_hd__xor2_1
X_14557_ _06761_ _06762_ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__xor2_1
XFILLER_0_126_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13508_ _05718_ _05720_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__nor2_4
XFILLER_0_99_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17276_ top0.matmul0.matmul_stage_inst.mult2\[4\] VGND VGND VPWR VPWR _09274_ sky130_fd_sc_hd__inv_2
X_14488_ _06661_ _06665_ _06662_ _06560_ VGND VGND VPWR VPWR _06695_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19015_ net435 _10985_ _10988_ net432 _07138_ VGND VGND VPWR VPWR _10989_ sky130_fd_sc_hd__a221o_1
XFILLER_0_153_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16227_ _08316_ _08318_ VGND VGND VPWR VPWR _08319_ sky130_fd_sc_hd__nand2_1
X_13439_ _05619_ _05628_ _05615_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16158_ _08231_ _08249_ VGND VGND VPWR VPWR _08250_ sky130_fd_sc_hd__nand2_1
X_15109_ _07204_ _07207_ VGND VGND VPWR VPWR _07208_ sky130_fd_sc_hd__xnor2_2
X_16089_ _08174_ _08181_ VGND VGND VPWR VPWR _08182_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_107_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19917_ _11761_ _11762_ _11777_ _11515_ VGND VGND VPWR VPWR _11790_ sky130_fd_sc_hd__o31a_1
X_19848_ _11725_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19779_ _11655_ _11560_ _11660_ VGND VGND VPWR VPWR _11661_ sky130_fd_sc_hd__a21oi_2
X_21810_ net155 net160 VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__nand2b_2
X_22790_ _02297_ _02304_ _06381_ VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__a21o_1
X_21741_ _01266_ _01177_ _01155_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__or3_1
XFILLER_0_148_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24460_ _03781_ _03815_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21672_ _01117_ _01120_ _01126_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__and3_1
XFILLER_0_148_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23411_ _02838_ _02842_ _01211_ VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__o21a_1
XFILLER_0_190_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20623_ net270 net258 VGND VGND VPWR VPWR _12472_ sky130_fd_sc_hd__nand2_1
X_24391_ _03738_ _03747_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26130_ spi0.data_packed\[25\] _05281_ _05282_ net952 VGND VGND VPWR VPWR _00806_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20554_ _12116_ _12171_ _12084_ VGND VGND VPWR VPWR _12403_ sky130_fd_sc_hd__or3b_1
X_23342_ net217 _11657_ _11658_ _02657_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26061_ top0.matmul0.alpha_pass\[7\] _05237_ _05247_ VGND VGND VPWR VPWR _05248_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20485_ net304 _12057_ VGND VGND VPWR VPWR _12334_ sky130_fd_sc_hd__nor2_1
X_23273_ _02720_ _02721_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25012_ _04278_ _04283_ _04276_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_15_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22224_ _01775_ _01776_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22155_ net90 _01716_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21106_ _12940_ _12951_ VGND VGND VPWR VPWR _12952_ sky130_fd_sc_hd__xor2_2
X_26963_ clknet_leaf_14_clk_sys _00580_ net617 VGND VGND VPWR VPWR top0.matmul0.b\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_22086_ _01647_ _01646_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout120 net121 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_4
Xfanout131 net134 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__buf_4
Xfanout142 net143 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__buf_2
X_25914_ top0.matmul0.alpha_pass\[11\] top0.matmul0.beta_pass\[11\] VGND VGND VPWR
+ VPWR _05130_ sky130_fd_sc_hd__nor2_1
X_21037_ _12736_ _12879_ _12881_ VGND VGND VPWR VPWR _12884_ sky130_fd_sc_hd__a21o_1
Xfanout153 net154 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_4
Xfanout164 net167 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__buf_2
X_26894_ clknet_leaf_106_clk_sys _00511_ net577 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_156_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout175 top0.cordic0.state\[0\] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_98_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout186 top0.cordic0.gm0.iter\[3\] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__buf_2
Xfanout197 net198 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_4
X_25845_ top0.matmul0.alpha_pass\[6\] top0.matmul0.beta_pass\[6\] VGND VGND VPWR VPWR
+ _05067_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13790_ _05999_ _06002_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__nand2_1
X_25776_ _12009_ net205 VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__or2_1
X_22988_ top0.svm0.counter\[9\] _02483_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24727_ _03983_ _03988_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21939_ _01102_ _01301_ _01136_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15460_ net493 net506 VGND VGND VPWR VPWR _07559_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24658_ _04009_ _04010_ _04007_ _04008_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14411_ _06615_ _06618_ VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__xnor2_4
X_23609_ _02971_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15391_ _07440_ _07441_ VGND VGND VPWR VPWR _07490_ sky130_fd_sc_hd__xor2_2
X_24589_ _03942_ _03943_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17130_ top0.pid_q.curr_int\[1\] top0.pid_q.prev_int\[1\] VGND VGND VPWR VPWR _09147_
+ sky130_fd_sc_hd__nand2_1
X_14342_ _06547_ _06550_ VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__nand2_4
XFILLER_0_181_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26328_ spi0.data_packed\[62\] spi0.data_packed\[63\] net696 VGND VGND VPWR VPWR
+ _05396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17061_ top0.pid_q.curr_error\[7\] _09100_ _09102_ _08974_ VGND VGND VPWR VPWR _00188_
+ sky130_fd_sc_hd__a22o_1
X_14273_ net1025 _06351_ _06403_ _06404_ VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26259_ _05361_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16012_ _08097_ _08105_ VGND VGND VPWR VPWR _08106_ sky130_fd_sc_hd__xnor2_1
X_13224_ net551 _05441_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17963_ _09869_ _09872_ VGND VGND VPWR VPWR _09949_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19702_ _11586_ _11587_ VGND VGND VPWR VPWR _11588_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16914_ _08971_ _08973_ VGND VGND VPWR VPWR _08974_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17894_ _09859_ _09879_ VGND VGND VPWR VPWR _09881_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19633_ _11452_ _11521_ VGND VGND VPWR VPWR _11522_ sky130_fd_sc_hd__xnor2_1
X_16845_ top0.pid_q.prev_error\[2\] top0.pid_q.curr_error\[2\] VGND VGND VPWR VPWR
+ _08910_ sky130_fd_sc_hd__xor2_1
XFILLER_0_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19564_ top0.cordic0.slte0.opB\[4\] top0.cordic0.slte0.opA\[4\] VGND VGND VPWR VPWR
+ _11453_ sky130_fd_sc_hd__and2b_1
X_16776_ _08858_ VGND VGND VPWR VPWR _08859_ sky130_fd_sc_hd__buf_2
X_13988_ _06143_ _06152_ _06153_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18515_ _09967_ VGND VGND VPWR VPWR _10495_ sky130_fd_sc_hd__buf_2
X_15727_ _07820_ _07823_ VGND VGND VPWR VPWR _07824_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_158_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19495_ _11289_ _11291_ VGND VGND VPWR VPWR _11388_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18446_ _10426_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__clkbuf_1
X_15658_ net451 net536 VGND VGND VPWR VPWR _07756_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14609_ _06800_ _06809_ VGND VGND VPWR VPWR _06814_ sky130_fd_sc_hd__nor2_1
XFILLER_0_173_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18377_ _10352_ _10357_ VGND VGND VPWR VPWR _10358_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15589_ _07677_ _07687_ VGND VGND VPWR VPWR _07688_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17328_ top0.matmul0.matmul_stage_inst.mult1\[12\] top0.matmul0.matmul_stage_inst.mult2\[12\]
+ VGND VGND VPWR VPWR _09319_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17259_ top0.matmul0.matmul_stage_inst.mult1\[2\] top0.matmul0.matmul_stage_inst.mult2\[2\]
+ VGND VGND VPWR VPWR _09260_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20270_ net289 _12102_ _12118_ VGND VGND VPWR VPWR _12119_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23960_ _02979_ _02980_ _03027_ _03028_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__o22a_1
X_22911_ _02317_ top0.svm0.tC\[13\] top0.svm0.tC\[12\] _02374_ _02428_ VGND VGND VPWR
+ VPWR _02429_ sky130_fd_sc_hd__o221a_1
XFILLER_0_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23891_ _03248_ _03120_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__nand2_1
X_25630_ net870 _04904_ _04907_ _04909_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__a22o_1
X_22842_ top0.svm0.counter\[4\] _02322_ _02330_ _02340_ _02333_ VGND VGND VPWR VPWR
+ _02362_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_78_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25561_ net987 top0.matmul0.matmul_stage_inst.e\[3\] _04867_ VGND VGND VPWR VPWR
+ _04868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22773_ _02296_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_151_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27300_ clknet_3_1__leaf_clk_mosi _00914_ VGND VGND VPWR VPWR spi0.opcode\[6\] sky130_fd_sc_hd__dfxtp_1
X_24512_ _03865_ _03866_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__xor2_2
XFILLER_0_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21724_ net122 net106 VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__nand2_2
X_25492_ top0.matmul0.matmul_stage_inst.mult1\[2\] _03855_ _04829_ VGND VGND VPWR
+ VPWR _04832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27231_ clknet_3_5__leaf_clk_mosi _00845_ VGND VGND VPWR VPWR spi0.data_packed\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24443_ _03103_ _03104_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21655_ net121 VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_47_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20606_ _12440_ _12445_ _12454_ VGND VGND VPWR VPWR _12455_ sky130_fd_sc_hd__a21o_1
X_27162_ clknet_leaf_10_clk_sys _00776_ net602 VGND VGND VPWR VPWR top0.a_in_matmul\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_191_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24374_ _03199_ _03205_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__nand2_1
X_21586_ net143 net164 VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__and2b_1
XFILLER_0_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26113_ net900 _05279_ _05280_ net40 VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__a22o_1
X_23325_ _11876_ _02712_ _02769_ _11612_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__a22o_1
X_27093_ clknet_leaf_17_clk_sys _00710_ net611 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.a\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_20537_ _12279_ _12266_ VGND VGND VPWR VPWR _12386_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26044_ top0.matmul0.alpha_pass\[3\] _05203_ _05234_ VGND VGND VPWR VPWR _05235_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20468_ net257 net248 VGND VGND VPWR VPWR _12317_ sky130_fd_sc_hd__nand2_1
X_23256_ _02702_ _02703_ _02704_ _02660_ VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__o31a_1
XFILLER_0_123_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22207_ _01412_ _01767_ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__xnor2_2
X_23187_ _02646_ _06682_ _02649_ net821 VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20399_ _12247_ VGND VGND VPWR VPWR _12248_ sky130_fd_sc_hd__inv_2
X_22138_ net138 _01076_ _01206_ _01458_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__o211a_1
X_14960_ spi0.data_packed\[22\] top0.kiq\[6\] _07097_ VGND VGND VPWR VPWR _07102_
+ sky130_fd_sc_hd__mux2_1
X_26946_ clknet_leaf_9_clk_sys _00563_ net595 VGND VGND VPWR VPWR top0.matmul0.a\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_22069_ _01563_ _01211_ _01564_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__mux2_1
Xhold9 _00440_ VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ _05772_ _05783_ _05770_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_199_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26877_ clknet_leaf_42_clk_sys _00494_ net684 VGND VGND VPWR VPWR top0.svm0.tB\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14891_ spi0.data_packed\[53\] top0.kpq\[5\] _07064_ VGND VGND VPWR VPWR _07066_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16630_ _08707_ _08715_ VGND VGND VPWR VPWR _08716_ sky130_fd_sc_hd__xnor2_1
X_25828_ _05050_ _05051_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__and2_1
X_13842_ net59 _05683_ _05894_ net62 VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__a22o_1
X_16561_ net458 _07213_ _08575_ VGND VGND VPWR VPWR _08648_ sky130_fd_sc_hd__a21oi_4
X_13773_ _05928_ _05943_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__xor2_1
X_25759_ net716 _04925_ _05000_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18300_ _10278_ _10281_ VGND VGND VPWR VPWR _10282_ sky130_fd_sc_hd__xnor2_1
X_15512_ _07255_ _07604_ VGND VGND VPWR VPWR _07611_ sky130_fd_sc_hd__nor2_1
X_19280_ _11121_ _11223_ _11123_ VGND VGND VPWR VPWR _11224_ sky130_fd_sc_hd__a21o_1
X_16492_ _08519_ VGND VGND VPWR VPWR _08580_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18231_ _10212_ _10213_ VGND VGND VPWR VPWR _10214_ sky130_fd_sc_hd__xnor2_4
X_15443_ net480 _07539_ _07541_ net514 VGND VGND VPWR VPWR _07542_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18162_ _10144_ _10145_ VGND VGND VPWR VPWR _10146_ sky130_fd_sc_hd__and2b_1
XFILLER_0_167_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15374_ net534 net493 net489 net537 VGND VGND VPWR VPWR _07473_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17113_ top0.pid_q.curr_error\[15\] _08860_ _09116_ VGND VGND VPWR VPWR _09133_ sky130_fd_sc_hd__and3_1
X_14325_ _06453_ _06533_ _06534_ VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18093_ _10075_ _10076_ VGND VGND VPWR VPWR _10077_ sky130_fd_sc_hd__xor2_2
XFILLER_0_20_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17044_ net443 _08861_ _09095_ _08930_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__o211a_1
X_14256_ _06349_ _06465_ _06466_ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13207_ top0.matmul0.done_pass top0.matmul0.state\[1\] VGND VGND VPWR VPWR _05433_
+ sky130_fd_sc_hd__and2_1
X_14187_ _06394_ _06397_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18995_ net383 _10494_ _10851_ VGND VGND VPWR VPWR _10969_ sky130_fd_sc_hd__or3b_2
XFILLER_0_178_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17946_ _09841_ _09842_ _09856_ VGND VGND VPWR VPWR _09932_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17877_ net355 net374 VGND VGND VPWR VPWR _09864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19616_ top0.cordic0.slte0.opB\[2\] VGND VGND VPWR VPWR _11505_ sky130_fd_sc_hd__inv_2
X_16828_ top0.currT_r\[1\] _08893_ VGND VGND VPWR VPWR _08894_ sky130_fd_sc_hd__xnor2_2
X_19547_ _11408_ _11432_ _11436_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16759_ top0.pid_q.out\[15\] _07704_ VGND VGND VPWR VPWR _08843_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19478_ _10831_ _11341_ VGND VGND VPWR VPWR _11373_ sky130_fd_sc_hd__and2_1
XFILLER_0_186_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18429_ _10400_ _10409_ VGND VGND VPWR VPWR _10410_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21440_ net236 net227 VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__or2_1
XFILLER_0_185_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21371_ _00936_ _00938_ net252 VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23110_ top0.svm0.delta\[4\] _02604_ _02595_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__o21a_1
X_20322_ _12077_ _12082_ _12076_ VGND VGND VPWR VPWR _12171_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24090_ _03434_ _03447_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__xor2_1
XFILLER_0_43_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23041_ net40 _02541_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__or2_1
X_20253_ net258 _12101_ VGND VGND VPWR VPWR _12102_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_101_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20184_ _12032_ _12026_ _12033_ net206 VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26800_ clknet_leaf_108_clk_sys _00417_ net606 VGND VGND VPWR VPWR top0.cordic0.gm0.iter\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_24992_ _04295_ _04297_ _04293_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__a21o_1
X_26731_ clknet_leaf_103_clk_sys _00348_ net576 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_23943_ _03299_ _03300_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__nor2_2
XFILLER_0_192_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26662_ clknet_leaf_75_clk_sys _00279_ net637 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_23874_ _03042_ _03052_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__xor2_2
X_25613_ net850 _04896_ _04891_ _04898_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__o22a_1
X_22825_ top0.svm0.counter\[11\] VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26593_ clknet_leaf_70_clk_sys _00216_ net662 VGND VGND VPWR VPWR top0.pid_q.curr_int\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25544_ top0.matmul0.b\[11\] top0.matmul0.matmul_stage_inst.f\[11\] _04856_ VGND
+ VGND VPWR VPWR _04859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22756_ net991 _02292_ _02295_ top0.pid_q.curr_int\[0\] VGND VGND VPWR VPWR _00419_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21707_ net152 net146 VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__xnor2_2
X_25475_ _04748_ _04817_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__nand2_1
XFILLER_0_192_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22687_ _02077_ _02135_ _02168_ _02170_ _02137_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__a221o_1
X_27214_ clknet_3_4__leaf_clk_mosi _00828_ VGND VGND VPWR VPWR spi0.data_packed\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_24426_ _03730_ _03731_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__nor2_1
X_21638_ net144 _01101_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27145_ clknet_leaf_31_clk_sys _00759_ net619 VGND VGND VPWR VPWR top0.b_in_matmul\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24357_ _03707_ _03708_ _03713_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__o21ai_1
X_21569_ net118 net114 VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__nand2_1
X_14110_ _05484_ _05486_ _06046_ _06320_ _06321_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__a41o_1
X_23308_ _02741_ _02742_ _11512_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__o21a_1
X_27076_ clknet_leaf_22_clk_sys _00693_ net607 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.c\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_15090_ net531 net464 VGND VGND VPWR VPWR _07189_ sky130_fd_sc_hd__nand2_1
X_24288_ _03299_ _03300_ _03624_ _03625_ _03630_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_160_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14041_ _06239_ _06253_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__xor2_2
XFILLER_0_127_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26027_ _05221_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__clkbuf_1
X_23239_ net272 net266 net260 net254 net198 net192 VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_26_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17800_ _09782_ _09786_ VGND VGND VPWR VPWR _09787_ sky130_fd_sc_hd__xor2_1
X_18780_ _10756_ _10596_ top0.pid_d.out\[9\] VGND VGND VPWR VPWR _10757_ sky130_fd_sc_hd__o21ba_1
X_15992_ _08083_ _08084_ VGND VGND VPWR VPWR _08086_ sky130_fd_sc_hd__nand2_1
X_17731_ _09716_ _09717_ VGND VGND VPWR VPWR _09718_ sky130_fd_sc_hd__and2_1
X_14943_ spi0.data_packed\[46\] top0.kid\[14\] _07086_ VGND VGND VPWR VPWR _07093_
+ sky130_fd_sc_hd__mux2_1
X_26929_ clknet_leaf_7_clk_sys _00546_ net593 VGND VGND VPWR VPWR top0.matmul0.cos\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_17662_ top0.pid_d.mult0.a\[3\] net329 VGND VGND VPWR VPWR _09649_ sky130_fd_sc_hd__nand2_1
X_14874_ spi0.data_packed\[77\] top0.kpd\[13\] _07053_ VGND VGND VPWR VPWR _07057_
+ sky130_fd_sc_hd__mux2_1
X_19401_ _11303_ _11304_ VGND VGND VPWR VPWR _11305_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16613_ _08630_ _08631_ _08632_ VGND VGND VPWR VPWR _08699_ sky130_fd_sc_hd__o21a_1
X_13825_ _05995_ _06037_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17593_ net422 net358 _09552_ VGND VGND VPWR VPWR _09580_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_35_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16544_ net510 net445 VGND VGND VPWR VPWR _08631_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19332_ net307 _11117_ _11270_ _10067_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13756_ _05967_ _05963_ _05964_ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16475_ net447 net510 VGND VGND VPWR VPWR _08563_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19263_ _11205_ _11206_ VGND VGND VPWR VPWR _11208_ sky130_fd_sc_hd__or2_1
X_13687_ _05872_ _05868_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__xor2_1
XFILLER_0_155_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18214_ _10185_ _10196_ VGND VGND VPWR VPWR _10197_ sky130_fd_sc_hd__nor2_1
X_15426_ _07523_ _07521_ _07522_ VGND VGND VPWR VPWR _07525_ sky130_fd_sc_hd__nand3_1
XFILLER_0_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19194_ top0.pid_d.curr_error\[2\] _11135_ _11144_ VGND VGND VPWR VPWR _11145_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_183_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18145_ _10097_ _10127_ VGND VGND VPWR VPWR _10129_ sky130_fd_sc_hd__and2_1
X_15357_ _07455_ VGND VGND VPWR VPWR _07456_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14308_ net36 _05551_ VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18076_ _09746_ _09821_ _10060_ VGND VGND VPWR VPWR _10061_ sky130_fd_sc_hd__a21o_1
Xhold206 top0.matmul0.matmul_stage_inst.b\[9\] VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__dlygate4sd3_1
X_15288_ _07320_ _07322_ _07374_ _07386_ _07321_ VGND VGND VPWR VPWR _07387_ sky130_fd_sc_hd__o32a_1
XPHY_EDGE_ROW_44_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold217 top0.pid_d.prev_int\[13\] VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold228 top0.cordic0.sin\[10\] VGND VGND VPWR VPWR net928 sky130_fd_sc_hd__dlygate4sd3_1
X_17027_ top0.currT_r\[13\] top0.currT_r\[14\] VGND VGND VPWR VPWR _09079_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14239_ _06417_ _06418_ _06448_ _06449_ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__a211o_1
Xhold239 top0.c_out_calc\[12\] VGND VGND VPWR VPWR net939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18978_ _10869_ _10871_ _10951_ VGND VGND VPWR VPWR _10952_ sky130_fd_sc_hd__o21a_1
X_17929_ _09909_ _09914_ VGND VGND VPWR VPWR _09915_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20940_ _12786_ _12787_ _11758_ VGND VGND VPWR VPWR _12788_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_53_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20871_ _12695_ _12718_ _12719_ VGND VGND VPWR VPWR _12720_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22610_ _02145_ _02163_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__xor2_1
XFILLER_0_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23590_ top0.matmul0.alpha_pass\[2\] _09261_ net559 VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22541_ _02095_ _02069_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25260_ _04537_ _04602_ _04601_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22472_ _02022_ _02028_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24211_ _03559_ _03566_ _03568_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__a21o_1
X_21423_ _00966_ _00989_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__xnor2_1
X_25191_ _04474_ _04532_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_62_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24142_ _03461_ _03499_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21354_ net763 _12813_ _00922_ _12963_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20305_ _12098_ _12099_ VGND VGND VPWR VPWR _12154_ sky130_fd_sc_hd__nand2_1
X_24073_ _03350_ _03428_ _03429_ _03430_ VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21285_ net248 net242 VGND VGND VPWR VPWR _13128_ sky130_fd_sc_hd__nand2_1
X_23024_ net168 top0.svm0.delta\[14\] VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__and2_1
X_20236_ net253 net249 VGND VGND VPWR VPWR _12085_ sky130_fd_sc_hd__nor2_1
XFILLER_0_200_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20167_ net207 net208 VGND VGND VPWR VPWR _12019_ sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_43_clk_sys clknet_3_7__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_43_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_200_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24975_ _04322_ _04324_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__or2_1
X_20098_ net194 _11730_ _11808_ _11936_ _11804_ VGND VGND VPWR VPWR _11957_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_71_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23926_ _03282_ _03283_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26714_ clknet_leaf_73_clk_sys _00331_ net655 VGND VGND VPWR VPWR top0.pid_d.curr_int\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26645_ clknet_leaf_75_clk_sys _00262_ net639 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_23857_ _03116_ _03117_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_197_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13610_ _05536_ _05822_ _05588_ net56 VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_196_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22808_ net170 top0.svm0.tA\[7\] VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__and2b_1
X_14590_ _06792_ _06795_ VGND VGND VPWR VPWR _06796_ sky130_fd_sc_hd__xnor2_2
X_26576_ clknet_leaf_52_clk_sys _00199_ net672 VGND VGND VPWR VPWR top0.pid_q.prev_error\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23788_ _03145_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__buf_4
XFILLER_0_67_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13541_ _05751_ _05752_ _05753_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_149_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25527_ top0.matmul0.b\[3\] top0.matmul0.matmul_stage_inst.f\[3\] _04846_ VGND VGND
+ VPWR VPWR _04850_ sky130_fd_sc_hd__mux2_1
X_22739_ net197 _02284_ net174 VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16260_ _07241_ net444 VGND VGND VPWR VPWR _08351_ sky130_fd_sc_hd__nand2_1
X_25458_ _04774_ _04800_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__xnor2_1
X_13472_ _05502_ _05503_ _05684_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__o21a_1
XFILLER_0_165_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15211_ net539 net470 VGND VGND VPWR VPWR _07310_ sky130_fd_sc_hd__nand2_2
X_24409_ _02978_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16191_ _08268_ _08282_ VGND VGND VPWR VPWR _08283_ sky130_fd_sc_hd__xnor2_4
X_25389_ _04673_ _04680_ _04681_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__o21a_1
XFILLER_0_152_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27128_ clknet_leaf_33_clk_sys _00742_ net666 VGND VGND VPWR VPWR top0.c_out_calc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_15142_ net523 VGND VGND VPWR VPWR _07241_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27059_ clknet_leaf_21_clk_sys _00676_ net610 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.d\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19950_ _11807_ _11808_ net195 net189 VGND VGND VPWR VPWR _11820_ sky130_fd_sc_hd__o211a_1
X_15073_ _07169_ _07170_ VGND VGND VPWR VPWR _07172_ sky130_fd_sc_hd__nor2_1
X_14024_ _06233_ _06236_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__xnor2_2
X_18901_ net324 net327 _10384_ VGND VGND VPWR VPWR _10876_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19881_ _11739_ _11755_ _11756_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__a21oi_1
X_18832_ _10787_ _10807_ VGND VGND VPWR VPWR _10808_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_184_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18763_ _10738_ _10739_ VGND VGND VPWR VPWR _10740_ sky130_fd_sc_hd__xnor2_1
X_15975_ _07983_ _07985_ VGND VGND VPWR VPWR _08070_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17714_ _09619_ _09700_ VGND VGND VPWR VPWR _09701_ sky130_fd_sc_hd__xnor2_2
X_14926_ spi0.data_packed\[38\] top0.kid\[6\] _07075_ VGND VGND VPWR VPWR _07084_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18694_ _10566_ _10567_ _10562_ VGND VGND VPWR VPWR _10672_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17645_ _09624_ _09631_ VGND VGND VPWR VPWR _09632_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_188_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14857_ spi0.data_packed\[69\] top0.kpd\[5\] _07042_ VGND VGND VPWR VPWR _07048_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13808_ _06019_ _06020_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__and2b_1
X_14788_ _06982_ _06988_ VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__xnor2_4
X_17576_ _09554_ _09557_ _09558_ _09562_ VGND VGND VPWR VPWR _09563_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19315_ top0.pid_d.prev_error\[14\] top0.pid_d.curr_error\[14\] VGND VGND VPWR VPWR
+ _11255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13739_ _05905_ _05904_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16527_ top0.pid_q.curr_int\[11\] _08614_ VGND VGND VPWR VPWR _08615_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19246_ _11121_ _11192_ _11125_ VGND VGND VPWR VPWR _11193_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16458_ _08543_ _08546_ VGND VGND VPWR VPWR _08547_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15409_ _07477_ _07504_ _07507_ VGND VGND VPWR VPWR _07508_ sky130_fd_sc_hd__o21a_1
X_16389_ _08411_ _08478_ VGND VGND VPWR VPWR _08479_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19177_ top0.matmul0.alpha_pass\[0\] top0.matmul0.alpha_pass\[1\] VGND VGND VPWR
+ VPWR _11130_ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18128_ _10102_ _10111_ VGND VGND VPWR VPWR _10112_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18059_ _09942_ _09944_ _10043_ VGND VGND VPWR VPWR _10044_ sky130_fd_sc_hd__a21o_1
X_21070_ _12094_ _12915_ net272 VGND VGND VPWR VPWR _12916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout505 top0.pid_q.mult0.a\[13\] VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__clkbuf_4
Xfanout516 top0.pid_q.mult0.a\[9\] VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__buf_4
X_20021_ _11880_ _11886_ VGND VGND VPWR VPWR _11887_ sky130_fd_sc_hd__xnor2_1
Xfanout527 top0.pid_q.mult0.a\[5\] VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_171_Right_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout538 net539 VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__buf_4
Xfanout549 net552 VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__clkbuf_4
X_24760_ _04021_ _04022_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__or2_1
X_21972_ _01474_ _01475_ net166 VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23711_ _03068_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__clkbuf_4
X_20923_ _12769_ _12770_ VGND VGND VPWR VPWR _12771_ sky130_fd_sc_hd__or2_1
XFILLER_0_179_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24691_ _04039_ _04041_ _04043_ _03935_ _04044_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__o32a_2
XFILLER_0_96_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26430_ clknet_leaf_77_clk_sys _00071_ net631 VGND VGND VPWR VPWR top0.kid\[3\] sky130_fd_sc_hd__dfrtp_1
X_23642_ _02999_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__clkbuf_4
X_20854_ net239 net235 VGND VGND VPWR VPWR _12703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26361_ _05412_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__clkbuf_1
X_23573_ _02953_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20785_ net300 net292 net278 VGND VGND VPWR VPWR _12634_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25312_ _04655_ _04657_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__nand2_1
X_22524_ _02077_ _02079_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26292_ net925 spi0.data_packed\[45\] net693 VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25243_ _04588_ _04589_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22455_ _01292_ net114 _01770_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21406_ _12762_ _12764_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__nand2_1
X_25174_ _04177_ _04521_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_150_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22386_ _01896_ _01944_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__xor2_1
X_24125_ _03323_ _03056_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21337_ _13176_ _13178_ VGND VGND VPWR VPWR _13179_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24056_ _03372_ _03375_ _03374_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__a21o_1
X_21268_ _13027_ _13033_ _13038_ VGND VGND VPWR VPWR _13111_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_198_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23007_ _06277_ _02511_ net171 VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20219_ _12065_ _12067_ VGND VGND VPWR VPWR _12068_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21199_ _13040_ _13042_ VGND VGND VPWR VPWR _13043_ sky130_fd_sc_hd__xnor2_1
X_15760_ _07739_ _07740_ _07856_ VGND VGND VPWR VPWR _07857_ sky130_fd_sc_hd__a21oi_2
X_24958_ _04226_ _04231_ _04308_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__a21o_1
X_14711_ _06889_ _06890_ VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__nand2_1
X_23909_ _03256_ _03262_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__xnor2_2
X_15691_ _07660_ _07787_ _07788_ VGND VGND VPWR VPWR _07789_ sky130_fd_sc_hd__a21oi_2
X_24889_ _04168_ _04240_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14642_ _06716_ _06846_ VGND VGND VPWR VPWR _06847_ sky130_fd_sc_hd__xor2_1
X_17430_ _09415_ _09416_ VGND VGND VPWR VPWR _09417_ sky130_fd_sc_hd__xor2_2
X_26628_ clknet_leaf_72_clk_sys _00245_ net655 VGND VGND VPWR VPWR top0.pid_d.out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_200_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14573_ _06640_ _06778_ net23 VGND VGND VPWR VPWR _06779_ sky130_fd_sc_hd__mux2_1
X_17361_ _09346_ _09347_ VGND VGND VPWR VPWR _09348_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_109_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26559_ clknet_leaf_51_clk_sys _00182_ net670 VGND VGND VPWR VPWR top0.pid_q.curr_error\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19100_ _11068_ _11071_ VGND VGND VPWR VPWR _11072_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13524_ net1025 _05602_ _05603_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__and3_1
X_16312_ _08402_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__clkbuf_1
X_17292_ _09286_ _09282_ _09287_ VGND VGND VPWR VPWR _09288_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16243_ _08304_ _08332_ _08333_ VGND VGND VPWR VPWR _08334_ sky130_fd_sc_hd__o21a_1
X_19031_ net314 net365 VGND VGND VPWR VPWR _11004_ sky130_fd_sc_hd__nand2_1
X_13455_ net63 _05619_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_180_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16174_ _08262_ _08265_ VGND VGND VPWR VPWR _08266_ sky130_fd_sc_hd__xnor2_2
X_13386_ top0.svm0.state\[1\] top0.svm0.state\[0\] top0.matmul0.alpha_pass\[10\] VGND
+ VGND VPWR VPWR _05599_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_24_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15125_ net514 net494 net490 net517 VGND VGND VPWR VPWR _07224_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19933_ net201 net184 net190 VGND VGND VPWR VPWR _11804_ sky130_fd_sc_hd__or3_1
X_15056_ net531 net470 VGND VGND VPWR VPWR _07155_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_118_Left_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14007_ _05894_ _05497_ _06215_ _06216_ _06219_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__o2111a_2
X_19864_ net82 _11535_ _11730_ VGND VGND VPWR VPWR _11740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18815_ _10790_ net368 net327 VGND VGND VPWR VPWR _10791_ sky130_fd_sc_hd__a21o_1
X_19795_ _11448_ _11442_ _11675_ VGND VGND VPWR VPWR _11676_ sky130_fd_sc_hd__o21a_1
XFILLER_0_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18746_ _10722_ VGND VGND VPWR VPWR _10723_ sky130_fd_sc_hd__inv_2
X_15958_ _08045_ _08052_ VGND VGND VPWR VPWR _08053_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_179_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14909_ _07041_ VGND VGND VPWR VPWR _07075_ sky130_fd_sc_hd__buf_4
X_18677_ _10629_ _10654_ VGND VGND VPWR VPWR _10655_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_144_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15889_ _07876_ _07878_ _07984_ VGND VGND VPWR VPWR _07985_ sky130_fd_sc_hd__a21o_1
XFILLER_0_187_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17628_ net1023 _09613_ _09614_ VGND VGND VPWR VPWR _09615_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_127_Left_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17559_ _09386_ _09545_ VGND VGND VPWR VPWR _09546_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20570_ _12359_ _12384_ _12401_ _12402_ _12418_ VGND VGND VPWR VPWR _12419_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_34_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19229_ _11175_ _11176_ VGND VGND VPWR VPWR _11177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22240_ _01221_ _01797_ _01800_ _01691_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_108_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22171_ _01165_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21122_ _12914_ _12919_ _12966_ VGND VGND VPWR VPWR _12967_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_111_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout302 net305 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25930_ _08899_ _05140_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__nor2_1
X_21053_ _12843_ _12898_ _12859_ VGND VGND VPWR VPWR _12899_ sky130_fd_sc_hd__a21oi_2
Xfanout313 top0.pid_d.mult0.b\[13\] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__buf_2
Xfanout324 net325 VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__clkbuf_2
Xfanout335 net336 VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__clkbuf_2
Xfanout346 top0.pid_d.mult0.b\[3\] VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_185_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout357 net358 VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__clkbuf_4
X_20004_ _11431_ _11870_ net177 VGND VGND VPWR VPWR _11871_ sky130_fd_sc_hd__o21ai_1
X_25861_ _05070_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__inv_2
Xfanout368 top0.pid_d.mult0.a\[14\] VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_185_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout379 net380 VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__buf_2
X_24812_ _04143_ _04163_ _04141_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__o21a_1
XFILLER_0_198_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25792_ net208 _05009_ _05021_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__and3_1
XFILLER_0_154_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24743_ _04013_ _04014_ _04095_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__o21a_1
XFILLER_0_201_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21955_ net156 net130 VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20906_ _12101_ _12715_ VGND VGND VPWR VPWR _12754_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24674_ _04011_ _04012_ _04027_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__a21boi_1
X_21886_ _01397_ _01403_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23625_ _02978_ _02982_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__nor2_2
X_26413_ clknet_leaf_61_clk_sys _00054_ net650 VGND VGND VPWR VPWR top0.kpq\[2\] sky130_fd_sc_hd__dfrtp_1
X_20837_ _12678_ _12679_ _12685_ VGND VGND VPWR VPWR _12686_ sky130_fd_sc_hd__a21o_1
X_26344_ spi0.data_packed\[70\] spi0.data_packed\[71\] net689 VGND VGND VPWR VPWR
+ _05404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23556_ _02944_ VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20768_ _12609_ _12610_ _12616_ VGND VGND VPWR VPWR _12617_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_92_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22507_ _01217_ _01784_ _02062_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_174_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26275_ _05369_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23487_ _02908_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20699_ net300 _12491_ VGND VGND VPWR VPWR _12548_ sky130_fd_sc_hd__xnor2_1
X_25226_ _04496_ _04502_ _04501_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__a21oi_2
X_13240_ top0.matmul0.matmul_stage_inst.state\[0\] top0.matmul0.matmul_stage_inst.start
+ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__nand2_4
X_22438_ _01987_ _01995_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_162_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25157_ _04492_ _04504_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22369_ _01923_ _01927_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24108_ _03463_ _03462_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__nor2_1
X_25088_ _03325_ _03908_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__nor2_2
XFILLER_0_202_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24039_ _03387_ _03392_ _03396_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__a21o_1
X_16930_ _08988_ _08977_ top0.pid_q.prev_error\[7\] VGND VGND VPWR VPWR _08989_ sky130_fd_sc_hd__o21ba_1
X_16861_ _08922_ _08924_ VGND VGND VPWR VPWR _08925_ sky130_fd_sc_hd__and2_1
X_18600_ _10573_ _10578_ VGND VGND VPWR VPWR _10579_ sky130_fd_sc_hd__xnor2_4
X_15812_ net474 net509 VGND VGND VPWR VPWR _07908_ sky130_fd_sc_hd__nand2_2
X_19580_ top0.cordic0.slte0.opB\[14\] top0.cordic0.slte0.opA\[14\] VGND VGND VPWR
+ VPWR _11469_ sky130_fd_sc_hd__and2b_1
X_16792_ net527 _08856_ _08859_ net793 _08869_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__a221o_1
XFILLER_0_172_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18531_ _05449_ _10510_ VGND VGND VPWR VPWR _10511_ sky130_fd_sc_hd__and2_1
X_15743_ net448 _07838_ _07839_ VGND VGND VPWR VPWR _07840_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_99_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18462_ _10346_ _10415_ VGND VGND VPWR VPWR _10442_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15674_ net481 _07771_ VGND VGND VPWR VPWR _07772_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17413_ net400 _09360_ _09399_ net352 VGND VGND VPWR VPWR _09400_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_200_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14625_ _06766_ _06771_ _06764_ VGND VGND VPWR VPWR _06830_ sky130_fd_sc_hd__o21ba_1
X_18393_ net324 net381 VGND VGND VPWR VPWR _10374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14556_ net25 _05640_ VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__nand2_1
X_17344_ _09332_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13507_ top0.matmul0.beta_pass\[14\] _05436_ _05719_ _05464_ top0.c_out_calc\[14\]
+ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__a32o_1
XFILLER_0_125_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14487_ _06661_ _06692_ VGND VGND VPWR VPWR _06694_ sky130_fd_sc_hd__nor2_1
X_17275_ _09273_ VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19014_ _10986_ _10987_ VGND VGND VPWR VPWR _10988_ sky130_fd_sc_hd__xnor2_1
X_13438_ _05643_ _05636_ _05650_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__o21ai_2
X_16226_ _08317_ VGND VGND VPWR VPWR _08318_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16157_ _08088_ _08161_ _08162_ _08232_ VGND VGND VPWR VPWR _08249_ sky130_fd_sc_hd__a211o_1
X_13369_ _05580_ _05581_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_139_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15108_ _07205_ _07206_ VGND VGND VPWR VPWR _07207_ sky130_fd_sc_hd__xnor2_1
X_16088_ _08179_ _08180_ VGND VGND VPWR VPWR _08181_ sky130_fd_sc_hd__or2_1
X_19916_ _11788_ VGND VGND VPWR VPWR _11789_ sky130_fd_sc_hd__buf_4
X_15039_ net990 _07140_ _07144_ top0.pid_d.curr_int\[9\] VGND VGND VPWR VPWR _00126_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19847_ _11723_ _11724_ net241 VGND VGND VPWR VPWR _11725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19778_ net181 net82 _11659_ net182 VGND VGND VPWR VPWR _11660_ sky130_fd_sc_hd__a22o_1
X_18729_ _10704_ _10705_ VGND VGND VPWR VPWR _10706_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21740_ _01266_ _01299_ _01301_ net152 _01102_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__a32o_1
XFILLER_0_188_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21671_ _01117_ _01120_ _01126_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__a21o_1
XFILLER_0_164_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23410_ _02847_ _02848_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20622_ _12469_ _12470_ VGND VGND VPWR VPWR _12471_ sky130_fd_sc_hd__nor2_2
XFILLER_0_171_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24390_ _03745_ _03746_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23341_ net128 _02774_ _02783_ _02784_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__o211a_1
X_20553_ _12399_ _12400_ VGND VGND VPWR VPWR _12402_ sky130_fd_sc_hd__nor2_1
X_26060_ top0.pid_d.out\[7\] _05232_ _05233_ spi0.data_packed\[71\] VGND VGND VPWR
+ VPWR _05247_ sky130_fd_sc_hd__a22o_1
X_23272_ _02707_ _02719_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20484_ _12059_ net302 _12057_ VGND VGND VPWR VPWR _12333_ sky130_fd_sc_hd__and3b_1
XFILLER_0_6_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25011_ _04352_ _04360_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22223_ _01777_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22154_ net114 _01075_ _01260_ _01715_ _01133_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__a221o_2
XFILLER_0_121_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21105_ _12808_ _12942_ _12950_ VGND VGND VPWR VPWR _12951_ sky130_fd_sc_hd__a21boi_2
X_26962_ clknet_leaf_14_clk_sys _00579_ net617 VGND VGND VPWR VPWR top0.matmul0.b\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_22085_ _01640_ _01645_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__nand2_1
Xfanout110 net112 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__buf_2
Xfanout121 top0.cordic0.vec\[1\]\[9\] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__buf_4
Xfanout132 net134 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
X_25913_ top0.matmul0.alpha_pass\[12\] top0.matmul0.beta_pass\[12\] VGND VGND VPWR
+ VPWR _05129_ sky130_fd_sc_hd__xnor2_2
Xfanout143 top0.cordic0.vec\[1\]\[4\] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_4
X_21036_ _12743_ VGND VGND VPWR VPWR _12883_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout154 net157 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_201_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout165 net167 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_2
X_26893_ clknet_leaf_107_clk_sys _00510_ net577 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout176 net178 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout187 net188 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_4
X_25844_ net76 top0.matmul0.beta_pass\[5\] _05058_ _05059_ VGND VGND VPWR VPWR _05066_
+ sky130_fd_sc_hd__nor4_1
Xfanout198 net200 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_4
XFILLER_0_199_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22987_ _06277_ _02494_ net172 VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__o21ai_1
X_25775_ _05008_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24726_ _03983_ _03988_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__nor2_1
X_21938_ _01495_ _01497_ _01499_ net162 VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__o22a_1
XFILLER_0_96_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24657_ _04007_ _04008_ _04009_ _04010_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_78_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21869_ _01409_ _01430_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__xor2_1
XFILLER_0_49_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14410_ _06616_ _06617_ VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_166_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23608_ top0.matmul0.alpha_pass\[11\] _09314_ net559 VGND VGND VPWR VPWR _02971_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15390_ _07482_ _07486_ _07476_ _07488_ VGND VGND VPWR VPWR _07489_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_182_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24588_ _03830_ _03940_ _03941_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14341_ _06549_ _06544_ _06543_ VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__o21ba_1
X_26327_ _05395_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__clkbuf_1
X_23539_ _02935_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17060_ top0.pid_q.curr_error\[6\] _09100_ _09102_ _08962_ VGND VGND VPWR VPWR _00187_
+ sky130_fd_sc_hd__a22o_1
X_14272_ _06408_ _06415_ _06416_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__a21boi_4
X_26258_ spi0.data_packed\[27\] spi0.data_packed\[28\] net699 VGND VGND VPWR VPWR
+ _05361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16011_ _08099_ _08104_ VGND VGND VPWR VPWR _08105_ sky130_fd_sc_hd__xor2_1
X_25209_ _03981_ _03123_ _03889_ _03758_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13223_ _05446_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__clkbuf_1
X_26189_ _05323_ top0.cordic0.slte0.opB\[13\] _12003_ VGND VGND VPWR VPWR _05324_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17962_ _09939_ _09947_ VGND VGND VPWR VPWR _09948_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19701_ _11544_ _11551_ _11567_ net292 VGND VGND VPWR VPWR _11587_ sky130_fd_sc_hd__a22oi_2
X_16913_ top0.currT_r\[7\] _08972_ VGND VGND VPWR VPWR _08973_ sky130_fd_sc_hd__xnor2_1
X_17893_ _09859_ _09879_ VGND VGND VPWR VPWR _09880_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19632_ _11424_ _11516_ _11520_ VGND VGND VPWR VPWR _11521_ sky130_fd_sc_hd__and3_1
X_16844_ top0.pid_q.prev_error\[1\] top0.pid_q.curr_error\[1\] top0.pid_q.prev_error\[0\]
+ top0.pid_q.curr_error\[0\] VGND VGND VPWR VPWR _08909_ sky130_fd_sc_hd__o211ai_2
Xclkbuf_leaf_91_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_91_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_192_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19563_ _11443_ _11445_ _11449_ _11450_ _11451_ VGND VGND VPWR VPWR _11452_ sky130_fd_sc_hd__a32oi_4
X_16775_ _08857_ VGND VGND VPWR VPWR _08858_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_87_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13987_ _06099_ _06199_ _06093_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18514_ _10103_ VGND VGND VPWR VPWR _10494_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15726_ _07821_ _07822_ VGND VGND VPWR VPWR _07823_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19494_ net441 _11386_ VGND VGND VPWR VPWR _11387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18445_ _05449_ _10425_ VGND VGND VPWR VPWR _10426_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15657_ net454 net532 VGND VGND VPWR VPWR _07755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14608_ _06800_ _06810_ _06697_ VGND VGND VPWR VPWR _06813_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18376_ _10355_ _10356_ VGND VGND VPWR VPWR _10357_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15588_ _07684_ _07686_ VGND VGND VPWR VPWR _07687_ sky130_fd_sc_hd__xor2_1
X_17327_ _09312_ _09316_ _09317_ VGND VGND VPWR VPWR _09318_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_161_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14539_ _06740_ _06745_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__xor2_2
XFILLER_0_172_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17258_ _09257_ _09258_ VGND VGND VPWR VPWR _09259_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16209_ _08298_ _08300_ VGND VGND VPWR VPWR _08301_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17189_ top0.pid_q.curr_int\[8\] _09140_ _09199_ _09135_ VGND VGND VPWR VPWR _09200_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22910_ _02374_ top0.svm0.tC\[12\] top0.svm0.tC\[11\] _02345_ _02427_ VGND VGND VPWR
+ VPWR _02428_ sky130_fd_sc_hd__a221o_1
X_23890_ _03061_ _03062_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__or2_2
X_22841_ top0.svm0.counter\[5\] _02323_ _02327_ _02328_ _02329_ VGND VGND VPWR VPWR
+ _02361_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_190_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25560_ _05456_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22772_ _07115_ _06276_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24511_ _03004_ _03005_ _03090_ _03091_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__o22a_1
XFILLER_0_52_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21723_ _01277_ _01284_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__nor2_1
X_25491_ _04831_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24442_ _03724_ _03729_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27230_ clknet_3_1__leaf_clk_mosi _00844_ VGND VGND VPWR VPWR spi0.data_packed\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21654_ net143 net139 VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_191_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20605_ _12447_ _12451_ _12453_ VGND VGND VPWR VPWR _12454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27161_ clknet_leaf_9_clk_sys _00775_ net596 VGND VGND VPWR VPWR top0.a_in_matmul\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_24373_ _03724_ _03729_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21585_ net164 net143 VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__and2b_1
XFILLER_0_34_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26112_ _05277_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_132_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23324_ _02709_ _02713_ net187 VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__mux2_1
X_27092_ clknet_leaf_22_clk_sys _00709_ net608 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_20536_ _12359_ _12384_ VGND VGND VPWR VPWR _12385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26043_ top0.pid_d.out\[3\] _05232_ _05233_ spi0.data_packed\[67\] VGND VGND VPWR
+ VPWR _05234_ sky130_fd_sc_hd__a22o_1
X_23255_ net165 _11511_ _02679_ _02683_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__a31o_1
X_20467_ _12296_ _12297_ _12315_ VGND VGND VPWR VPWR _12316_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22206_ _01102_ _01100_ _01766_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23186_ _02646_ _06612_ _02649_ net823 VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__a22o_1
X_20398_ _11727_ _12246_ VGND VGND VPWR VPWR _12247_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22137_ _01139_ _01208_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22068_ net118 net106 net102 _01563_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__a31o_1
X_26945_ clknet_leaf_8_clk_sys _00562_ net595 VGND VGND VPWR VPWR top0.matmul0.a\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13910_ _06119_ _06120_ _06121_ _06122_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__o211a_1
X_21019_ _12782_ _12800_ VGND VGND VPWR VPWR _12866_ sky130_fd_sc_hd__nor2_1
X_26876_ clknet_leaf_42_clk_sys _00493_ net684 VGND VGND VPWR VPWR top0.svm0.tB\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14890_ _07065_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25827_ _05043_ _05044_ _05047_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__a21o_1
X_13841_ net62 net59 _06047_ _05497_ net68 VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__a32o_1
XFILLER_0_159_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16560_ _08554_ _08555_ _08646_ VGND VGND VPWR VPWR _08647_ sky130_fd_sc_hd__a21o_1
X_13772_ _05968_ _05984_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__or2_1
X_25758_ net70 top0.matmul0.cos\[7\] _05458_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15511_ _07255_ _07601_ VGND VGND VPWR VPWR _07610_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24709_ top0.matmul0.matmul_stage_inst.mult2\[4\] _04062_ _03642_ VGND VGND VPWR
+ VPWR _04063_ sky130_fd_sc_hd__mux2_1
X_16491_ _08567_ _08578_ VGND VGND VPWR VPWR _08579_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_139_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25689_ top0.matmul0.sin\[13\] _04955_ _04956_ net72 _04896_ VGND VGND VPWR VPWR
+ _04957_ sky130_fd_sc_hd__o221a_1
XFILLER_0_183_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18230_ net415 top0.pid_d.mult0.b\[14\] VGND VGND VPWR VPWR _10213_ sky130_fd_sc_hd__nand2_2
XFILLER_0_155_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15442_ net480 _07540_ VGND VGND VPWR VPWR _07541_ sky130_fd_sc_hd__nand2_1
X_18161_ _10137_ _10143_ VGND VGND VPWR VPWR _10145_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15373_ _07469_ _07471_ VGND VGND VPWR VPWR _07472_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_38_clk_sys clknet_3_7__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_38_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17112_ net728 _09114_ _09132_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__a21o_1
X_14324_ _06455_ _06456_ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__and2b_1
XFILLER_0_135_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18092_ net405 net318 VGND VGND VPWR VPWR _10076_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14255_ _06349_ _06465_ _06348_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_151_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17043_ net546 _09090_ _09094_ _08882_ VGND VGND VPWR VPWR _09095_ sky130_fd_sc_hd__a211o_1
XFILLER_0_52_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13206_ top0.matmul0.start VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14186_ _06395_ _06396_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__xor2_1
XFILLER_0_150_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18994_ _10965_ _10967_ net380 VGND VGND VPWR VPWR _10968_ sky130_fd_sc_hd__mux2_1
X_17945_ _09916_ _09930_ VGND VGND VPWR VPWR _09931_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17876_ net361 net372 VGND VGND VPWR VPWR _09863_ sky130_fd_sc_hd__nand2_2
X_19615_ _11491_ _11493_ _11495_ _11496_ _11503_ VGND VGND VPWR VPWR _11504_ sky130_fd_sc_hd__o221a_4
X_16827_ _05439_ _08892_ VGND VGND VPWR VPWR _08893_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19546_ net306 _11424_ _11435_ VGND VGND VPWR VPWR _11436_ sky130_fd_sc_hd__and3_1
X_16758_ _08840_ _08841_ _08745_ VGND VGND VPWR VPWR _08842_ sky130_fd_sc_hd__mux2_2
XFILLER_0_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15709_ top0.pid_q.out\[2\] _07801_ _07805_ VGND VGND VPWR VPWR _07806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19477_ net441 _11370_ _11371_ _11231_ VGND VGND VPWR VPWR _11372_ sky130_fd_sc_hd__a31o_1
X_16689_ _08648_ _08773_ VGND VGND VPWR VPWR _08774_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_146_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18428_ _10402_ _10408_ VGND VGND VPWR VPWR _10409_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_186_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18359_ top0.pid_d.out\[6\] top0.pid_d.curr_int\[6\] VGND VGND VPWR VPWR _10340_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21370_ _00937_ _12820_ _13170_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20321_ _12153_ _12169_ VGND VGND VPWR VPWR _12170_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23040_ net46 net44 top0.periodTop_r\[9\] _02540_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__or4_1
X_20252_ net271 net265 VGND VGND VPWR VPWR _12101_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_12_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20183_ top0.state\[1\] _12026_ VGND VGND VPWR VPWR _12033_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24991_ _04069_ _04340_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__xnor2_1
X_26730_ clknet_leaf_100_clk_sys _00347_ net576 VGND VGND VPWR VPWR top0.cordic0.vec\[0\]\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_192_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23942_ _03229_ _03230_ _03298_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__and3_1
XFILLER_0_193_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23873_ _03098_ _03134_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__xnor2_4
X_26661_ clknet_leaf_75_clk_sys _00278_ net637 VGND VGND VPWR VPWR top0.pid_d.mult0.b\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_193_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22824_ _02340_ _02341_ _02342_ _02343_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__or4b_1
X_25612_ net70 top0.matmul0.cos\[9\] VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26592_ clknet_leaf_65_clk_sys _00215_ net657 VGND VGND VPWR VPWR top0.pid_q.curr_int\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25543_ _04858_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__clkbuf_1
X_22755_ _02294_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21706_ net152 net146 VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__and2b_1
X_25474_ _04717_ _04814_ _04816_ _04712_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22686_ _02223_ _02236_ _02206_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_176_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24425_ _03774_ _03780_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27213_ clknet_leaf_87_clk_sys _00827_ net642 VGND VGND VPWR VPWR top0.ready sky130_fd_sc_hd__dfstp_1
X_21637_ _01106_ _01107_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__nor2_1
XFILLER_0_191_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24356_ _03709_ _03712_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__xnor2_2
X_27144_ clknet_leaf_31_clk_sys _00758_ net617 VGND VGND VPWR VPWR top0.b_in_matmul\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21568_ _01099_ _01129_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_185_Right_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23307_ _11425_ net215 _02750_ _11576_ _02752_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__o221a_2
X_27075_ clknet_leaf_22_clk_sys _00692_ net607 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.c\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_20519_ _12363_ _12365_ _12266_ VGND VGND VPWR VPWR _12368_ sky130_fd_sc_hd__mux2_1
X_24287_ _03624_ _03625_ _03630_ _03300_ _03299_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__a2111oi_1
X_21499_ _12037_ _01060_ _01061_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__o21ai_1
X_14040_ _06251_ _06252_ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__and2b_1
X_26026_ top0.b_in_matmul\[15\] _05220_ _05196_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__mux2_1
X_23238_ net249 net244 net243 net237 net198 net192 VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__mux4_2
XFILLER_0_105_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23169_ _02641_ _06799_ _02645_ net788 VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__a22o_1
X_15991_ _08083_ _08084_ VGND VGND VPWR VPWR _08085_ sky130_fd_sc_hd__or2_1
X_17730_ _09714_ _09715_ _09686_ VGND VGND VPWR VPWR _09717_ sky130_fd_sc_hd__o21ai_1
X_14942_ _07092_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__clkbuf_1
X_26928_ clknet_leaf_7_clk_sys _00545_ net592 VGND VGND VPWR VPWR top0.matmul0.cos\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_17661_ net322 net424 VGND VGND VPWR VPWR _09648_ sky130_fd_sc_hd__nand2_1
X_26859_ clknet_leaf_36_clk_sys _00476_ net678 VGND VGND VPWR VPWR top0.svm0.tA\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14873_ _07056_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__clkbuf_1
X_19400_ top0.pid_d.curr_int\[2\] top0.pid_d.prev_int\[2\] VGND VGND VPWR VPWR _11304_
+ sky130_fd_sc_hd__xnor2_1
X_16612_ _08695_ _08697_ VGND VGND VPWR VPWR _08698_ sky130_fd_sc_hd__xor2_1
XFILLER_0_199_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13824_ _06016_ _06015_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__and2_1
X_17592_ _09522_ _09575_ _09577_ net347 _09578_ VGND VGND VPWR VPWR _09579_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19331_ net438 _11268_ _11269_ _11120_ _11123_ VGND VGND VPWR VPWR _11270_ sky130_fd_sc_hd__a221o_1
XFILLER_0_187_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16543_ net1029 net444 VGND VGND VPWR VPWR _08630_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_97_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13755_ _05963_ _05964_ _05967_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_202_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19262_ _11205_ _11206_ VGND VGND VPWR VPWR _11207_ sky130_fd_sc_hd__nand2_1
X_16474_ net1029 top0.pid_q.mult0.b\[14\] VGND VGND VPWR VPWR _08562_ sky130_fd_sc_hd__nand2_1
X_13686_ _05889_ _05892_ _05898_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18213_ _10190_ _10195_ VGND VGND VPWR VPWR _10196_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15425_ _07521_ _07522_ _07523_ VGND VGND VPWR VPWR _07524_ sky130_fd_sc_hd__a21o_1
XFILLER_0_183_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19193_ top0.pid_d.curr_error\[2\] _11133_ _11134_ top0.pid_d.prev_error\[2\] VGND
+ VGND VPWR VPWR _11144_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18144_ _10097_ _10127_ VGND VGND VPWR VPWR _10128_ sky130_fd_sc_hd__nor2_1
X_15356_ net531 net493 VGND VGND VPWR VPWR _07455_ sky130_fd_sc_hd__and2_1
XFILLER_0_198_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14307_ net31 _05586_ VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18075_ _09972_ _09974_ _09822_ _09891_ VGND VGND VPWR VPWR _10060_ sky130_fd_sc_hd__a211o_1
X_15287_ _07385_ net525 _07374_ VGND VGND VPWR VPWR _07386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold207 top0.currT_r\[0\] VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold218 top0.currT_r\[4\] VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17026_ net445 _08890_ _09078_ _08930_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__o211a_1
Xhold229 top0.pid_q.curr_error\[4\] VGND VGND VPWR VPWR net929 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ _06446_ _06447_ _06419_ _06420_ VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_145_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14169_ _05465_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18977_ net365 _10863_ _10869_ _10871_ VGND VGND VPWR VPWR _10951_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17928_ _09910_ _09913_ VGND VGND VPWR VPWR _09914_ sky130_fd_sc_hd__xnor2_2
X_17859_ net342 net388 VGND VGND VPWR VPWR _09846_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20870_ _12717_ _12711_ _12712_ VGND VGND VPWR VPWR _12719_ sky130_fd_sc_hd__nand3_1
XFILLER_0_178_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19529_ net187 VGND VGND VPWR VPWR _11419_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22540_ _02053_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22471_ _02026_ _02027_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24210_ _03567_ _03552_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_161_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21422_ _00987_ _00988_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__nand2_1
X_25190_ _04474_ _04532_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24141_ _03462_ _03465_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21353_ _13155_ _00921_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20304_ _12125_ _12152_ VGND VGND VPWR VPWR _12153_ sky130_fd_sc_hd__xnor2_1
X_24072_ _03424_ _03426_ _03374_ VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__and3_1
X_21284_ _13123_ _13126_ VGND VGND VPWR VPWR _13127_ sky130_fd_sc_hd__xnor2_2
X_23023_ net168 _02524_ _02525_ _02523_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__a22o_1
X_20235_ _12070_ _12071_ _12083_ VGND VGND VPWR VPWR _12084_ sky130_fd_sc_hd__a21oi_2
X_20166_ _12017_ VGND VGND VPWR VPWR _12018_ sky130_fd_sc_hd__inv_2
XFILLER_0_200_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24974_ _04322_ _04324_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__nand2_1
X_20097_ _11956_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__clkbuf_1
X_26713_ clknet_leaf_72_clk_sys _00330_ net663 VGND VGND VPWR VPWR top0.pid_d.curr_int\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_23925_ _03144_ _03153_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26644_ clknet_leaf_86_clk_sys _00261_ net640 VGND VGND VPWR VPWR top0.pid_d.out_valid
+ sky130_fd_sc_hd__dfrtp_1
X_23856_ _03116_ _03117_ _03112_ _03113_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_54_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22807_ _02325_ _02326_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__or2_1
X_26575_ clknet_leaf_52_clk_sys _00198_ net671 VGND VGND VPWR VPWR top0.pid_q.prev_error\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23787_ net571 net575 VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__or2_1
X_20999_ _11592_ _12844_ _12845_ VGND VGND VPWR VPWR _12846_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13540_ _05708_ _05693_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__or2_1
X_25526_ _04849_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22738_ net197 _11526_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13471_ net35 _05683_ _05503_ _05505_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__a31o_1
X_25457_ _04796_ _04799_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__xnor2_1
X_22669_ _02219_ _02220_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15210_ _07305_ _07306_ _07308_ VGND VGND VPWR VPWR _07309_ sky130_fd_sc_hd__a21o_1
X_24408_ _03502_ _03158_ _03681_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16190_ _08270_ _08281_ VGND VGND VPWR VPWR _08282_ sky130_fd_sc_hd__xor2_2
X_25388_ _04726_ _04731_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_35_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27127_ clknet_leaf_33_clk_sys _00741_ net666 VGND VGND VPWR VPWR top0.c_out_calc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15141_ _07186_ _07237_ _07239_ VGND VGND VPWR VPWR _07240_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24339_ _03184_ _03190_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15072_ _07169_ _07170_ VGND VGND VPWR VPWR _07171_ sky130_fd_sc_hd__nand2_1
X_27058_ clknet_leaf_20_clk_sys _00675_ net610 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.d\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14023_ _06109_ _06234_ _06235_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_121_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18900_ _10861_ _10874_ VGND VGND VPWR VPWR _10875_ sky130_fd_sc_hd__xnor2_4
X_26009_ top0.matmul0.beta_pass\[11\] _05203_ _05207_ VGND VGND VPWR VPWR _05208_
+ sky130_fd_sc_hd__a21o_1
X_19880_ net232 _11435_ _11754_ VGND VGND VPWR VPWR _11756_ sky130_fd_sc_hd__and3_1
X_18831_ _10789_ _10806_ VGND VGND VPWR VPWR _10807_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18762_ _09688_ _09459_ _10228_ VGND VGND VPWR VPWR _10739_ sky130_fd_sc_hd__or3_2
XFILLER_0_93_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15974_ _07985_ _07983_ VGND VGND VPWR VPWR _08069_ sky130_fd_sc_hd__or2b_1
XFILLER_0_175_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17713_ _09632_ _09633_ VGND VGND VPWR VPWR _09700_ sky130_fd_sc_hd__xor2_1
X_14925_ _07083_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__clkbuf_1
X_18693_ _10559_ _10571_ _10570_ VGND VGND VPWR VPWR _10671_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold90 top0.svm0.tB\[11\] VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__dlygate4sd3_1
X_17644_ _09627_ _09630_ VGND VGND VPWR VPWR _09631_ sky130_fd_sc_hd__xnor2_1
X_14856_ _07047_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13807_ _06003_ _06009_ _05995_ VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__a21bo_1
X_17575_ net359 _09560_ _09431_ _09561_ VGND VGND VPWR VPWR _09562_ sky130_fd_sc_hd__a22oi_4
X_14787_ _06964_ _06985_ _06987_ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_133_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19314_ top0.pid_d.prev_error\[14\] top0.pid_d.curr_error\[14\] VGND VGND VPWR VPWR
+ _11254_ sky130_fd_sc_hd__and2_1
XFILLER_0_202_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16526_ _08486_ _08612_ _08613_ VGND VGND VPWR VPWR _08614_ sky130_fd_sc_hd__o21ai_2
X_13738_ _05905_ _05904_ _05878_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19245_ _11190_ _11191_ VGND VGND VPWR VPWR _11192_ sky130_fd_sc_hd__and2_1
X_16457_ _08467_ _08471_ _08545_ _08142_ VGND VGND VPWR VPWR _08546_ sky130_fd_sc_hd__o2bb2a_1
X_13669_ _05832_ _05844_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15408_ net541 _07505_ _07506_ _07478_ VGND VGND VPWR VPWR _07507_ sky130_fd_sc_hd__a22o_1
X_19176_ _11127_ _11128_ net439 VGND VGND VPWR VPWR _11129_ sky130_fd_sc_hd__o21a_1
X_16388_ _08474_ _08477_ VGND VGND VPWR VPWR _08478_ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18127_ _10105_ _10110_ VGND VGND VPWR VPWR _10111_ sky130_fd_sc_hd__xnor2_1
X_15339_ net534 net487 VGND VGND VPWR VPWR _07438_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18058_ _09942_ _09944_ _09943_ VGND VGND VPWR VPWR _10043_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17009_ net547 _09062_ VGND VGND VPWR VPWR _09063_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout506 top0.pid_q.mult0.a\[12\] VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20020_ _11883_ _11885_ VGND VGND VPWR VPWR _11886_ sky130_fd_sc_hd__nor2_1
Xfanout517 net518 VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__clkbuf_4
Xfanout528 top0.pid_q.mult0.a\[4\] VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__buf_4
Xfanout539 top0.pid_q.mult0.a\[1\] VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__buf_4
XFILLER_0_67_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21971_ _01528_ _01532_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23710_ net571 net574 top0.matmul0.matmul_stage_inst.f\[8\] VGND VGND VPWR VPWR _03068_
+ sky130_fd_sc_hd__o21a_1
X_20922_ net218 net224 VGND VGND VPWR VPWR _12770_ sky130_fd_sc_hd__and2b_1
XFILLER_0_83_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24690_ _04042_ VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__inv_2
XFILLER_0_178_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23641_ net572 top0.matmul0.matmul_stage_inst.d\[6\] top0.matmul0.matmul_stage_inst.c\[6\]
+ net558 VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__a22o_1
X_20853_ net229 net221 VGND VGND VPWR VPWR _12702_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23572_ top0.b_in_matmul\[9\] top0.matmul0.b\[9\] _02948_ VGND VGND VPWR VPWR _02953_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26360_ spi0.data_packed\[78\] spi0.data_packed\[79\] net690 VGND VGND VPWR VPWR
+ _05412_ sky130_fd_sc_hd__mux2_1
X_20784_ top0.cordic0.vec\[0\]\[2\] net285 net278 VGND VGND VPWR VPWR _12633_ sky130_fd_sc_hd__o21a_1
XFILLER_0_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25311_ _04656_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__inv_2
X_22523_ _02042_ _02078_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__nand2_2
XFILLER_0_135_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26291_ _05377_ VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25242_ _04517_ _04587_ _04475_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__a21oi_1
X_22454_ _01966_ _01969_ _02010_ VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_91_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21405_ _00942_ _12696_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__and2b_1
X_25173_ _04518_ _04520_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__nor2_4
X_22385_ _01942_ _01943_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24124_ _03480_ _03481_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__and2_1
XFILLER_0_161_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21336_ net213 _12705_ _13177_ net222 VGND VGND VPWR VPWR _13178_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24055_ _03372_ _03374_ _03375_ VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__nand3_2
XFILLER_0_124_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21267_ _13049_ _13109_ VGND VGND VPWR VPWR _13110_ sky130_fd_sc_hd__nand2_2
XFILLER_0_103_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23006_ top0.svm0.delta\[12\] _02510_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__xnor2_1
X_20218_ net264 _12066_ VGND VGND VPWR VPWR _12067_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_25_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21198_ net213 _12697_ _13041_ VGND VGND VPWR VPWR _13042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_198_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20149_ _11433_ top0.cordic0.in_valid VGND VGND VPWR VPWR _12003_ sky130_fd_sc_hd__nand2_4
X_24957_ _04226_ _04231_ _04216_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__o21a_1
X_14710_ _06873_ _06911_ _06912_ VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__a21oi_2
X_23908_ _03233_ _03265_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__xnor2_4
X_15690_ _07671_ _07675_ VGND VGND VPWR VPWR _07788_ sky130_fd_sc_hd__nor2_1
X_24888_ _04237_ _04239_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__xnor2_1
X_14641_ _06837_ _06845_ VGND VGND VPWR VPWR _06846_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_197_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26627_ clknet_leaf_25_clk_sys _00244_ net628 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_23839_ net566 net560 top0.matmul0.matmul_stage_inst.e\[13\] VGND VGND VPWR VPWR
+ _03197_ sky130_fd_sc_hd__o21a_2
XFILLER_0_200_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17360_ net418 net340 VGND VGND VPWR VPWR _09347_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14572_ _05822_ _06640_ VGND VGND VPWR VPWR _06778_ sky130_fd_sc_hd__nor2_1
X_26558_ clknet_leaf_52_clk_sys _00181_ net670 VGND VGND VPWR VPWR top0.pid_q.curr_error\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16311_ _07800_ _08401_ VGND VGND VPWR VPWR _08402_ sky130_fd_sc_hd__and2_1
X_25509_ _04840_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__clkbuf_1
X_13523_ _05735_ _05629_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17291_ _09286_ _09282_ top0.matmul0.matmul_stage_inst.mult1\[6\] VGND VGND VPWR
+ VPWR _09287_ sky130_fd_sc_hd__a21bo_1
X_26489_ clknet_leaf_61_clk_sys _00009_ net651 VGND VGND VPWR VPWR top0.pid_q.state\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_193_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19030_ net356 _11000_ _11001_ _11002_ net363 VGND VGND VPWR VPWR _11003_ sky130_fd_sc_hd__o2111a_2
X_16242_ _08305_ _08331_ VGND VGND VPWR VPWR _08333_ sky130_fd_sc_hd__nand2_1
X_13454_ net65 _05666_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13385_ _05578_ _05594_ _05597_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__o21a_1
X_16173_ _08263_ _08264_ VGND VGND VPWR VPWR _08265_ sky130_fd_sc_hd__xor2_1
XFILLER_0_112_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15124_ net517 net514 net494 net490 VGND VGND VPWR VPWR _07223_ sky130_fd_sc_hd__and4_1
XFILLER_0_51_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19932_ _11576_ _11427_ VGND VGND VPWR VPWR _11803_ sky130_fd_sc_hd__nor2_1
X_15055_ _07150_ _07151_ _07153_ VGND VGND VPWR VPWR _07154_ sky130_fd_sc_hd__a21bo_1
X_14006_ _06217_ _05501_ _05497_ _05686_ _06218_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__o32a_1
X_19863_ net229 VGND VGND VPWR VPWR _11739_ sky130_fd_sc_hd__clkinv_4
X_18814_ net373 VGND VGND VPWR VPWR _10790_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19794_ _11674_ _11448_ VGND VGND VPWR VPWR _11675_ sky130_fd_sc_hd__nand2_1
X_18745_ _10484_ _10721_ VGND VGND VPWR VPWR _10722_ sky130_fd_sc_hd__xor2_2
X_15957_ _08050_ _08051_ VGND VGND VPWR VPWR _08052_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14908_ _07074_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__clkbuf_1
X_18676_ _10652_ _10653_ VGND VGND VPWR VPWR _10654_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15888_ _07876_ _07878_ _07871_ VGND VGND VPWR VPWR _07984_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_53_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17627_ net1023 _09612_ VGND VGND VPWR VPWR _09614_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14839_ _06824_ _06955_ _06867_ VGND VGND VPWR VPWR _07037_ sky130_fd_sc_hd__a21o_1
XFILLER_0_188_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17558_ _09404_ _09392_ VGND VGND VPWR VPWR _09545_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16509_ _08492_ _08540_ _08493_ VGND VGND VPWR VPWR _08597_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_191_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17489_ net419 net330 net333 net422 VGND VGND VPWR VPWR _09476_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19228_ top0.pid_d.prev_error\[6\] top0.pid_d.curr_error\[6\] VGND VGND VPWR VPWR
+ _11176_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_86_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_86_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_144_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19159_ top0.kid\[14\] _11097_ _11099_ top0.kpd\[14\] VGND VGND VPWR VPWR _11115_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22170_ _01250_ _01731_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21121_ _12914_ _12919_ _12908_ VGND VGND VPWR VPWR _12966_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout303 net305 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__clkbuf_2
X_21052_ _12849_ _12857_ VGND VGND VPWR VPWR _12898_ sky130_fd_sc_hd__nand2_1
Xfanout314 net315 VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_4
Xfanout325 net326 VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_4
X_20003_ _11865_ _11869_ VGND VGND VPWR VPWR _11870_ sky130_fd_sc_hd__xnor2_1
Xfanout336 top0.pid_d.mult0.b\[6\] VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__clkbuf_4
Xfanout347 net348 VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__clkbuf_4
X_25860_ net888 _05029_ _05076_ _05080_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__a22o_1
Xfanout358 net359 VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__buf_2
Xfanout369 top0.pid_d.mult0.a\[14\] VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_94_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24811_ _04035_ _04032_ _04142_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__o21a_1
X_25791_ _12009_ net205 VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__nand2_1
XFILLER_0_158_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24742_ _03106_ _03826_ _04014_ _04015_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__a31o_1
XFILLER_0_154_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21954_ _01267_ _01102_ _01515_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__or3b_1
XFILLER_0_90_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20905_ net271 _12095_ _12713_ VGND VGND VPWR VPWR _12753_ sky130_fd_sc_hd__o21ba_1
X_24673_ _04017_ _04026_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__xnor2_1
X_21885_ _01429_ _01446_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__and2b_1
XFILLER_0_90_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26412_ clknet_leaf_62_clk_sys _00053_ net646 VGND VGND VPWR VPWR top0.kpq\[1\] sky130_fd_sc_hd__dfrtp_1
X_23624_ _02981_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__buf_4
X_20836_ _12681_ _12684_ VGND VGND VPWR VPWR _12685_ sky130_fd_sc_hd__xor2_2
XFILLER_0_194_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26343_ _05403_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23555_ top0.b_in_matmul\[1\] top0.matmul0.b\[1\] _02937_ VGND VGND VPWR VPWR _02944_
+ sky130_fd_sc_hd__mux2_1
X_20767_ _11608_ _12611_ _12615_ net306 VGND VGND VPWR VPWR _12616_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_193_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22506_ net119 net104 _01643_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26274_ net975 spi0.data_packed\[36\] net688 VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__mux2_1
X_23486_ net996 top0.matmul0.sin\[12\] _02904_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__mux2_1
X_20698_ _12347_ _12309_ VGND VGND VPWR VPWR _12547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25225_ _04411_ _04571_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__nor2_4
X_22437_ _01885_ _01989_ _01993_ _01994_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_116_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25156_ _04496_ _04503_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__xnor2_2
X_22368_ _11444_ _01926_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24107_ _03463_ _03464_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__or2_1
X_21319_ _13121_ _13127_ _13160_ VGND VGND VPWR VPWR _13161_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25087_ _04354_ _04359_ _04435_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22299_ _01839_ _01858_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_130_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24038_ _03394_ _03395_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__xnor2_4
X_16860_ _08921_ _08908_ _08909_ _08923_ VGND VGND VPWR VPWR _08924_ sky130_fd_sc_hd__a31o_1
X_15811_ net477 net506 VGND VGND VPWR VPWR _07907_ sky130_fd_sc_hd__nand2_2
X_16791_ top0.kiq\[5\] _08863_ _08866_ VGND VGND VPWR VPWR _08869_ sky130_fd_sc_hd__and3_1
X_25989_ top0.matmul0.beta_pass\[7\] _05169_ _05191_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__a21o_1
X_18530_ top0.pid_d.out\[7\] _10509_ net14 VGND VGND VPWR VPWR _10510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15742_ net448 net536 VGND VGND VPWR VPWR _07839_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18461_ _10439_ _10440_ VGND VGND VPWR VPWR _10441_ sky130_fd_sc_hd__or2_1
X_15673_ net508 _07770_ VGND VGND VPWR VPWR _07771_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17412_ _09353_ net396 VGND VGND VPWR VPWR _09399_ sky130_fd_sc_hd__nor2_1
X_14624_ _06823_ _06828_ VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18392_ net1023 net386 VGND VGND VPWR VPWR _10373_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17343_ top0.matmul0.beta_pass\[14\] _09331_ net562 VGND VGND VPWR VPWR _09332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14555_ net33 _05626_ VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13506_ _05470_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__buf_6
XFILLER_0_126_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17274_ top0.matmul0.beta_pass\[4\] _09272_ net562 VGND VGND VPWR VPWR _09273_ sky130_fd_sc_hd__mux2_1
X_14486_ _06661_ _06692_ _06664_ VGND VGND VPWR VPWR _06693_ sky130_fd_sc_hd__a21oi_1
X_19013_ top0.pid_d.out\[13\] top0.pid_d.curr_int\[13\] VGND VGND VPWR VPWR _10987_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_181_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16225_ _08315_ _08251_ _08252_ VGND VGND VPWR VPWR _08317_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13437_ _05643_ _05636_ _05645_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16156_ _08245_ _08246_ VGND VGND VPWR VPWR _08248_ sky130_fd_sc_hd__or2_1
X_13368_ _05549_ _05550_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15107_ net517 net485 VGND VGND VPWR VPWR _07206_ sky130_fd_sc_hd__nand2_1
X_16087_ _08176_ _08178_ VGND VGND VPWR VPWR _08180_ sky130_fd_sc_hd__nor2_1
X_13299_ _05510_ _05511_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__xnor2_2
X_19915_ _11787_ VGND VGND VPWR VPWR _11788_ sky130_fd_sc_hd__buf_6
X_15038_ top0.pid_d.prev_int\[8\] _07140_ _07144_ top0.pid_d.curr_int\[8\] VGND VGND
+ VPWR VPWR _00125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19846_ _11435_ _11722_ VGND VGND VPWR VPWR _11724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16989_ _09042_ _05438_ _09041_ VGND VGND VPWR VPWR _09044_ sky130_fd_sc_hd__and3_1
X_19777_ net82 _11657_ _11658_ _11575_ VGND VGND VPWR VPWR _11659_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18728_ _10700_ _10703_ VGND VGND VPWR VPWR _10705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18659_ net320 net376 VGND VGND VPWR VPWR _10637_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21670_ _11444_ _01066_ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20621_ _12262_ _12429_ VGND VGND VPWR VPWR _12470_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_188_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23340_ net134 _02755_ _02780_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__or3_1
X_20552_ _12399_ _12400_ VGND VGND VPWR VPWR _12401_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23271_ _02707_ _02719_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__and2_1
X_20483_ _12257_ _12331_ VGND VGND VPWR VPWR _12332_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_131_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25010_ _04354_ _04359_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22222_ _01777_ _01781_ _01782_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22153_ net124 _01065_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21104_ _12802_ _12875_ _12944_ _12947_ _12949_ VGND VGND VPWR VPWR _12950_ sky130_fd_sc_hd__a311oi_2
X_26961_ clknet_leaf_31_clk_sys _00578_ net617 VGND VGND VPWR VPWR top0.matmul0.b\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_22084_ _01640_ _01645_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout100 net101 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout111 net112 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout122 net125 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_8
X_25912_ _05102_ _05126_ _05127_ _05110_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__a22o_1
X_21035_ _12808_ _12881_ _12879_ VGND VGND VPWR VPWR _12882_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout133 net134 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_8
Xfanout144 net145 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_2
XFILLER_0_195_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26892_ clknet_leaf_105_clk_sys _00509_ net577 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout155 net156 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__buf_2
Xfanout166 net167 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_2
Xfanout177 net178 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_4
X_25843_ net76 _05059_ _05063_ _05064_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__a31o_1
Xfanout188 top0.cordic0.gm0.iter\[2\] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_4
Xfanout199 net200 VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_199_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25774_ top0.matmul0.op_in\[1\] net70 _05460_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__mux2_1
X_22986_ top0.svm0.delta\[9\] _02493_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24725_ _04069_ _04077_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__xnor2_4
X_21937_ _01267_ net147 _01216_ _01498_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__o31a_1
XFILLER_0_167_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24656_ _03868_ _03877_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__or2_1
X_21868_ net145 net129 _01122_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23607_ _02970_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20819_ _12543_ _12667_ VGND VGND VPWR VPWR _12668_ sky130_fd_sc_hd__or2b_1
X_24587_ _03940_ _03941_ _03830_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_154_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21799_ _01102_ _01360_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__xnor2_2
X_14340_ _06386_ _06548_ _06470_ VGND VGND VPWR VPWR _06549_ sky130_fd_sc_hd__a21oi_1
X_26326_ spi0.data_packed\[61\] spi0.data_packed\[62\] net699 VGND VGND VPWR VPWR
+ _05395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23538_ top0.a_in_matmul\[9\] top0.matmul0.a\[9\] _02926_ VGND VGND VPWR VPWR _02935_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_146_Left_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14271_ _06417_ _06418_ _06479_ _06480_ VGND VGND VPWR VPWR _06481_ sky130_fd_sc_hd__a31oi_4
X_26257_ _05360_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__clkbuf_1
X_23469_ net727 top0.matmul0.sin\[4\] _05461_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__mux2_1
X_16010_ _08100_ _08103_ VGND VGND VPWR VPWR _08104_ sky130_fd_sc_hd__xnor2_2
X_25208_ _04483_ _04488_ _04554_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__o21ai_1
X_13222_ top0.pid_d.state\[3\] _05441_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__and2_1
X_26188_ spi0.data_packed\[11\] _05322_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25139_ _04485_ _04486_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17961_ _09941_ _09946_ VGND VGND VPWR VPWR _09947_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16912_ top0.matmul0.beta_pass\[7\] _05436_ VGND VGND VPWR VPWR _08972_ sky130_fd_sc_hd__nand2_1
X_19700_ net291 _11567_ VGND VGND VPWR VPWR _11586_ sky130_fd_sc_hd__nor2_1
X_17892_ _09861_ _09878_ VGND VGND VPWR VPWR _09879_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_155_Left_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16843_ top0.pid_q.prev_error\[1\] top0.pid_q.curr_error\[1\] VGND VGND VPWR VPWR
+ _08908_ sky130_fd_sc_hd__nand2_1
X_19631_ net306 _11519_ VGND VGND VPWR VPWR _11520_ sky130_fd_sc_hd__nand2_1
X_19562_ net188 _11448_ VGND VGND VPWR VPWR _11451_ sky130_fd_sc_hd__nor2_2
X_16774_ net547 _05442_ _08854_ VGND VGND VPWR VPWR _08857_ sky130_fd_sc_hd__and3_1
X_13986_ _06092_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__inv_2
XFILLER_0_189_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18513_ _10348_ _10361_ _10362_ VGND VGND VPWR VPWR _10493_ sky130_fd_sc_hd__o21ai_2
X_15725_ net492 net502 VGND VGND VPWR VPWR _07822_ sky130_fd_sc_hd__nand2_1
X_19493_ _11384_ _11385_ VGND VGND VPWR VPWR _11386_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18444_ top0.pid_d.out\[6\] _10424_ net14 VGND VGND VPWR VPWR _10425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15656_ net457 net529 VGND VGND VPWR VPWR _07754_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_199_Right_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14607_ _06792_ _06808_ _06811_ VGND VGND VPWR VPWR _06812_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18375_ net405 net310 VGND VGND VPWR VPWR _10356_ sky130_fd_sc_hd__nand2_1
X_15587_ _07543_ _07544_ _07685_ VGND VGND VPWR VPWR _07686_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_164_Left_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17326_ top0.matmul0.matmul_stage_inst.mult1\[11\] top0.matmul0.matmul_stage_inst.mult2\[11\]
+ VGND VGND VPWR VPWR _09317_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14538_ _06742_ _06744_ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_173_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17257_ top0.matmul0.matmul_stage_inst.mult2\[1\] top0.matmul0.matmul_stage_inst.mult1\[0\]
+ top0.matmul0.matmul_stage_inst.mult2\[0\] top0.matmul0.matmul_stage_inst.mult1\[1\]
+ VGND VGND VPWR VPWR _09258_ sky130_fd_sc_hd__a31o_1
X_14469_ _06556_ VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__clkinvlp_2
X_16208_ _08167_ _08172_ _08299_ VGND VGND VPWR VPWR _08300_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17188_ net554 _09197_ _09198_ _08994_ VGND VGND VPWR VPWR _09199_ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16139_ _08165_ _08230_ VGND VGND VPWR VPWR _08232_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_173_Left_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19829_ _11430_ _11707_ net175 VGND VGND VPWR VPWR _11708_ sky130_fd_sc_hd__o21a_1
XFILLER_0_194_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22840_ top0.svm0.counter\[9\] VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_196_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22771_ top0.pid_q.prev_int\[15\] _02291_ _02294_ net772 VGND VGND VPWR VPWR _00434_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24510_ _02998_ _03000_ _03093_ _03094_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__o22a_2
X_21722_ _01278_ _01279_ _01283_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25490_ top0.matmul0.matmul_stage_inst.mult1\[1\] _03756_ _04829_ VGND VGND VPWR
+ VPWR _04831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_182_Left_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_166_Right_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24441_ _03795_ _03796_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__and2_1
X_21653_ _01212_ _01214_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20604_ _12428_ _12452_ VGND VGND VPWR VPWR _12453_ sky130_fd_sc_hd__xnor2_2
X_27160_ clknet_leaf_90_clk_sys _00774_ net602 VGND VGND VPWR VPWR top0.a_in_matmul\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_24372_ _03725_ _03728_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__xnor2_2
X_21584_ _01142_ _01145_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_163_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26111_ _05275_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__clkbuf_4
X_20535_ _12377_ _12383_ VGND VGND VPWR VPWR _12384_ sky130_fd_sc_hd__xnor2_2
X_23323_ _02768_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27091_ clknet_leaf_22_clk_sys _00708_ net607 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26042_ _05013_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__buf_2
X_20466_ _12296_ _12297_ _12295_ VGND VGND VPWR VPWR _12315_ sky130_fd_sc_hd__o21ba_1
X_23254_ net161 _11511_ _02679_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__and3_1
XFILLER_0_162_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22205_ net124 net126 net144 VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__and3b_1
X_23185_ _02646_ _06546_ _02649_ net837 VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__a22o_1
X_20397_ net262 net252 VGND VGND VPWR VPWR _12246_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_191_Left_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22136_ _01205_ _01696_ _01697_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_100_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22067_ _01619_ _01628_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__xor2_2
X_26944_ clknet_leaf_6_clk_sys _00561_ net594 VGND VGND VPWR VPWR top0.matmul0.a\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_21018_ _12835_ _12864_ VGND VGND VPWR VPWR _12865_ sky130_fd_sc_hd__xnor2_4
X_26875_ clknet_leaf_40_clk_sys _00492_ net682 VGND VGND VPWR VPWR top0.svm0.tB\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25826_ _05043_ _05044_ _05047_ _05046_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__a31o_1
X_13840_ _06051_ _06052_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13771_ _05970_ _05981_ _05983_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__a21o_1
X_25757_ _04999_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22969_ _02478_ _02474_ _02324_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__a21o_1
XFILLER_0_168_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15510_ _07607_ _07608_ _07220_ VGND VGND VPWR VPWR _07609_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24708_ _03963_ _04061_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__xnor2_1
X_16490_ _08569_ _08577_ VGND VGND VPWR VPWR _08578_ sky130_fd_sc_hd__xor2_1
X_25688_ top0.matmul0.sin\[13\] _04954_ _04886_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15441_ net489 net484 net511 VGND VGND VPWR VPWR _07540_ sky130_fd_sc_hd__and3_1
X_24639_ _03991_ _03992_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__nand2_2
XFILLER_0_33_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18160_ _10137_ _10143_ VGND VGND VPWR VPWR _10144_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15372_ _07436_ _07437_ _07470_ VGND VGND VPWR VPWR _07471_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17111_ top0.pid_q.curr_error\[14\] _08860_ _09116_ VGND VGND VPWR VPWR _09132_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14323_ net56 _06268_ _06455_ VGND VGND VPWR VPWR _06533_ sky130_fd_sc_hd__nand3_1
X_26309_ _05386_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18091_ net365 _10074_ VGND VGND VPWR VPWR _10075_ sky130_fd_sc_hd__nand2_2
XFILLER_0_68_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27289_ clknet_3_3__leaf_clk_mosi _00903_ VGND VGND VPWR VPWR spi0.data_packed\[75\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17042_ net551 _09093_ VGND VGND VPWR VPWR _09094_ sky130_fd_sc_hd__and2_1
X_14254_ _06191_ _06193_ _06350_ net60 VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13205_ _05431_ top0.matmul0.state\[1\] net748 VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14185_ net41 _05611_ _05612_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18993_ net309 _10966_ _10964_ VGND VGND VPWR VPWR _10967_ sky130_fd_sc_hd__a21oi_1
X_17944_ _09918_ _09929_ VGND VGND VPWR VPWR _09930_ sky130_fd_sc_hd__xor2_1
XFILLER_0_178_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17875_ net420 net319 VGND VGND VPWR VPWR _09862_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19614_ _11473_ _11501_ _11502_ _11472_ _11476_ VGND VGND VPWR VPWR _11503_ sky130_fd_sc_hd__o221a_1
X_16826_ top0.matmul0.beta_pass\[1\] _08891_ VGND VGND VPWR VPWR _08892_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16757_ _08788_ _08839_ VGND VGND VPWR VPWR _08841_ sky130_fd_sc_hd__and2_1
X_19545_ _11434_ VGND VGND VPWR VPWR _11435_ sky130_fd_sc_hd__clkbuf_4
X_13969_ net48 _05605_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__nand2_1
XFILLER_0_177_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15708_ top0.pid_q.curr_int\[2\] _07804_ VGND VGND VPWR VPWR _07805_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16688_ net452 net455 net498 _08772_ VGND VGND VPWR VPWR _08773_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19476_ _11368_ _11369_ VGND VGND VPWR VPWR _11371_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_185_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18427_ _10406_ _10407_ VGND VGND VPWR VPWR _10408_ sky130_fd_sc_hd__xor2_1
X_15639_ _07734_ _07736_ VGND VGND VPWR VPWR _07737_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18358_ _10337_ _10246_ _10338_ VGND VGND VPWR VPWR _10339_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17309_ top0.matmul0.beta_pass\[9\] _09302_ net562 VGND VGND VPWR VPWR _09303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18289_ net338 net373 VGND VGND VPWR VPWR _10271_ sky130_fd_sc_hd__nand2_1
X_20320_ _12161_ _12168_ VGND VGND VPWR VPWR _12169_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20251_ net301 net276 VGND VGND VPWR VPWR _12100_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_102_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20182_ _12031_ VGND VGND VPWR VPWR _12032_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24990_ _04252_ _04338_ _04339_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__a21oi_1
X_23941_ _03229_ _03230_ _03298_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__a21oi_2
X_26660_ clknet_leaf_77_clk_sys _00277_ net635 VGND VGND VPWR VPWR top0.pid_d.mult0.a\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_23872_ _03227_ _03228_ _03131_ _03137_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__a211o_1
X_25611_ net739 _04896_ _04891_ _04897_ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__o22a_1
X_22823_ top0.svm0.tA\[10\] net169 VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__or2b_1
XFILLER_0_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26591_ clknet_leaf_65_clk_sys _00214_ net657 VGND VGND VPWR VPWR top0.pid_q.curr_int\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_25542_ net951 top0.matmul0.matmul_stage_inst.f\[10\] _04856_ VGND VGND VPWR VPWR
+ _04858_ sky130_fd_sc_hd__mux2_1
X_22754_ _02293_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__buf_2
XFILLER_0_17_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21705_ _01266_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__clkbuf_4
X_25473_ _04717_ _04815_ _04814_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22685_ _02138_ _02171_ _02173_ _02209_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__o211a_1
X_27212_ clknet_leaf_6_clk_sys _00826_ net598 VGND VGND VPWR VPWR top0.cordic0.slte0.opB\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_24424_ _03777_ _03779_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__xor2_1
XFILLER_0_136_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21636_ net138 _01101_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27143_ clknet_leaf_31_clk_sys _00757_ net619 VGND VGND VPWR VPWR top0.b_in_matmul\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_191_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24355_ _03710_ _03711_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__xor2_1
XFILLER_0_105_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21567_ _01110_ _01128_ VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__xor2_1
X_23306_ _11448_ _02751_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__or2_1
X_27074_ clknet_leaf_21_clk_sys _00691_ net607 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.c\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20518_ _12279_ _12366_ VGND VGND VPWR VPWR _12367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24286_ _03643_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21498_ net863 _12034_ _12037_ VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__nand3_1
XFILLER_0_132_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26025_ top0.matmul0.beta_pass\[15\] _05203_ _05219_ VGND VGND VPWR VPWR _05220_
+ sky130_fd_sc_hd__a21o_1
X_20449_ _12296_ _12297_ VGND VGND VPWR VPWR _12298_ sky130_fd_sc_hd__xnor2_1
X_23237_ net233 net228 net223 net220 net203 net196 VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__mux4_2
XFILLER_0_63_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23168_ _02641_ _06748_ _02645_ net780 VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22119_ _01640_ _01660_ _01645_ _01653_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__a211o_1
X_23099_ top0.svm0.delta\[1\] _02597_ _02599_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__a21o_1
X_15990_ top0.pid_q.out\[5\] top0.pid_q.curr_int\[5\] VGND VGND VPWR VPWR _08084_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14941_ spi0.data_packed\[45\] top0.kid\[13\] _07086_ VGND VGND VPWR VPWR _07092_
+ sky130_fd_sc_hd__mux2_1
X_26927_ clknet_leaf_7_clk_sys _00544_ net593 VGND VGND VPWR VPWR top0.matmul0.cos\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_202_Right_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17660_ _09641_ _09646_ VGND VGND VPWR VPWR _09647_ sky130_fd_sc_hd__xnor2_1
X_26858_ clknet_leaf_40_clk_sys _00475_ net678 VGND VGND VPWR VPWR top0.svm0.tA\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14872_ spi0.data_packed\[76\] top0.kpd\[12\] _07053_ VGND VGND VPWR VPWR _07056_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16611_ net498 _08696_ VGND VGND VPWR VPWR _08697_ sky130_fd_sc_hd__nand2_1
X_25809_ _05033_ _05034_ _05035_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__a21oi_1
X_13823_ _06024_ _06026_ _06035_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__or3_1
XFILLER_0_187_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17591_ net347 _09524_ net340 VGND VGND VPWR VPWR _09578_ sky130_fd_sc_hd__and3b_1
XFILLER_0_173_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26789_ clknet_leaf_3_clk_sys _00406_ net583 VGND VGND VPWR VPWR top0.cordic0.sin\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_187_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16542_ _08567_ _08577_ _08628_ VGND VGND VPWR VPWR _08629_ sky130_fd_sc_hd__a21o_1
X_19330_ top0.matmul0.alpha_pass\[15\] _11262_ VGND VGND VPWR VPWR _11269_ sky130_fd_sc_hd__xnor2_1
X_13754_ _05965_ _05966_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__or2b_1
XFILLER_0_85_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19261_ top0.pid_d.prev_error\[9\] top0.pid_d.curr_error\[9\] VGND VGND VPWR VPWR
+ _11206_ sky130_fd_sc_hd__xnor2_1
X_16473_ net516 top0.pid_q.mult0.b\[15\] VGND VGND VPWR VPWR _08561_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_155_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13685_ _05889_ _05892_ _05897_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__o21a_1
X_18212_ _10192_ _10194_ VGND VGND VPWR VPWR _10195_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15424_ _07392_ _07396_ VGND VGND VPWR VPWR _07523_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19192_ _11125_ _11139_ _11142_ _11143_ _07800_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__o311a_1
XFILLER_0_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18143_ _10112_ _10126_ VGND VGND VPWR VPWR _10127_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15355_ _07432_ _07453_ VGND VGND VPWR VPWR _07454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_198_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14306_ _06514_ _06515_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_202_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18074_ _09972_ _09974_ _09902_ VGND VGND VPWR VPWR _10059_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15286_ net525 _07366_ VGND VGND VPWR VPWR _07385_ sky130_fd_sc_hd__nand2_1
Xhold208 top0.svm0.tA\[14\] VGND VGND VPWR VPWR net908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17025_ top0.pid_q.state\[3\] _09070_ _09077_ net551 _08881_ VGND VGND VPWR VPWR
+ _09078_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold219 top0.currT_r\[1\] VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ _06419_ _06420_ _06446_ _06447_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14168_ _06370_ _06379_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14099_ _06222_ _06224_ VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__or2_1
X_18976_ _10944_ _10949_ VGND VGND VPWR VPWR _10950_ sky130_fd_sc_hd__xnor2_2
X_17927_ _09911_ _09912_ VGND VGND VPWR VPWR _09913_ sky130_fd_sc_hd__xnor2_1
X_17858_ net346 net383 VGND VGND VPWR VPWR _09845_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_0__f_clk_sys clknet_0_clk_sys VGND VGND VPWR VPWR clknet_3_0__leaf_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_178_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16809_ top0.kiq\[14\] _05448_ _08854_ VGND VGND VPWR VPWR _08878_ sky130_fd_sc_hd__and3_1
X_17789_ net399 net339 VGND VGND VPWR VPWR _09776_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19528_ net165 net160 net157 top0.cordic0.vec\[1\]\[3\] net197 net191 VGND VGND VPWR
+ VPWR _11418_ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19459_ net431 _10679_ _11355_ net441 _11209_ VGND VGND VPWR VPWR _11356_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22470_ net85 _02025_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21421_ _00984_ _00986_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24140_ _03495_ _03497_ VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__nand2_1
X_21352_ _00917_ _00920_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20303_ _12150_ _12151_ VGND VGND VPWR VPWR _12152_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24071_ _03426_ _03374_ _03371_ _03424_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__o211a_1
X_21283_ _13124_ _13125_ VGND VGND VPWR VPWR _13126_ sky130_fd_sc_hd__xor2_1
Xfanout2 _11548_ VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__buf_4
XFILLER_0_97_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23022_ net168 _02483_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__nor2_1
X_20234_ _12078_ _12082_ VGND VGND VPWR VPWR _12083_ sky130_fd_sc_hd__xnor2_2
X_20165_ net205 _05425_ VGND VGND VPWR VPWR _12017_ sky130_fd_sc_hd__or2_2
XFILLER_0_200_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24973_ _04237_ _04239_ _04323_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__a21oi_1
X_20096_ _11953_ _11955_ top0.cordic0.slte0.opA\[12\] VGND VGND VPWR VPWR _11956_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26712_ clknet_leaf_72_clk_sys _00329_ net655 VGND VGND VPWR VPWR top0.pid_d.curr_int\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_157_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23924_ _03279_ _03281_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26643_ clknet_leaf_78_clk_sys _00260_ net632 VGND VGND VPWR VPWR top0.pid_d.out\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23855_ _03209_ _03212_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_169_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22806_ _02324_ top0.svm0.tA\[6\] VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__and2_1
X_26574_ clknet_leaf_52_clk_sys _00197_ net670 VGND VGND VPWR VPWR top0.pid_q.prev_error\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23786_ _03047_ _02982_ _03142_ _03143_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__o31ai_2
X_20998_ net277 net259 net255 VGND VGND VPWR VPWR _12845_ sky130_fd_sc_hd__or3b_1
XFILLER_0_196_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25525_ top0.matmul0.b\[2\] top0.matmul0.matmul_stage_inst.f\[2\] _04846_ VGND VGND
+ VPWR VPWR _04849_ sky130_fd_sc_hd__mux2_1
X_22737_ top0.state\[1\] net206 top0.start_svm _02283_ VGND VGND VPWR VPWR _00412_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_137_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25456_ _04733_ _04797_ _04798_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13470_ _05682_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22668_ _02197_ _02196_ _02192_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24407_ _03759_ _03762_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_152_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21619_ _01150_ _01152_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_192_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25387_ _04728_ _04730_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22599_ net114 _02149_ _02152_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27126_ clknet_3_6__leaf_clk_sys _00740_ net665 VGND VGND VPWR VPWR top0.c_out_calc\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_129_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15140_ _07236_ _07238_ VGND VGND VPWR VPWR _07239_ sky130_fd_sc_hd__and2b_1
X_24338_ _03184_ _03190_ _03181_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27057_ clknet_leaf_20_clk_sys _00674_ net609 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.d\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15071_ top0.pid_q.mult0.a\[2\] net471 VGND VGND VPWR VPWR _07170_ sky130_fd_sc_hd__nand2_2
X_24269_ _03623_ _03626_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__or2b_1
XFILLER_0_22_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14022_ _06111_ _06116_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__nand2_1
X_26008_ top0.pid_q.out\[11\] _05198_ _05199_ spi0.data_packed\[59\] VGND VGND VPWR
+ VPWR _05207_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18830_ _10804_ _10805_ VGND VGND VPWR VPWR _10806_ sky130_fd_sc_hd__nand2_1
XFILLER_0_175_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18761_ net390 _10734_ _10735_ _10737_ VGND VGND VPWR VPWR _10738_ sky130_fd_sc_hd__o31ai_4
X_15973_ _08063_ _08067_ VGND VGND VPWR VPWR _08068_ sky130_fd_sc_hd__xnor2_1
X_17712_ _09696_ _09698_ VGND VGND VPWR VPWR _09699_ sky130_fd_sc_hd__xnor2_2
X_14924_ spi0.data_packed\[37\] top0.kid\[5\] _07075_ VGND VGND VPWR VPWR _07083_
+ sky130_fd_sc_hd__mux2_1
X_18692_ _10655_ _10669_ VGND VGND VPWR VPWR _10670_ sky130_fd_sc_hd__xnor2_2
Xhold80 top0.svm0.tA\[6\] VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 top0.matmul0.matmul_stage_inst.c\[8\] VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17643_ _09483_ _09628_ _09629_ VGND VGND VPWR VPWR _09630_ sky130_fd_sc_hd__o21a_1
X_14855_ spi0.data_packed\[68\] top0.kpd\[4\] _07042_ VGND VGND VPWR VPWR _07047_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13806_ _05981_ _06018_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__xnor2_1
X_17574_ net410 net352 VGND VGND VPWR VPWR _09561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14786_ _06986_ _06983_ _06952_ VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19313_ net313 _11117_ _11253_ _10067_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16525_ top0.pid_q.out\[10\] top0.pid_q.curr_int\[10\] VGND VGND VPWR VPWR _08613_
+ sky130_fd_sc_hd__or2_1
X_13737_ _05881_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16456_ _08467_ _08469_ _08544_ _08386_ VGND VGND VPWR VPWR _08545_ sky130_fd_sc_hd__o2bb2a_1
X_19244_ top0.matmul0.alpha_pass\[7\] _11180_ VGND VGND VPWR VPWR _11191_ sky130_fd_sc_hd__nand2_1
X_13668_ _05879_ _05880_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15407_ net481 _07459_ VGND VGND VPWR VPWR _07506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19175_ top0.pid_d.prev_error\[0\] top0.pid_d.curr_error\[0\] _11126_ VGND VGND VPWR
+ VPWR _11128_ sky130_fd_sc_hd__a21oi_1
X_16387_ _08334_ _08475_ _08476_ VGND VGND VPWR VPWR _08477_ sky130_fd_sc_hd__a21oi_2
X_13599_ _05735_ _05531_ _05532_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__or3_2
XFILLER_0_14_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18126_ _10106_ _10109_ VGND VGND VPWR VPWR _10110_ sky130_fd_sc_hd__xnor2_2
X_15338_ net531 net491 VGND VGND VPWR VPWR _07437_ sky130_fd_sc_hd__nand2_2
X_18057_ _09951_ _09954_ _10041_ VGND VGND VPWR VPWR _10042_ sky130_fd_sc_hd__o21ai_1
X_15269_ net479 _07323_ _07367_ _07322_ VGND VGND VPWR VPWR _07368_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17008_ _09059_ _09061_ VGND VGND VPWR VPWR _09062_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire9 _02593_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
Xfanout507 top0.pid_q.mult0.a\[12\] VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__buf_2
XFILLER_0_111_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout518 net1028 VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__buf_2
XFILLER_0_10_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout529 net530 VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__clkbuf_2
X_18959_ _10875_ _10931_ _10932_ VGND VGND VPWR VPWR _10933_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_82_clk_sys clknet_3_4__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_82_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_21970_ _01523_ _01527_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__or2_1
X_20921_ net223 net218 VGND VGND VPWR VPWR _12769_ sky130_fd_sc_hd__and2b_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23640_ _02997_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__clkbuf_4
X_20852_ _12698_ _12700_ VGND VGND VPWR VPWR _12701_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_194_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_190_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23571_ _02952_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20783_ _11408_ _12631_ VGND VGND VPWR VPWR _12632_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25310_ _04610_ _04654_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22522_ _02038_ _02040_ _02036_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26290_ net942 net925 net690 VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25241_ _04517_ _04587_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22453_ _01966_ _01969_ _01962_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_106_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21404_ net232 _12696_ _12761_ _00942_ _00970_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__a221o_1
X_25172_ _04069_ _04412_ _04519_ _03765_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__o22a_1
X_22384_ _01898_ _01941_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__nand2_1
XFILLER_0_199_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24123_ _03479_ _03408_ _03400_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__o21ai_1
X_21335_ net242 net236 _11759_ _12697_ VGND VGND VPWR VPWR _13177_ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24054_ _03404_ _03405_ _03410_ _03411_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__o211a_1
X_21266_ _13044_ _13051_ VGND VGND VPWR VPWR _13109_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23005_ _02508_ _02504_ _02509_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20217_ net279 net269 VGND VGND VPWR VPWR _12066_ sky130_fd_sc_hd__and2b_2
X_21197_ _12180_ _12990_ VGND VGND VPWR VPWR _13041_ sky130_fd_sc_hd__nor2_1
XFILLER_0_198_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20148_ _11999_ _12000_ _12001_ _12002_ top0.cordic0.slte0.opA\[17\] VGND VGND VPWR
+ VPWR _00377_ sky130_fd_sc_hd__a32o_1
XFILLER_0_99_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24956_ _04071_ _04076_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__nor2_1
X_20079_ _11937_ _11939_ VGND VGND VPWR VPWR _11940_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23907_ _03247_ _03260_ _03263_ _03264_ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__o22a_2
XFILLER_0_99_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24887_ _04130_ _04135_ _04238_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__o21a_1
X_14640_ _06839_ _06844_ VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__xor2_1
X_26626_ clknet_leaf_25_clk_sys _00243_ net627 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[14\]
+ sky130_fd_sc_hd__dfrtp_2
X_23838_ net570 net575 top0.matmul0.matmul_stage_inst.f\[13\] VGND VGND VPWR VPWR
+ _03196_ sky130_fd_sc_hd__o21a_2
XFILLER_0_185_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14571_ _06323_ VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__inv_2
X_26557_ clknet_leaf_49_clk_sys _00180_ net687 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_23769_ _03078_ _03079_ _03080_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__o21a_1
X_16310_ top0.pid_q.out\[8\] _08400_ _07700_ VGND VGND VPWR VPWR _08401_ sky130_fd_sc_hd__mux2_1
X_25508_ top0.matmul0.matmul_stage_inst.mult1\[10\] _04535_ _03148_ VGND VGND VPWR
+ VPWR _04840_ sky130_fd_sc_hd__mux2_1
X_13522_ net57 VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__inv_2
X_17290_ top0.matmul0.matmul_stage_inst.mult2\[6\] VGND VGND VPWR VPWR _09286_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26488_ clknet_leaf_55_clk_sys _00008_ net667 VGND VGND VPWR VPWR top0.pid_q.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16241_ _08305_ _08331_ VGND VGND VPWR VPWR _08332_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13453_ _05665_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__buf_4
X_25439_ _04190_ _04097_ _04781_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16172_ net453 net516 VGND VGND VPWR VPWR _08264_ sky130_fd_sc_hd__nand2_1
X_13384_ _05578_ _05594_ _05596_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15123_ _07161_ _07175_ VGND VGND VPWR VPWR _07222_ sky130_fd_sc_hd__nor2_2
X_27109_ clknet_leaf_89_clk_sys _00015_ net603 VGND VGND VPWR VPWR top0.matmul0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_181_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19931_ top0.cordic0.slte0.opA\[0\] _11799_ VGND VGND VPWR VPWR _11802_ sky130_fd_sc_hd__and2_1
X_15054_ _07150_ _07151_ _07152_ VGND VGND VPWR VPWR _07153_ sky130_fd_sc_hd__o21ai_1
X_14005_ net1030 _06211_ _06212_ _05894_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__o22a_1
XFILLER_0_142_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19862_ net175 _11727_ _11737_ _11738_ VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18813_ _10718_ _10716_ _10723_ _10788_ VGND VGND VPWR VPWR _10789_ sky130_fd_sc_hd__a31o_1
X_19793_ _11444_ VGND VGND VPWR VPWR _11674_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18744_ net362 _10720_ VGND VGND VPWR VPWR _10721_ sky130_fd_sc_hd__nand2_1
X_15956_ _08047_ _08049_ VGND VGND VPWR VPWR _08051_ sky130_fd_sc_hd__nand2_1
X_14907_ spi0.data_packed\[61\] top0.kpq\[13\] _07064_ VGND VGND VPWR VPWR _07074_
+ sky130_fd_sc_hd__mux2_1
X_18675_ _10649_ _10651_ VGND VGND VPWR VPWR _10653_ sky130_fd_sc_hd__nand2_1
X_15887_ _07867_ _07981_ _07982_ VGND VGND VPWR VPWR _07983_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17626_ net1022 _09609_ _09612_ VGND VGND VPWR VPWR _09613_ sky130_fd_sc_hd__o21a_1
X_14838_ _07013_ _07014_ net26 _06867_ VGND VGND VPWR VPWR _07036_ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14769_ _06947_ _06970_ VGND VGND VPWR VPWR _06971_ sky130_fd_sc_hd__xnor2_2
X_17557_ _09537_ _09539_ _09543_ VGND VGND VPWR VPWR _09544_ sky130_fd_sc_hd__o21a_1
XFILLER_0_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16508_ _08592_ _08595_ VGND VGND VPWR VPWR _08596_ sky130_fd_sc_hd__xnor2_1
X_17488_ _09414_ _09473_ _09474_ VGND VGND VPWR VPWR _09475_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19227_ _11173_ _11166_ _11174_ VGND VGND VPWR VPWR _11175_ sky130_fd_sc_hd__a21o_1
XFILLER_0_171_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16439_ _08525_ _08527_ VGND VGND VPWR VPWR _08528_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_29_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_29_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19158_ net372 _11095_ _11114_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18109_ _10090_ _10091_ VGND VGND VPWR VPWR _10093_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19089_ net371 _11054_ _11055_ _11060_ VGND VGND VPWR VPWR _11061_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21120_ _12897_ _12933_ _12964_ VGND VGND VPWR VPWR _12965_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_41_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21051_ _11789_ _12896_ VGND VGND VPWR VPWR _12897_ sky130_fd_sc_hd__or2_1
Xfanout304 net305 VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout315 top0.pid_d.mult0.b\[12\] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20002_ _11867_ _11868_ VGND VGND VPWR VPWR _11869_ sky130_fd_sc_hd__nand2_1
Xfanout326 top0.pid_d.mult0.b\[9\] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__buf_2
Xfanout337 net339 VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__clkbuf_4
Xfanout348 net350 VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__clkbuf_4
Xfanout359 net360 VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__clkbuf_4
X_24810_ _04141_ _04143_ VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25790_ _12009_ _05019_ _05020_ top0.cordic0.in_valid VGND VGND VPWR VPWR _00728_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24741_ _04090_ _04093_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__xnor2_2
X_21953_ net156 net130 VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20904_ _12717_ _12750_ _12751_ VGND VGND VPWR VPWR _12752_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_167_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24672_ _04020_ _04025_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__xnor2_1
X_21884_ _01432_ _01435_ _01445_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26411_ clknet_leaf_62_clk_sys _00052_ net650 VGND VGND VPWR VPWR top0.kpq\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23623_ _02979_ _02980_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20835_ _12682_ _12683_ VGND VGND VPWR VPWR _12684_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_59_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_182_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26342_ spi0.data_packed\[69\] spi0.data_packed\[70\] net689 VGND VGND VPWR VPWR
+ _05403_ sky130_fd_sc_hd__mux2_1
X_23554_ _02943_ VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20766_ _12612_ _12613_ _12614_ VGND VGND VPWR VPWR _12615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22505_ _01069_ _01924_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__xor2_4
X_26273_ net945 VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23485_ _02907_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__clkbuf_1
X_20697_ _12544_ _12545_ VGND VGND VPWR VPWR _12546_ sky130_fd_sc_hd__nor2_2
XFILLER_0_190_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25224_ _04069_ _04339_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__and2_2
XFILLER_0_73_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22436_ _01896_ _01943_ _01988_ net210 VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__a211o_1
XFILLER_0_165_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25155_ _04501_ _04502_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__or2b_1
XFILLER_0_32_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22367_ _01924_ _01925_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24106_ _02978_ _03195_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__nor2_2
X_21318_ _13121_ _13127_ _13132_ VGND VGND VPWR VPWR _13160_ sky130_fd_sc_hd__o21ba_1
X_25086_ _04354_ _04359_ _04352_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22298_ _01856_ _01857_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_68_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24037_ _03354_ _03356_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__xnor2_2
X_21249_ _12535_ _12539_ VGND VGND VPWR VPWR _13093_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15810_ net469 net512 VGND VGND VPWR VPWR _07906_ sky130_fd_sc_hd__nand2_2
X_16790_ net1026 _08856_ _08859_ net751 _08868_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__a221o_1
X_25988_ top0.pid_q.out\[7\] _12032_ _05014_ spi0.data_packed\[55\] VGND VGND VPWR
+ VPWR _05191_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15741_ net538 net446 VGND VGND VPWR VPWR _07838_ sky130_fd_sc_hd__nand2_2
X_24939_ _03112_ _03280_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__nor2_1
XFILLER_0_198_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18460_ _10436_ _10438_ VGND VGND VPWR VPWR _10440_ sky130_fd_sc_hd__and2_1
X_15672_ net511 _07769_ VGND VGND VPWR VPWR _07770_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_77_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14623_ _06826_ _06827_ VGND VGND VPWR VPWR _06828_ sky130_fd_sc_hd__xnor2_1
X_17411_ net400 _09395_ _09397_ net405 VGND VGND VPWR VPWR _09398_ sky130_fd_sc_hd__a22o_1
X_18391_ net1022 net378 VGND VGND VPWR VPWR _10372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26609_ clknet_leaf_86_clk_sys _00004_ net641 VGND VGND VPWR VPWR top0.pid_d.state\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_96_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17342_ _09329_ _09330_ VGND VGND VPWR VPWR _09331_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_157_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_200_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14554_ net30 _05605_ VGND VGND VPWR VPWR _06760_ sky130_fd_sc_hd__nand2_2
XFILLER_0_82_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13505_ top0.matmul0.alpha_pass\[14\] _05436_ _05717_ VGND VGND VPWR VPWR _05718_
+ sky130_fd_sc_hd__and3_1
X_17273_ _09270_ _09271_ VGND VGND VPWR VPWR _09272_ sky130_fd_sc_hd__xnor2_1
X_14485_ _06560_ _06663_ _06665_ VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_30_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_30_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16224_ _08251_ _08252_ _08315_ VGND VGND VPWR VPWR _08316_ sky130_fd_sc_hd__a21o_1
X_19012_ _10911_ _10915_ _10910_ VGND VGND VPWR VPWR _10986_ sky130_fd_sc_hd__a21o_1
XFILLER_0_180_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13436_ _05559_ _05598_ _05648_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_130_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16155_ _08245_ _08246_ VGND VGND VPWR VPWR _08247_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13367_ net57 _05579_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15106_ net514 net490 VGND VGND VPWR VPWR _07205_ sky130_fd_sc_hd__nand2_1
X_16086_ _08176_ _08178_ VGND VGND VPWR VPWR _08179_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13298_ _05487_ _05492_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__xor2_1
XFILLER_0_107_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19914_ net214 VGND VGND VPWR VPWR _11787_ sky130_fd_sc_hd__inv_2
X_15037_ top0.pid_d.prev_int\[7\] _07140_ _07144_ net911 VGND VGND VPWR VPWR _00124_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19845_ _11430_ _11722_ net175 VGND VGND VPWR VPWR _11723_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19776_ net181 _11657_ VGND VGND VPWR VPWR _11658_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16988_ _05438_ _09041_ _09042_ VGND VGND VPWR VPWR _09043_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18727_ _10700_ _10703_ VGND VGND VPWR VPWR _10704_ sky130_fd_sc_hd__nor2_1
X_15939_ _07948_ _07950_ _07949_ VGND VGND VPWR VPWR _08034_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18658_ net327 net368 VGND VGND VPWR VPWR _10636_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_171_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17609_ _09562_ _09595_ VGND VGND VPWR VPWR _09596_ sky130_fd_sc_hd__xnor2_1
X_18589_ _10566_ _10567_ VGND VGND VPWR VPWR _10568_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20620_ net282 _12466_ _12467_ _11525_ _12468_ VGND VGND VPWR VPWR _12469_ sky130_fd_sc_hd__a221o_2
XFILLER_0_175_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20551_ _12377_ _12381_ _12382_ VGND VGND VPWR VPWR _12400_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_188_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23270_ _02717_ _02718_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20482_ _12251_ _12249_ VGND VGND VPWR VPWR _12331_ sky130_fd_sc_hd__xor2_1
XFILLER_0_54_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22221_ _01716_ _01780_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22152_ _01213_ net99 _01223_ _01712_ _01713_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__a311o_1
X_21103_ _12945_ _12948_ _12875_ VGND VGND VPWR VPWR _12949_ sky130_fd_sc_hd__o21a_1
XFILLER_0_160_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26960_ clknet_leaf_14_clk_sys _00577_ net617 VGND VGND VPWR VPWR top0.matmul0.b\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22083_ _01616_ _01642_ _01644_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__a21oi_2
Xfanout101 net102 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
Xfanout112 net113 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_196_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_195_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25911_ net429 _05114_ _05115_ top0.matmul0.alpha_pass\[10\] VGND VGND VPWR VPWR
+ _05127_ sky130_fd_sc_hd__a22oi_2
X_21034_ _12804_ _12805_ VGND VGND VPWR VPWR _12881_ sky130_fd_sc_hd__and2_1
Xfanout123 net124 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26891_ clknet_leaf_105_clk_sys _00508_ net577 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout134 top0.cordic0.vec\[1\]\[6\] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_2
Xfanout145 top0.cordic0.vec\[1\]\[4\] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_4
Xfanout156 net157 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_4
Xfanout167 top0.cordic0.vec\[1\]\[0\] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_2
X_25842_ net76 _05059_ _05058_ top0.matmul0.beta_pass\[5\] VGND VGND VPWR VPWR _05064_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout178 top0.cordic0.state\[0\] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__buf_2
Xfanout189 net190 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25773_ _05007_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22985_ _02491_ _02487_ _02492_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__a21o_1
XFILLER_0_198_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24724_ _04071_ _04076_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21936_ _01267_ _01330_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24655_ _03868_ _03877_ _03872_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_167_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21867_ _01422_ _01427_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__and2_1
XFILLER_0_171_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23606_ top0.matmul0.alpha_pass\[10\] _09308_ net559 VGND VGND VPWR VPWR _02970_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20818_ _12535_ _12539_ _12661_ _12663_ _12666_ VGND VGND VPWR VPWR _12667_ sky130_fd_sc_hd__a221o_1
X_24586_ _03768_ _03769_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__nand2_1
X_21798_ _01357_ _01359_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26325_ _05394_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__clkbuf_1
X_23537_ _02934_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20749_ _12593_ _12594_ _12596_ _12597_ VGND VGND VPWR VPWR _12598_ sky130_fd_sc_hd__or4_4
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14270_ _06419_ _06420_ _06477_ _06478_ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__o22a_1
X_26256_ spi0.data_packed\[26\] spi0.data_packed\[27\] net699 VGND VGND VPWR VPWR
+ _05360_ sky130_fd_sc_hd__mux2_1
X_23468_ _02898_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25207_ _04483_ _04488_ _04480_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__a21bo_1
X_13221_ _05445_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__clkbuf_1
X_22419_ _01971_ _01976_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__xnor2_1
X_26187_ net18 _05321_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23399_ net112 _02827_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25138_ _03900_ _04190_ _03889_ _03758_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25069_ _04411_ _04417_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17960_ _09942_ _09945_ VGND VGND VPWR VPWR _09946_ sky130_fd_sc_hd__xnor2_2
X_16911_ top0.currT_r\[6\] _08959_ _08970_ VGND VGND VPWR VPWR _08971_ sky130_fd_sc_hd__a21o_1
X_17891_ _09874_ _09877_ VGND VGND VPWR VPWR _09878_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19630_ _11518_ VGND VGND VPWR VPWR _11519_ sky130_fd_sc_hd__buf_4
X_16842_ _08905_ _08906_ net547 VGND VGND VPWR VPWR _08907_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout690 net692 VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19561_ net160 net156 net150 net144 net197 net191 VGND VGND VPWR VPWR _11450_ sky130_fd_sc_hd__mux4_2
X_13985_ _06186_ _06197_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__xnor2_2
X_16773_ _08855_ VGND VGND VPWR VPWR _08856_ sky130_fd_sc_hd__buf_2
XFILLER_0_176_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18512_ _10394_ _10397_ _10491_ VGND VGND VPWR VPWR _10492_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15724_ net505 net488 VGND VGND VPWR VPWR _07821_ sky130_fd_sc_hd__nand2_1
X_19492_ top0.pid_d.curr_int\[13\] top0.pid_d.prev_int\[13\] VGND VGND VPWR VPWR _11385_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_198_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18443_ net434 _10341_ _10342_ _10423_ net436 VGND VGND VPWR VPWR _10424_ sky130_fd_sc_hd__a32o_1
XFILLER_0_197_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15655_ _07751_ _07752_ VGND VGND VPWR VPWR _07753_ sky130_fd_sc_hd__xor2_1
X_14606_ _06697_ _06809_ _06810_ VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__o21ai_1
X_18374_ _10353_ _10354_ VGND VGND VPWR VPWR _10355_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15586_ _07543_ _07544_ _07533_ _07534_ VGND VGND VPWR VPWR _07685_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14537_ _06652_ _06614_ _06743_ VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__o21ai_4
X_17325_ top0.matmul0.matmul_stage_inst.mult1\[11\] top0.matmul0.matmul_stage_inst.mult2\[11\]
+ VGND VGND VPWR VPWR _09316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14468_ _06554_ _06608_ _06609_ VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__o21ba_1
X_17256_ top0.matmul0.matmul_stage_inst.mult1\[0\] top0.matmul0.matmul_stage_inst.mult2\[0\]
+ top0.matmul0.matmul_stage_inst.mult2\[1\] VGND VGND VPWR VPWR _09257_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13419_ _05621_ _05622_ net65 VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__a21o_1
X_16207_ _08167_ _08172_ _08049_ VGND VGND VPWR VPWR _08299_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17187_ _09195_ _09196_ VGND VGND VPWR VPWR _09198_ sky130_fd_sc_hd__or2_1
X_14399_ _06603_ _06607_ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16138_ _08165_ _08230_ VGND VGND VPWR VPWR _08231_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16069_ _08153_ _08155_ VGND VGND VPWR VPWR _08162_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19828_ _11705_ _11706_ VGND VGND VPWR VPWR _11707_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19759_ _11518_ _11641_ VGND VGND VPWR VPWR _11642_ sky130_fd_sc_hd__or2_1
X_22770_ top0.pid_q.prev_int\[14\] _02291_ _02294_ top0.pid_q.curr_int\[14\] VGND
+ VGND VPWR VPWR _00433_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21721_ net153 _01280_ _01281_ _01282_ net167 VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24440_ _03794_ _03788_ _03789_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__or3_1
XFILLER_0_115_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21652_ _01213_ _01112_ net105 VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20603_ _12430_ _12431_ VGND VGND VPWR VPWR _12452_ sky130_fd_sc_hd__nor2_1
X_24371_ _03726_ _03727_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21583_ _01144_ _01115_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_191_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26110_ top0.periodTop\[9\] _05276_ _05278_ net42 VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__a22o_1
X_23322_ _02766_ _02767_ _01105_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__mux2_1
X_27090_ clknet_leaf_1_clk_sys _00707_ net584 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.b\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_20534_ _12381_ _12382_ VGND VGND VPWR VPWR _12383_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26041_ _12031_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__buf_2
XFILLER_0_90_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23253_ net165 net1016 _02669_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__and3_1
X_20465_ _12292_ _12299_ _12313_ VGND VGND VPWR VPWR _12314_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_104_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22204_ _01756_ _01764_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__xnor2_4
X_23184_ _02646_ _06473_ _02649_ net835 VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__a22o_1
X_20396_ net264 net253 net240 VGND VGND VPWR VPWR _12245_ sky130_fd_sc_hd__and3_1
X_22135_ _01210_ _01227_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__nand2_1
X_22066_ _01620_ _01624_ _01625_ _01626_ _01627_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__o2111a_2
X_26943_ clknet_leaf_9_clk_sys _00560_ net594 VGND VGND VPWR VPWR top0.matmul0.a\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_21017_ _12861_ _12863_ VGND VGND VPWR VPWR _12864_ sky130_fd_sc_hd__xnor2_2
X_26874_ clknet_leaf_40_clk_sys _00491_ net682 VGND VGND VPWR VPWR top0.svm0.tB\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25825_ top0.c_out_calc\[3\] _05029_ _05031_ _05049_ VGND VGND VPWR VPWR _00734_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13770_ _05941_ _05982_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__xnor2_1
X_25756_ top0.matmul0.matmul_stage_inst.a\[6\] _04894_ _05458_ VGND VGND VPWR VPWR
+ _04999_ sky130_fd_sc_hd__mux2_1
X_22968_ top0.svm0.delta\[6\] VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__inv_2
X_24707_ _04059_ _04060_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__or2b_1
X_21919_ _01458_ _01393_ net165 VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__a21oi_1
X_25687_ _04885_ _04954_ _04883_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__mux2_1
X_22899_ _02324_ top0.svm0.tC\[6\] top0.svm0.tC\[5\] _02415_ _02416_ VGND VGND VPWR
+ VPWR _02417_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15440_ _07274_ _07276_ net484 VGND VGND VPWR VPWR _07539_ sky130_fd_sc_hd__o21a_1
XFILLER_0_167_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24638_ _03990_ _03970_ _03971_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__nand3_2
XFILLER_0_195_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15371_ _07436_ _07437_ _07438_ VGND VGND VPWR VPWR _07470_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24569_ _03797_ _03812_ _03923_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_26_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14322_ _06481_ _06531_ VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__xnor2_1
X_17110_ net873 _09114_ _09131_ VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18090_ net356 net361 VGND VGND VPWR VPWR _10074_ sky130_fd_sc_hd__xor2_4
X_26308_ spi0.data_packed\[52\] spi0.data_packed\[53\] net697 VGND VGND VPWR VPWR
+ _05386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27288_ clknet_3_0__leaf_clk_mosi _00902_ VGND VGND VPWR VPWR spi0.data_packed\[74\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17041_ _09091_ _09092_ VGND VGND VPWR VPWR _09093_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14253_ _06462_ _06463_ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__or2_2
XFILLER_0_29_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26239_ _05351_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13204_ top0.matmul0.done_pass VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14184_ net44 _05602_ _05603_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18992_ _10865_ _10866_ VGND VGND VPWR VPWR _10966_ sky130_fd_sc_hd__nand2_1
X_17943_ _09923_ _09928_ VGND VGND VPWR VPWR _09929_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_178_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17874_ _09764_ _09761_ _09860_ VGND VGND VPWR VPWR _09861_ sky130_fd_sc_hd__a21o_1
X_19613_ _11469_ _11471_ VGND VGND VPWR VPWR _11502_ sky130_fd_sc_hd__nor2_1
X_16825_ top0.currT_r\[0\] top0.matmul0.beta_pass\[0\] VGND VGND VPWR VPWR _08891_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19544_ _11433_ _11430_ VGND VGND VPWR VPWR _11434_ sky130_fd_sc_hd__nor2_1
X_16756_ _08787_ _08839_ VGND VGND VPWR VPWR _08840_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13968_ _06118_ _06180_ _06102_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_158_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15707_ _07802_ _07803_ VGND VGND VPWR VPWR _07804_ sky130_fd_sc_hd__nand2_1
X_19475_ _11368_ _11369_ VGND VGND VPWR VPWR _11370_ sky130_fd_sc_hd__nand2_1
X_13899_ net40 _05472_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__nand2_1
X_16687_ net452 net455 net500 net449 VGND VGND VPWR VPWR _08772_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_201_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18426_ net416 _09365_ _10228_ VGND VGND VPWR VPWR _10407_ sky130_fd_sc_hd__or3_2
XFILLER_0_75_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15638_ _07623_ _07628_ _07735_ VGND VGND VPWR VPWR _07736_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18357_ _10337_ _10246_ top0.pid_d.out\[5\] VGND VGND VPWR VPWR _10338_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15569_ net511 _07667_ VGND VGND VPWR VPWR _07668_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17308_ _09300_ _09301_ VGND VGND VPWR VPWR _09302_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18288_ _10256_ _10269_ VGND VGND VPWR VPWR _10270_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17239_ _08791_ _09192_ _09242_ net1019 _09243_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20250_ _12097_ _12092_ _12093_ VGND VGND VPWR VPWR _12099_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20181_ _12009_ _12030_ VGND VGND VPWR VPWR _12031_ sky130_fd_sc_hd__nor2_2
XFILLER_0_177_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23940_ _03292_ _03295_ _03296_ _03297_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__and4bb_1
X_23871_ _03131_ _03137_ _03227_ _03228_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__o211ai_4
X_25610_ net70 top0.matmul0.cos\[8\] VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__and2_1
X_22822_ top0.svm0.counter\[10\] top0.svm0.tA\[10\] VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__and2b_1
XFILLER_0_193_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26590_ clknet_leaf_65_clk_sys _00213_ net660 VGND VGND VPWR VPWR top0.pid_q.curr_int\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_17_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25541_ _04857_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__clkbuf_1
X_22753_ net549 _05442_ net13 net545 VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__and4b_1
XFILLER_0_39_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21704_ net158 VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__inv_2
X_25472_ _04721_ _04750_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__nand2_1
XFILLER_0_177_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22684_ _12963_ _02234_ _02235_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24423_ _03713_ _03708_ _03778_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27211_ clknet_leaf_6_clk_sys _00825_ net591 VGND VGND VPWR VPWR top0.cordic0.slte0.opB\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_21635_ _01087_ _01172_ _01196_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27142_ clknet_leaf_14_clk_sys _00756_ net620 VGND VGND VPWR VPWR top0.b_in_matmul\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24354_ _03004_ _03005_ _03061_ _03062_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__o22a_1
X_21566_ _01114_ _01127_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_77_clk_sys clknet_3_1__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_77_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_23305_ _02688_ _02689_ _11573_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__mux2_1
X_27073_ clknet_leaf_21_clk_sys _00690_ net610 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.c\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_20517_ _12266_ _12362_ _12365_ VGND VGND VPWR VPWR _12366_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_7_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24285_ top0.matmul0.matmul_stage_inst.mult2\[0\] _03641_ _03642_ VGND VGND VPWR
+ VPWR _03643_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21497_ _01058_ _12883_ _01057_ VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__mux2_1
X_26024_ top0.pid_q.out\[15\] _05198_ _05199_ spi0.data_packed\[63\] VGND VGND VPWR
+ VPWR _05219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23236_ _02678_ _02682_ _02684_ _02685_ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__nand4_2
XFILLER_0_132_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20448_ net283 _12065_ VGND VGND VPWR VPWR _12297_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23167_ _02641_ _06682_ _02645_ net894 VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__a22o_1
X_20379_ _12218_ _12219_ _12227_ VGND VGND VPWR VPWR _12228_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22118_ _01653_ _01645_ _01660_ _01640_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__a211oi_1
X_23098_ top0.svm0.delta\[1\] net555 _02598_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__and3b_1
XFILLER_0_98_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22049_ _01599_ _01604_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__nand2_1
X_14940_ _07091_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__clkbuf_1
X_26926_ clknet_leaf_4_clk_sys _00543_ net580 VGND VGND VPWR VPWR top0.matmul0.cos\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26857_ clknet_leaf_38_clk_sys _00474_ net677 VGND VGND VPWR VPWR top0.svm0.calc_ready
+ sky130_fd_sc_hd__dfrtp_1
X_14871_ _07055_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__clkbuf_1
X_16610_ net452 net455 VGND VGND VPWR VPWR _08696_ sky130_fd_sc_hd__xor2_1
X_25808_ top0.matmul0.alpha_pass\[0\] top0.matmul0.beta_pass\[0\] VGND VGND VPWR VPWR
+ _05035_ sky130_fd_sc_hd__nor2_1
X_13822_ _06029_ _06034_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17590_ net425 _09550_ _09576_ net418 VGND VGND VPWR VPWR _09577_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26788_ clknet_leaf_3_clk_sys _00405_ net583 VGND VGND VPWR VPWR top0.cordic0.sin\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_13753_ net67 _05587_ _05534_ _05607_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__a211o_1
X_16541_ _08567_ _08577_ _08569_ VGND VGND VPWR VPWR _08628_ sky130_fd_sc_hd__o21a_1
X_25739_ net786 _04890_ _04913_ _04990_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19260_ _11203_ _11196_ _11204_ VGND VGND VPWR VPWR _11205_ sky130_fd_sc_hd__a21o_1
X_16472_ _08501_ _08503_ _08559_ VGND VGND VPWR VPWR _08560_ sky130_fd_sc_hd__a21oi_2
X_13684_ net1027 _05497_ _05895_ _05896_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18211_ _10098_ _10100_ _10193_ VGND VGND VPWR VPWR _10194_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_39_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15423_ _07380_ _07381_ _07376_ VGND VGND VPWR VPWR _07522_ sky130_fd_sc_hd__a21o_1
X_19191_ net351 _11094_ VGND VGND VPWR VPWR _11143_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18142_ _10114_ _10125_ VGND VGND VPWR VPWR _10126_ sky130_fd_sc_hd__xnor2_1
X_15354_ _07442_ _07449_ _07450_ _07452_ VGND VGND VPWR VPWR _07453_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14305_ net28 net1015 VGND VGND VPWR VPWR _06515_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18073_ _10053_ _10057_ VGND VGND VPWR VPWR _10058_ sky130_fd_sc_hd__xnor2_1
X_15285_ _07321_ _07374_ _07383_ VGND VGND VPWR VPWR _07384_ sky130_fd_sc_hd__a21o_1
XFILLER_0_202_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_184_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14236_ _06444_ _06445_ _06433_ _06434_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__a211o_1
Xhold209 top0.pid_q.prev_error\[12\] VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__dlygate4sd3_1
X_17024_ _09073_ _09076_ VGND VGND VPWR VPWR _09077_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14167_ _06178_ _06372_ _06378_ VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_1_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14098_ _06306_ _06309_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__xor2_1
X_18975_ net316 _10946_ _10948_ VGND VGND VPWR VPWR _10949_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_13_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17926_ net1023 net413 VGND VGND VPWR VPWR _09912_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17857_ net351 net380 VGND VGND VPWR VPWR _09844_ sky130_fd_sc_hd__nand2_2
X_16808_ net505 _08855_ _08858_ net703 _08877_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__a221o_1
X_17788_ _09767_ _09774_ VGND VGND VPWR VPWR _09775_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_191_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19527_ net144 net138 net133 net128 net197 net191 VGND VGND VPWR VPWR _11417_ sky130_fd_sc_hd__mux4_1
X_16739_ net445 net444 net504 VGND VGND VPWR VPWR _08823_ sky130_fd_sc_hd__and3b_1
XFILLER_0_89_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19458_ _11353_ _11354_ VGND VGND VPWR VPWR _11355_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18409_ _10383_ _10389_ VGND VGND VPWR VPWR _10390_ sky130_fd_sc_hd__xnor2_1
X_19389_ net439 _11118_ _11294_ net442 VGND VGND VPWR VPWR _11295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_189_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21420_ _00984_ _00986_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21351_ _13110_ _00918_ _00919_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20302_ _12148_ _12149_ _12133_ VGND VGND VPWR VPWR _12151_ sky130_fd_sc_hd__a21o_1
X_24070_ _03426_ _03374_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__nor2_1
X_21282_ net251 net229 VGND VGND VPWR VPWR _13125_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_188_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout3 _11439_ VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__clkbuf_4
X_23021_ _06277_ _02523_ net172 VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20233_ _12041_ _12079_ _12081_ VGND VGND VPWR VPWR _12082_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_31_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20164_ net207 _12015_ VGND VGND VPWR VPWR _12016_ sky130_fd_sc_hd__nand2_1
X_24972_ _04237_ _04239_ _04168_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__o21a_1
XFILLER_0_157_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20095_ _11649_ _11952_ _11954_ VGND VGND VPWR VPWR _11955_ sky130_fd_sc_hd__a21o_1
X_26711_ clknet_leaf_72_clk_sys _00328_ net655 VGND VGND VPWR VPWR top0.pid_d.curr_int\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_23923_ _03280_ _03149_ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23854_ _03210_ _03211_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__xor2_1
X_26642_ clknet_leaf_80_clk_sys _00259_ net634 VGND VGND VPWR VPWR top0.pid_d.out\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_22805_ _02324_ top0.svm0.tA\[6\] VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23785_ _03049_ _03050_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__nand2_1
X_26573_ clknet_leaf_55_clk_sys _00196_ net667 VGND VGND VPWR VPWR top0.pid_q.curr_error\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_40_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20997_ net255 net259 VGND VGND VPWR VPWR _12844_ sky130_fd_sc_hd__or2b_1
X_25524_ _04848_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__clkbuf_1
X_22736_ _02282_ _12012_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25455_ _04733_ _04797_ _04732_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__o21a_1
X_22667_ _01223_ _02218_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24406_ _03760_ _03761_ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_180_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21618_ _01176_ _01177_ _01175_ _01179_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_180_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25386_ _04518_ _04729_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__nor2_1
XFILLER_0_180_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22598_ _02146_ _02151_ _01074_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_27125_ clknet_leaf_33_clk_sys _00739_ net665 VGND VGND VPWR VPWR top0.c_out_calc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_24337_ _03684_ _03693_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__xor2_4
XFILLER_0_129_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21549_ net77 net102 VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__xor2_1
X_27056_ clknet_leaf_20_clk_sys _00673_ net609 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.d\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_15070_ net533 net475 VGND VGND VPWR VPWR _07169_ sky130_fd_sc_hd__nand2_2
X_24268_ _03624_ _03625_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14021_ _06111_ _06116_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__nor2_1
X_26007_ _05206_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__clkbuf_1
X_23219_ _01320_ _11515_ VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__nor2_1
X_24199_ _03500_ _03556_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__xnor2_1
X_18760_ _09771_ _10495_ _10736_ net309 _09493_ VGND VGND VPWR VPWR _10737_ sky130_fd_sc_hd__a221o_1
X_15972_ _08064_ _08066_ VGND VGND VPWR VPWR _08067_ sky130_fd_sc_hd__xor2_1
X_17711_ _09475_ _09478_ _09697_ VGND VGND VPWR VPWR _09698_ sky130_fd_sc_hd__o21ai_2
X_14923_ _07082_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__clkbuf_1
X_26909_ clknet_leaf_110_clk_sys _00526_ net579 VGND VGND VPWR VPWR top0.matmul0.sin\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_117_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18691_ _10667_ _10668_ VGND VGND VPWR VPWR _10669_ sky130_fd_sc_hd__nor2_1
Xhold70 top0.matmul0.matmul_stage_inst.a\[3\] VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 top0.svm0.tA\[10\] VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold92 top0.matmul0.matmul_stage_inst.b\[7\] VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__dlygate4sd3_1
X_17642_ net419 net330 net337 net412 VGND VGND VPWR VPWR _09629_ sky130_fd_sc_hd__a22o_1
X_14854_ _07046_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13805_ _05983_ _05970_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__xor2_1
XFILLER_0_187_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17573_ _09529_ _09559_ net415 _09401_ VGND VGND VPWR VPWR _09560_ sky130_fd_sc_hd__a2bb2o_1
X_14785_ net34 _06867_ _06984_ VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__and3_1
XFILLER_0_202_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19312_ _11247_ _11123_ _11252_ VGND VGND VPWR VPWR _11253_ sky130_fd_sc_hd__or3b_1
XFILLER_0_86_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16524_ top0.pid_q.out\[10\] top0.pid_q.curr_int\[10\] VGND VGND VPWR VPWR _08612_
+ sky130_fd_sc_hd__and2_1
X_13736_ _05924_ _05926_ _05948_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19243_ top0.matmul0.alpha_pass\[7\] _11180_ VGND VGND VPWR VPWR _11190_ sky130_fd_sc_hd__or2_1
X_16455_ _08467_ _08470_ VGND VGND VPWR VPWR _08544_ sky130_fd_sc_hd__nor2_1
X_13667_ _05863_ _05874_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_171_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15406_ net484 _07473_ _07474_ VGND VGND VPWR VPWR _07505_ sky130_fd_sc_hd__a21o_1
X_19174_ top0.pid_d.prev_error\[0\] top0.pid_d.curr_error\[0\] _11126_ VGND VGND VPWR
+ VPWR _11127_ sky130_fd_sc_hd__and3_1
X_13598_ _05657_ _05543_ _05545_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__or3_2
XFILLER_0_143_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16386_ _08334_ _08475_ _08307_ VGND VGND VPWR VPWR _08476_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_27_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18125_ _10107_ _10108_ VGND VGND VPWR VPWR _10109_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15337_ net528 net495 VGND VGND VPWR VPWR _07436_ sky130_fd_sc_hd__nand2_4
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1 _01123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18056_ _09951_ _09954_ _09948_ VGND VGND VPWR VPWR _10041_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_41_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15268_ _07366_ net479 VGND VGND VPWR VPWR _07367_ sky130_fd_sc_hd__nor2_1
X_17007_ top0.currT_r\[13\] _09060_ VGND VGND VPWR VPWR _09061_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14219_ _06306_ _06308_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__and2b_1
XFILLER_0_50_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15199_ _07281_ _07297_ VGND VGND VPWR VPWR _07298_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_1_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout508 net509 VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__clkbuf_4
Xfanout519 top0.pid_q.mult0.a\[8\] VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__clkbuf_2
X_18958_ _10875_ _10931_ _10804_ VGND VGND VPWR VPWR _10932_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_174_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_25_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_25_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_17909_ _09895_ _07138_ VGND VGND VPWR VPWR _09896_ sky130_fd_sc_hd__nor2_1
X_18889_ net365 _10863_ VGND VGND VPWR VPWR _10864_ sky130_fd_sc_hd__nand2_1
X_20920_ _11726_ _12763_ _12766_ _12767_ VGND VGND VPWR VPWR _12768_ sky130_fd_sc_hd__o31a_1
XFILLER_0_179_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_clk_mosi clk_mosi VGND VGND VPWR VPWR clknet_0_clk_mosi sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20851_ net229 _12699_ VGND VGND VPWR VPWR _12700_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23570_ top0.b_in_matmul\[8\] top0.matmul0.b\[8\] _02948_ VGND VGND VPWR VPWR _02952_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20782_ _12142_ _12623_ _12468_ net299 _12630_ VGND VGND VPWR VPWR _12631_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22521_ _02051_ _02076_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25240_ _04515_ _04521_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__xor2_1
XFILLER_0_123_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22452_ _01979_ _01982_ _02008_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_17_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21403_ _00969_ _12764_ _00942_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25171_ _03355_ _04252_ _04258_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__a21oi_1
X_22383_ _01898_ _01941_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24122_ _03400_ _03479_ _03408_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__or3_1
XFILLER_0_130_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21334_ _13173_ _13175_ VGND VGND VPWR VPWR _13176_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24053_ _03398_ _03400_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__nand2_1
X_21265_ net762 _12034_ _12037_ _13108_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23004_ _02508_ _02504_ _02345_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__a21o_1
XFILLER_0_198_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20216_ net297 net290 VGND VGND VPWR VPWR _12065_ sky130_fd_sc_hd__nand2_4
XFILLER_0_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21196_ _13027_ _13039_ VGND VGND VPWR VPWR _13040_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_159_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20147_ _11983_ _11649_ _11954_ VGND VGND VPWR VPWR _12002_ sky130_fd_sc_hd__a21o_1
X_24955_ _03549_ _04176_ _03829_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__o21ai_4
X_20078_ _11715_ _11938_ VGND VGND VPWR VPWR _11939_ sky130_fd_sc_hd__nor2_1
X_23906_ _03237_ _03242_ _03246_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__o21a_1
XFILLER_0_169_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24886_ _04130_ _04135_ _04138_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26625_ clknet_leaf_31_clk_sys _00242_ net619 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_23837_ _03088_ _03089_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__nor2_4
XFILLER_0_197_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14570_ _05586_ _06640_ VGND VGND VPWR VPWR _06776_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_197_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26556_ clknet_leaf_49_clk_sys _00179_ net675 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_23768_ _03078_ _03079_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__and2_1
XFILLER_0_178_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25507_ _04839_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__clkbuf_1
X_13521_ _05656_ _05732_ _05733_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__o21a_1
XFILLER_0_137_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22719_ _12036_ _02269_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__nor2_1
X_23699_ net574 net566 top0.matmul0.matmul_stage_inst.a\[3\] VGND VGND VPWR VPWR _03057_
+ sky130_fd_sc_hd__o21a_2
X_26487_ clknet_leaf_66_clk_sys _00007_ net660 VGND VGND VPWR VPWR top0.pid_q.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13452_ _05663_ _05664_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__and2_1
X_16240_ _08309_ VGND VGND VPWR VPWR _08331_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25438_ _03123_ _03889_ _03124_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_165_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25369_ _04406_ _04698_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__and2_1
X_13383_ _05527_ _05595_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__xnor2_4
X_16171_ net450 net1028 VGND VGND VPWR VPWR _08263_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15122_ _07217_ _07218_ _07196_ VGND VGND VPWR VPWR _07221_ sky130_fd_sc_hd__a21oi_1
X_27108_ clknet_leaf_8_clk_sys _00725_ net592 VGND VGND VPWR VPWR top0.matmul0.op\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19930_ net901 _11800_ _11801_ _11799_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__a22o_1
X_15053_ net534 net470 VGND VGND VPWR VPWR _07152_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27039_ clknet_leaf_7_clk_sys _00656_ net592 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14004_ net1030 VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19861_ net1013 _11736_ _11727_ VGND VGND VPWR VPWR _11738_ sky130_fd_sc_hd__a21oi_1
X_18812_ _10718_ _10716_ _10723_ VGND VGND VPWR VPWR _10788_ sky130_fd_sc_hd__nor3_1
XFILLER_0_128_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19792_ _11672_ VGND VGND VPWR VPWR _11673_ sky130_fd_sc_hd__buf_2
XFILLER_0_179_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18743_ _09377_ _10719_ VGND VGND VPWR VPWR _10720_ sky130_fd_sc_hd__or2_1
X_15955_ _08047_ _08049_ VGND VGND VPWR VPWR _08050_ sky130_fd_sc_hd__nor2_1
X_14906_ _07073_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__clkbuf_1
X_18674_ _10649_ _10651_ VGND VGND VPWR VPWR _10652_ sky130_fd_sc_hd__nor2_1
X_15886_ _07980_ _07880_ VGND VGND VPWR VPWR _07982_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17625_ net1022 net420 VGND VGND VPWR VPWR _09612_ sky130_fd_sc_hd__nand2_2
XFILLER_0_76_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14837_ _06955_ _07013_ _07014_ VGND VGND VPWR VPWR _07035_ sky130_fd_sc_hd__and3b_1
XFILLER_0_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_175_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17556_ _09537_ _09539_ _09542_ VGND VGND VPWR VPWR _09543_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14768_ _06949_ _06969_ VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16507_ _08593_ _08594_ VGND VGND VPWR VPWR _08595_ sky130_fd_sc_hd__xnor2_1
X_13719_ net1027 _05488_ _05490_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17487_ net408 net343 net347 net403 VGND VGND VPWR VPWR _09474_ sky130_fd_sc_hd__a22o_1
X_14699_ _06866_ _06902_ VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_184_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19226_ _11173_ _11166_ top0.pid_d.prev_error\[5\] VGND VGND VPWR VPWR _11174_ sky130_fd_sc_hd__o21ba_1
X_16438_ _08453_ _08526_ VGND VGND VPWR VPWR _08527_ sky130_fd_sc_hd__nor2_4
XFILLER_0_2_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19157_ top0.kid\[13\] _11097_ _11099_ top0.kpd\[13\] VGND VGND VPWR VPWR _11114_
+ sky130_fd_sc_hd__a22o_1
X_16369_ _08442_ _08458_ VGND VGND VPWR VPWR _08459_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18108_ _10090_ _10091_ VGND VGND VPWR VPWR _10092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19088_ net365 _11059_ VGND VGND VPWR VPWR _11060_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18039_ _09909_ _09914_ _10023_ VGND VGND VPWR VPWR _10024_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21050_ net222 _12827_ _12894_ _12773_ _12895_ VGND VGND VPWR VPWR _12896_ sky130_fd_sc_hd__o221a_1
Xfanout305 net306 VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__clkbuf_2
Xfanout316 net317 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__buf_2
X_20001_ top0.cordic0.slte0.opA\[4\] net1012 VGND VGND VPWR VPWR _11868_ sky130_fd_sc_hd__or2_1
Xfanout327 net1022 VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__clkbuf_4
Xfanout338 net339 VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__buf_4
XFILLER_0_185_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout349 net350 VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__buf_2
XFILLER_0_185_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24740_ _04091_ _04092_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__xnor2_1
X_21952_ _01511_ _01513_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__nor2_1
X_20903_ _12717_ _12750_ _12695_ VGND VGND VPWR VPWR _12751_ sky130_fd_sc_hd__o21a_1
X_24671_ _04021_ _04024_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__xnor2_1
X_21883_ _01432_ _01435_ _01444_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23622_ net570 top0.matmul0.matmul_stage_inst.b\[8\] top0.matmul0.matmul_stage_inst.a\[8\]
+ net567 VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__a22o_4
XFILLER_0_77_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26410_ clknet_leaf_85_clk_sys _00051_ net640 VGND VGND VPWR VPWR top0.kpd\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_20834_ net229 net221 VGND VGND VPWR VPWR _12683_ sky130_fd_sc_hd__nand2_4
XFILLER_0_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23553_ top0.b_in_matmul\[0\] top0.matmul0.b\[0\] _02937_ VGND VGND VPWR VPWR _02943_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26341_ _05402_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20765_ _12348_ _12584_ VGND VGND VPWR VPWR _12614_ sky130_fd_sc_hd__or2_2
XFILLER_0_175_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22504_ net107 _01312_ _02054_ _02055_ _02059_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__a311o_2
XFILLER_0_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26272_ net944 spi0.data_packed\[35\] net688 VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23484_ top0.cordic0.sin\[11\] top0.matmul0.sin\[11\] _02904_ VGND VGND VPWR VPWR
+ _02907_ sky130_fd_sc_hd__mux2_1
X_20696_ _12515_ _12531_ _12532_ VGND VGND VPWR VPWR _12545_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25223_ _04492_ _04504_ _04569_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__o21a_1
XFILLER_0_165_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22435_ _01885_ _01898_ _01941_ _01992_ _01877_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__a311o_1
XFILLER_0_162_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25154_ _04498_ _04500_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__nand2_1
X_22366_ net86 _01248_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24105_ _03355_ _03324_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__nand2_1
X_21317_ _13112_ _13134_ _13158_ VGND VGND VPWR VPWR _13159_ sky130_fd_sc_hd__a21o_1
X_25085_ _04424_ _04433_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__xnor2_1
X_22297_ _01843_ _01855_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__nand2_1
X_24036_ _03355_ _03217_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__nand2_2
X_21248_ _13088_ _13090_ _13091_ _12541_ VGND VGND VPWR VPWR _13092_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_102_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21179_ _11689_ _12982_ VGND VGND VPWR VPWR _13023_ sky130_fd_sc_hd__nand2_1
X_25987_ _05190_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15740_ _07833_ _07836_ VGND VGND VPWR VPWR _07837_ sky130_fd_sc_hd__xnor2_1
X_24938_ _03325_ _04288_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15671_ net490 net486 net508 _07768_ VGND VGND VPWR VPWR _07769_ sky130_fd_sc_hd__a31o_1
X_24869_ _04219_ _04220_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_198_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17410_ net400 net395 _09396_ VGND VGND VPWR VPWR _09397_ sky130_fd_sc_hd__a21o_1
X_14622_ net41 _06268_ VGND VGND VPWR VPWR _06827_ sky130_fd_sc_hd__nand2_1
X_26608_ clknet_leaf_83_clk_sys _00003_ net641 VGND VGND VPWR VPWR top0.pid_d.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_18390_ _10278_ _10280_ _10370_ VGND VGND VPWR VPWR _10371_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_200_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17341_ top0.matmul0.matmul_stage_inst.mult1\[14\] top0.matmul0.matmul_stage_inst.mult2\[14\]
+ VGND VGND VPWR VPWR _09330_ sky130_fd_sc_hd__xor2_1
X_14553_ net23 _05579_ _06643_ VGND VGND VPWR VPWR _06759_ sky130_fd_sc_hd__and3_1
X_26539_ clknet_leaf_60_clk_sys _00162_ net668 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13504_ _05474_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__buf_6
XFILLER_0_165_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17272_ top0.matmul0.matmul_stage_inst.mult1\[4\] top0.matmul0.matmul_stage_inst.mult2\[4\]
+ VGND VGND VPWR VPWR _09271_ sky130_fd_sc_hd__xor2_1
XFILLER_0_55_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14484_ _06685_ _06690_ VGND VGND VPWR VPWR _06691_ sky130_fd_sc_hd__and2_2
XFILLER_0_125_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19011_ _10927_ _10984_ VGND VGND VPWR VPWR _10985_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16223_ _08254_ _08314_ VGND VGND VPWR VPWR _08315_ sky130_fd_sc_hd__xnor2_1
X_13435_ _05559_ _05598_ _05647_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_64_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13366_ _05551_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16154_ top0.pid_q.out\[7\] top0.pid_q.curr_int\[7\] VGND VGND VPWR VPWR _08246_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15105_ net494 net511 VGND VGND VPWR VPWR _07204_ sky130_fd_sc_hd__nand2_2
X_13297_ net42 _05497_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__nand2_1
X_16085_ _08123_ _08128_ _08177_ VGND VGND VPWR VPWR _08178_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19913_ net224 _11782_ _11786_ _11781_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__a22o_1
X_15036_ net938 _07140_ _07144_ top0.pid_d.curr_int\[6\] VGND VGND VPWR VPWR _00123_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19844_ _11713_ _11721_ VGND VGND VPWR VPWR _11722_ sky130_fd_sc_hd__xor2_1
X_19775_ _11656_ VGND VGND VPWR VPWR _11657_ sky130_fd_sc_hd__buf_2
X_16987_ top0.currT_r\[12\] VGND VGND VPWR VPWR _09042_ sky130_fd_sc_hd__inv_2
X_18726_ _10701_ _10702_ net362 VGND VGND VPWR VPWR _10703_ sky130_fd_sc_hd__o21a_1
X_15938_ _07938_ _07940_ _08032_ VGND VGND VPWR VPWR _08033_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_79_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18657_ _10537_ _10539_ _10634_ VGND VGND VPWR VPWR _10635_ sky130_fd_sc_hd__a21bo_1
X_15869_ _07832_ _07864_ _07865_ VGND VGND VPWR VPWR _07965_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_188_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17608_ _09551_ _09553_ VGND VGND VPWR VPWR _09595_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18588_ net406 _09353_ _09351_ _10228_ VGND VGND VPWR VPWR _10567_ sky130_fd_sc_hd__or4_2
XFILLER_0_153_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17539_ net340 _09524_ _09525_ VGND VGND VPWR VPWR _09526_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20550_ _12386_ _12388_ _12395_ _12398_ VGND VGND VPWR VPWR _12399_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_156_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19209_ _11158_ VGND VGND VPWR VPWR _11159_ sky130_fd_sc_hd__inv_2
X_20481_ net304 _12329_ VGND VGND VPWR VPWR _12330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22220_ _01716_ _01780_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22151_ net99 _01223_ net110 net105 VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__and4bb_1
XPHY_EDGE_ROW_5_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21102_ _12746_ _12943_ _12749_ VGND VGND VPWR VPWR _12948_ sky130_fd_sc_hd__a21oi_1
X_22082_ _01641_ _01643_ _01615_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout102 top0.cordic0.vec\[1\]\[13\] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_4
X_25910_ _05120_ _05121_ _05601_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__a21o_1
X_21033_ _12675_ _12807_ VGND VGND VPWR VPWR _12880_ sky130_fd_sc_hd__or2_1
Xfanout113 top0.cordic0.vec\[1\]\[11\] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_4
XFILLER_0_201_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout124 net125 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_4
Xfanout135 net137 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_4
X_26890_ clknet_leaf_105_clk_sys _00507_ net577 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout146 net148 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_201_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout157 top0.cordic0.vec\[1\]\[2\] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
Xfanout168 top0.svm0.counter\[14\] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_4
X_25841_ top0.matmul0.beta_pass\[5\] _05058_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__or2_1
Xfanout179 net180 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_198_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22984_ _02491_ _02487_ _02367_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__o21a_1
X_25772_ top0.matmul0.op_in\[0\] net74 _05460_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__mux2_1
X_24723_ _04072_ _04075_ VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_201_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21935_ net136 _01496_ _01267_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24654_ _04005_ _04006_ _04000_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__a21oi_1
X_21866_ _01422_ _01427_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23605_ _02969_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__clkbuf_1
X_20817_ _12460_ _12461_ _12540_ _12533_ _12665_ VGND VGND VPWR VPWR _12666_ sky130_fd_sc_hd__a32o_1
XFILLER_0_166_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24585_ _03768_ _03769_ _03770_ VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__o21ai_2
X_21797_ _01177_ _01358_ net162 VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__o21a_1
XFILLER_0_194_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26324_ spi0.data_packed\[60\] spi0.data_packed\[61\] net699 VGND VGND VPWR VPWR
+ _05394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20748_ _11408_ _12491_ _12590_ _12595_ VGND VGND VPWR VPWR _12597_ sky130_fd_sc_hd__and4_1
X_23536_ net985 top0.matmul0.a\[8\] _02926_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26255_ _05359_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__clkbuf_1
X_23467_ net1010 top0.matmul0.sin\[3\] _05461_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20679_ _12525_ _12527_ net274 VGND VGND VPWR VPWR _12528_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13220_ top0.pid_d.state\[0\] top0.pid_d.iterate_enable net1019 VGND VGND VPWR VPWR
+ _05445_ sky130_fd_sc_hd__and3_1
X_25206_ _04544_ _04552_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__xnor2_2
X_22418_ net93 _01973_ _01974_ _01975_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__o211a_1
X_23398_ _02835_ _02837_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__xor2_2
X_26186_ spi0.data_packed\[9\] spi0.data_packed\[10\] _05314_ VGND VGND VPWR VPWR
+ _05321_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25137_ _03280_ _04097_ _03123_ _03981_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22349_ _01852_ _01907_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25068_ _03765_ _04414_ _04416_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__a21o_1
X_24019_ _03350_ _03376_ VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__xnor2_1
X_16910_ top0.currT_r\[6\] _08959_ _08960_ VGND VGND VPWR VPWR _08970_ sky130_fd_sc_hd__o21ba_1
X_17890_ _09795_ _09875_ _09876_ VGND VGND VPWR VPWR _09877_ sky130_fd_sc_hd__a21oi_2
X_16841_ top0.currT_r\[2\] _08900_ _08904_ VGND VGND VPWR VPWR _08906_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout680 net681 VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__clkbuf_4
X_19560_ net188 _11446_ _11448_ VGND VGND VPWR VPWR _11449_ sky130_fd_sc_hd__a21o_1
Xfanout691 net692 VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__clkbuf_2
X_16772_ net15 _08854_ VGND VGND VPWR VPWR _08855_ sky130_fd_sc_hd__nor2_4
X_13984_ _06189_ _06196_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__xnor2_1
X_18511_ _10394_ _10397_ _10364_ VGND VGND VPWR VPWR _10491_ sky130_fd_sc_hd__a21o_1
X_15723_ net496 net499 VGND VGND VPWR VPWR _07820_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19491_ top0.pid_d.curr_int\[12\] top0.pid_d.prev_int\[12\] _11383_ VGND VGND VPWR
+ VPWR _11384_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18442_ _10344_ _10422_ VGND VGND VPWR VPWR _10423_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_197_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15654_ net448 net538 VGND VGND VPWR VPWR _07752_ sky130_fd_sc_hd__nand2_1
XFILLER_0_185_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14605_ _06740_ _06742_ VGND VGND VPWR VPWR _06810_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_200_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18373_ net396 net314 VGND VGND VPWR VPWR _10354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15585_ _07679_ _07681_ _07682_ _07683_ _07585_ VGND VGND VPWR VPWR _07684_ sky130_fd_sc_hd__o32a_1
XFILLER_0_185_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17324_ _09315_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__clkbuf_1
X_14536_ _06652_ _06614_ _06659_ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_154_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17255_ _09256_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__clkbuf_1
X_14467_ _06674_ VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16206_ _08207_ _08209_ _08297_ VGND VGND VPWR VPWR _08298_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13418_ _05621_ _05622_ _05619_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__a21o_1
X_17186_ _09195_ _09196_ VGND VGND VPWR VPWR _09197_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14398_ _06535_ _06532_ _06606_ VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_180_Right_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16137_ _08225_ _08229_ VGND VGND VPWR VPWR _08230_ sky130_fd_sc_hd__xor2_1
X_13349_ net47 _05523_ _05524_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16068_ _08153_ _08155_ VGND VGND VPWR VPWR _08161_ sky130_fd_sc_hd__nand2_1
X_15019_ spi0.data_packed\[15\] net1006 _07125_ VGND VGND VPWR VPWR _07135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19827_ net251 _11695_ _11696_ VGND VGND VPWR VPWR _11706_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19758_ _11616_ _11617_ VGND VGND VPWR VPWR _11641_ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18709_ _10671_ _10673_ _10685_ VGND VGND VPWR VPWR _10686_ sky130_fd_sc_hd__a21o_1
X_19689_ net88 net83 net203 VGND VGND VPWR VPWR _11575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21720_ _01155_ _01123_ net142 _01280_ _01266_ net153 VGND VGND VPWR VPWR _01282_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_182_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21651_ net109 VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_177_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_176_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20602_ net302 _12057_ _12448_ net298 _12450_ VGND VGND VPWR VPWR _12451_ sky130_fd_sc_hd__o221a_1
XFILLER_0_192_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24370_ _03207_ _03208_ _03093_ _03094_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__o22a_1
X_21582_ net109 _01143_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_163_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23321_ _11784_ _02765_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_96_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20533_ _12378_ _12379_ _12380_ VGND VGND VPWR VPWR _12382_ sky130_fd_sc_hd__and3_1
XFILLER_0_172_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23252_ net155 _02700_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__or2_1
X_26040_ _05231_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20464_ _12306_ _12312_ VGND VGND VPWR VPWR _12313_ sky130_fd_sc_hd__or2b_1
XFILLER_0_171_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22203_ _01758_ _01763_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__xnor2_2
X_23183_ _02646_ _06380_ _02649_ net831 VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20395_ _12172_ _12173_ _12243_ VGND VGND VPWR VPWR _12244_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22134_ _01210_ _01227_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22065_ _01621_ _01622_ _01558_ _01557_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__a211o_1
X_26942_ clknet_leaf_6_clk_sys _00559_ net594 VGND VGND VPWR VPWR top0.matmul0.a\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_21016_ _12775_ _12780_ _12862_ VGND VGND VPWR VPWR _12863_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26873_ clknet_leaf_37_clk_sys _00490_ net679 VGND VGND VPWR VPWR top0.svm0.tA\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_25824_ _05045_ _05048_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_73_clk_sys clknet_3_5__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_73_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25755_ net767 _04925_ _04998_ VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__a21o_1
XFILLER_0_202_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22967_ _02324_ _02297_ _02475_ _02477_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_179_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24706_ _04058_ _03965_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__or2b_1
X_21918_ _01468_ _01479_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__nor2_1
X_25686_ top0.matmul0.sin\[12\] _04951_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__or2_1
X_22898_ top0.svm0.tC\[5\] _02415_ _02331_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__o21a_1
XFILLER_0_167_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24637_ _03970_ _03971_ _03990_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__a21o_1
X_21849_ net141 net122 VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__and2b_1
XFILLER_0_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15370_ net479 _07468_ VGND VGND VPWR VPWR _07469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24568_ _03795_ _03796_ _03812_ _03798_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__a31o_1
X_14321_ _06487_ _06530_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__xor2_1
XFILLER_0_81_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26307_ _05385_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23519_ top0.a_in_matmul\[0\] top0.matmul0.a\[0\] _02915_ VGND VGND VPWR VPWR _02925_
+ sky130_fd_sc_hd__mux2_1
X_27287_ clknet_3_3__leaf_clk_mosi _00901_ VGND VGND VPWR VPWR spi0.data_packed\[73\]
+ sky130_fd_sc_hd__dfxtp_1
X_24499_ _03846_ _03854_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__xnor2_1
X_17040_ top0.pid_q.prev_error\[15\] top0.pid_q.curr_error\[15\] VGND VGND VPWR VPWR
+ _09092_ sky130_fd_sc_hd__xnor2_1
X_14252_ _06461_ _06459_ _06460_ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__and3_1
X_26238_ spi0.data_packed\[17\] spi0.data_packed\[18\] net697 VGND VGND VPWR VPWR
+ _05351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13203_ net744 top0.ready state\[0\] _05425_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__a22o_1
X_14183_ net45 _05625_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26169_ spi0.data_packed\[7\] _05307_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18991_ net307 _10964_ VGND VGND VPWR VPWR _10965_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17942_ _09925_ _09927_ VGND VGND VPWR VPWR _09928_ sky130_fd_sc_hd__xnor2_1
X_17873_ _09764_ _09761_ _09765_ VGND VGND VPWR VPWR _09860_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16824_ _08861_ VGND VGND VPWR VPWR _08890_ sky130_fd_sc_hd__buf_2
X_19612_ _11497_ _11498_ _11500_ _11468_ VGND VGND VPWR VPWR _11501_ sky130_fd_sc_hd__o22a_1
X_19543_ net176 VGND VGND VPWR VPWR _11433_ sky130_fd_sc_hd__inv_2
X_16755_ _08799_ _08838_ VGND VGND VPWR VPWR _08839_ sky130_fd_sc_hd__xnor2_1
X_13967_ _06103_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15706_ top0.pid_q.out\[1\] top0.pid_q.curr_int\[1\] VGND VGND VPWR VPWR _07803_
+ sky130_fd_sc_hd__or2_1
X_19474_ top0.pid_d.curr_int\[11\] top0.pid_d.prev_int\[11\] VGND VGND VPWR VPWR _11369_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16686_ _08700_ _08705_ _08770_ VGND VGND VPWR VPWR _08771_ sky130_fd_sc_hd__o21a_1
XFILLER_0_159_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13898_ _05756_ _05757_ _06110_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18425_ _10404_ _10405_ net411 VGND VGND VPWR VPWR _10406_ sky130_fd_sc_hd__mux2_1
X_15637_ _07623_ _07628_ _07621_ VGND VGND VPWR VPWR _07735_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18356_ top0.pid_d.curr_int\[5\] VGND VGND VPWR VPWR _10337_ sky130_fd_sc_hd__inv_2
XFILLER_0_185_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15568_ _07540_ _07666_ net514 VGND VGND VPWR VPWR _07667_ sky130_fd_sc_hd__o21ai_2
X_17307_ top0.matmul0.matmul_stage_inst.mult1\[9\] top0.matmul0.matmul_stage_inst.mult2\[9\]
+ VGND VGND VPWR VPWR _09301_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14519_ _06723_ _06725_ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__xor2_1
X_18287_ _10266_ _10268_ VGND VGND VPWR VPWR _10269_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15499_ _07544_ _07597_ VGND VGND VPWR VPWR _07598_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17238_ net551 _09077_ _09135_ VGND VGND VPWR VPWR _09243_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17169_ net553 _09180_ _09181_ _08968_ VGND VGND VPWR VPWR _09182_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20180_ net205 net208 VGND VGND VPWR VPWR _12030_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_110_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23870_ _03225_ _03226_ _03168_ _03169_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22821_ _02339_ top0.svm0.tA\[3\] VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25540_ top0.matmul0.b\[9\] top0.matmul0.matmul_stage_inst.f\[9\] _04856_ VGND VGND
+ VPWR VPWR _04857_ sky130_fd_sc_hd__mux2_1
X_22752_ _02291_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21703_ net146 _01081_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__nor2_2
X_25471_ _04721_ _04750_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22683_ top0.cordic0.sin\[10\] _12004_ _12036_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__and3_1
XFILLER_0_164_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27210_ clknet_leaf_93_clk_sys _00824_ net591 VGND VGND VPWR VPWR top0.cordic0.slte0.opB\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24422_ _03703_ _03704_ _03705_ _03706_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__a211o_1
X_21634_ _01087_ _01172_ _01195_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_165_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27141_ clknet_leaf_13_clk_sys _00755_ net616 VGND VGND VPWR VPWR top0.b_in_matmul\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_24353_ _02998_ _03000_ _03069_ _03071_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21565_ _01121_ _01126_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__xor2_1
XFILLER_0_173_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20516_ _12280_ _12361_ VGND VGND VPWR VPWR _12365_ sky130_fd_sc_hd__nand2_1
X_23304_ _11573_ net215 _11613_ _02687_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__o22a_1
X_24284_ _03146_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__clkbuf_4
X_27072_ clknet_leaf_2_clk_sys _00689_ net582 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.c\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_21496_ net761 _12813_ _01059_ _12963_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26023_ _05218_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__clkbuf_1
X_23235_ _01267_ _02660_ _02679_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__or3_1
XFILLER_0_166_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20447_ _12102_ _12267_ VGND VGND VPWR VPWR _12296_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23166_ _02641_ _06612_ _02645_ net883 VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__a22o_1
X_20378_ _12223_ _12226_ VGND VGND VPWR VPWR _12227_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22117_ _01452_ _01547_ _01638_ _01668_ _01678_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__a311o_1
XFILLER_0_98_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23097_ net171 _02306_ _02594_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__and3_2
X_22048_ _01591_ _01605_ _01609_ _01363_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__o22a_1
X_26925_ clknet_leaf_5_clk_sys _00542_ net598 VGND VGND VPWR VPWR top0.matmul0.cos\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_26856_ clknet_leaf_36_clk_sys _00473_ net686 VGND VGND VPWR VPWR top0.svm0.rising
+ sky130_fd_sc_hd__dfstp_1
X_14870_ spi0.data_packed\[75\] top0.kpd\[11\] _07053_ VGND VGND VPWR VPWR _07055_
+ sky130_fd_sc_hd__mux2_1
X_25807_ top0.matmul0.alpha_pass\[1\] top0.matmul0.beta_pass\[1\] VGND VGND VPWR VPWR
+ _05034_ sky130_fd_sc_hd__nand2_1
X_13821_ _06030_ _06032_ _06033_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26787_ clknet_leaf_3_clk_sys _00404_ net583 VGND VGND VPWR VPWR top0.cordic0.sin\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23999_ _03355_ _03216_ _03356_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16540_ _08620_ _08623_ _08626_ VGND VGND VPWR VPWR _08627_ sky130_fd_sc_hd__mux2_1
X_13752_ _05607_ _05534_ _05587_ net67 VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25738_ top0.matmul0.sin\[13\] _04989_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16471_ _08501_ _08503_ _08502_ VGND VGND VPWR VPWR _08559_ sky130_fd_sc_hd__o21a_1
XFILLER_0_195_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13683_ net50 net47 _05682_ _05894_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__and4_1
X_25669_ top0.matmul0.sin\[7\] top0.matmul0.sin\[8\] _04931_ VGND VGND VPWR VPWR _04941_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18210_ _10098_ _10100_ _10099_ VGND VGND VPWR VPWR _10193_ sky130_fd_sc_hd__o21a_1
XFILLER_0_70_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15422_ _07380_ _07381_ _07376_ VGND VGND VPWR VPWR _07521_ sky130_fd_sc_hd__nand3_1
X_19190_ _11120_ _11140_ _11141_ VGND VGND VPWR VPWR _11142_ sky130_fd_sc_hd__and3_1
XFILLER_0_167_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18141_ _10119_ _10124_ VGND VGND VPWR VPWR _10125_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15353_ _07442_ _07451_ _07449_ VGND VGND VPWR VPWR _07452_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14304_ net23 _06025_ VGND VGND VPWR VPWR _06514_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18072_ _10054_ _10056_ VGND VGND VPWR VPWR _10057_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15284_ _07233_ _07374_ _07322_ net487 VGND VGND VPWR VPWR _07383_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17023_ _09074_ _09075_ VGND VGND VPWR VPWR _09076_ sky130_fd_sc_hd__or2b_1
XFILLER_0_124_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14235_ _06433_ _06434_ _06444_ _06445_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_34_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14166_ _06256_ _06376_ _06377_ VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14097_ _06307_ _06308_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__xnor2_1
X_18974_ net356 _10947_ net363 VGND VGND VPWR VPWR _10948_ sky130_fd_sc_hd__o21ai_1
X_17925_ net325 net408 VGND VGND VPWR VPWR _09911_ sky130_fd_sc_hd__nand2_1
X_17856_ _09841_ _09842_ VGND VGND VPWR VPWR _09843_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16807_ top0.kiq\[13\] _05448_ _08854_ VGND VGND VPWR VPWR _08877_ sky130_fd_sc_hd__and3_1
X_17787_ _09770_ _09773_ VGND VGND VPWR VPWR _09774_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14999_ _07124_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16738_ net447 _07781_ VGND VGND VPWR VPWR _08822_ sky130_fd_sc_hd__and2_1
X_19526_ net123 net120 net1031 net113 net197 net191 VGND VGND VPWR VPWR _11416_ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19457_ top0.pid_d.curr_int\[9\] top0.pid_d.prev_int\[9\] VGND VGND VPWR VPWR _11354_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16669_ _08527_ _08753_ VGND VGND VPWR VPWR _08754_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_147_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18408_ net341 _10386_ _10388_ VGND VGND VPWR VPWR _10389_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19388_ top0.pid_d.curr_int\[0\] top0.pid_d.prev_int\[0\] VGND VGND VPWR VPWR _11294_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_91_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18339_ _10225_ _10230_ _10320_ VGND VGND VPWR VPWR _10321_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_clk_sys clknet_3_2__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_21_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_173_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21350_ _13141_ _13146_ VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20301_ _12133_ _12148_ _12149_ VGND VGND VPWR VPWR _12150_ sky130_fd_sc_hd__nand3_2
XFILLER_0_130_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21281_ net214 _12853_ VGND VGND VPWR VPWR _13124_ sky130_fd_sc_hd__xnor2_2
Xfanout4 _05518_ VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__buf_4
X_23020_ top0.svm0.delta\[14\] _02522_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__xor2_1
X_20232_ _12051_ _12046_ _12080_ _12043_ VGND VGND VPWR VPWR _12081_ sky130_fd_sc_hd__and4b_1
XFILLER_0_4_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20163_ net205 net208 VGND VGND VPWR VPWR _12015_ sky130_fd_sc_hd__and2b_1
XFILLER_0_110_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_200_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24971_ _04315_ _04321_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__xnor2_1
X_20094_ _11433_ VGND VGND VPWR VPWR _11954_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26710_ clknet_leaf_71_clk_sys _00327_ net657 VGND VGND VPWR VPWR top0.pid_d.curr_int\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_23922_ _03029_ _03030_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_179_Left_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26641_ clknet_leaf_80_clk_sys _00258_ net634 VGND VGND VPWR VPWR top0.pid_d.out\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_23853_ _03004_ _03005_ _03069_ _03071_ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22804_ top0.svm0.counter\[6\] VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__inv_2
X_26572_ clknet_leaf_54_clk_sys _00195_ net667 VGND VGND VPWR VPWR top0.pid_q.curr_error\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_23784_ _03049_ _03050_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__nor2_1
X_20996_ _12778_ _12836_ _12840_ net284 _12842_ VGND VGND VPWR VPWR _12843_ sky130_fd_sc_hd__a221o_2
XFILLER_0_79_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25523_ top0.matmul0.b\[1\] top0.matmul0.matmul_stage_inst.f\[1\] _04846_ VGND VGND
+ VPWR VPWR _04848_ sky130_fd_sc_hd__mux2_1
X_22735_ _08900_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25454_ _04737_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22666_ _01211_ _02216_ _02217_ _01230_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24405_ _02994_ _02996_ _03024_ _03025_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__o22a_1
X_21617_ net152 _01178_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__or2_1
X_25385_ _03889_ _04677_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_188_Left_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22597_ _02147_ _02150_ net98 VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__o21a_1
X_27124_ clknet_leaf_33_clk_sys _00738_ net665 VGND VGND VPWR VPWR top0.c_out_calc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_24336_ _03686_ _03692_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21548_ _01101_ _01109_ VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27055_ clknet_leaf_20_clk_sys _00672_ net609 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.d\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24267_ net8 _03447_ _03434_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_65_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21479_ _12963_ _01042_ _01043_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14020_ _06226_ _06232_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__xnor2_2
X_26006_ top0.b_in_matmul\[10\] _05205_ _05196_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23218_ _11425_ _02667_ _02668_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__a21bo_2
X_24198_ _03505_ _03508_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23149_ top0.svm0.delta\[14\] _02632_ _02595_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15971_ _07969_ _07973_ _08065_ VGND VGND VPWR VPWR _08066_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17710_ _09475_ _09478_ _09472_ VGND VGND VPWR VPWR _09697_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_41_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14922_ spi0.data_packed\[36\] top0.kid\[4\] _07075_ VGND VGND VPWR VPWR _07082_
+ sky130_fd_sc_hd__mux2_1
X_26908_ clknet_leaf_109_clk_sys _00525_ net579 VGND VGND VPWR VPWR top0.matmul0.sin\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_18690_ _10657_ _10665_ VGND VGND VPWR VPWR _10668_ sky130_fd_sc_hd__nor2_1
XFILLER_0_175_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold60 top0.pid_d.curr_error\[11\] VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 top0.cordic0.cos\[8\] VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 top0.periodTop\[3\] VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17641_ net412 net419 net330 net337 VGND VGND VPWR VPWR _09628_ sky130_fd_sc_hd__and4_1
X_26839_ clknet_leaf_47_clk_sys _00456_ net680 VGND VGND VPWR VPWR top0.svm0.counter\[14\]
+ sky130_fd_sc_hd__dfrtp_2
X_14853_ spi0.data_packed\[67\] top0.kpd\[3\] _07042_ VGND VGND VPWR VPWR _07046_
+ sky130_fd_sc_hd__mux2_1
Xhold93 top0.kpq\[5\] VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13804_ _05995_ _06015_ _06016_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__a21bo_1
X_17572_ net415 net410 VGND VGND VPWR VPWR _09559_ sky130_fd_sc_hd__or2b_1
X_14784_ _06952_ _06983_ _06984_ VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_58_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19311_ net437 _11251_ VGND VGND VPWR VPWR _11252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16523_ top0.pid_q.out\[11\] _07704_ VGND VGND VPWR VPWR _08611_ sky130_fd_sc_hd__nor2_1
X_13735_ _05924_ _05926_ _05947_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19242_ net440 _11187_ _11188_ VGND VGND VPWR VPWR _11189_ sky130_fd_sc_hd__and3_1
XFILLER_0_195_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16454_ _08542_ VGND VGND VPWR VPWR _08543_ sky130_fd_sc_hd__inv_2
XFILLER_0_183_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13666_ _05863_ _05874_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15405_ net537 net486 _07503_ net481 VGND VGND VPWR VPWR _07504_ sky130_fd_sc_hd__a31o_1
X_19173_ top0.pid_d.prev_error\[1\] top0.pid_d.curr_error\[1\] VGND VGND VPWR VPWR
+ _11126_ sky130_fd_sc_hd__xnor2_1
X_16385_ _08388_ VGND VGND VPWR VPWR _08475_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_183_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13597_ net63 _05551_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__nand2_1
X_18124_ net325 net398 VGND VGND VPWR VPWR _10108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15336_ _07414_ _07433_ VGND VGND VPWR VPWR _07435_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18055_ _09931_ _09957_ _09958_ VGND VGND VPWR VPWR _10040_ sky130_fd_sc_hd__o21ai_1
X_15267_ net484 VGND VGND VPWR VPWR _07366_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_2 _01211_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17006_ top0.matmul0.beta_pass\[13\] _05437_ VGND VGND VPWR VPWR _09060_ sky130_fd_sc_hd__nand2_1
X_14218_ _05688_ _05822_ _06308_ _06307_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__o31a_1
XFILLER_0_1_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15198_ _07293_ _07296_ VGND VGND VPWR VPWR _07297_ sky130_fd_sc_hd__xor2_2
XFILLER_0_22_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14149_ _06155_ _06247_ VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__nand2_1
Xfanout509 net510 VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__buf_2
XFILLER_0_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18957_ _10880_ _10886_ VGND VGND VPWR VPWR _10931_ sky130_fd_sc_hd__xor2_1
X_17908_ top0.pid_d.curr_int\[0\] VGND VGND VPWR VPWR _09895_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18888_ _09395_ _10778_ _10862_ VGND VGND VPWR VPWR _10863_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_174_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17839_ _09809_ _09824_ _09825_ VGND VGND VPWR VPWR _09826_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_178_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20850_ net238 net234 VGND VGND VPWR VPWR _12699_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_7_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19509_ top0.pid_d.curr_int\[14\] top0.pid_d.prev_int\[14\] _11393_ VGND VGND VPWR
+ VPWR _11400_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20781_ _12344_ _12623_ _11438_ VGND VGND VPWR VPWR _12630_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22520_ _02073_ _02075_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22451_ _01979_ _01982_ _01978_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21402_ net232 _11759_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__nand2_1
X_25170_ _04039_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22382_ _01934_ _01940_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24121_ _03393_ _03397_ _03406_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21333_ _12819_ _13174_ top0.cordic0.vec\[0\]\[10\] VGND VGND VPWR VPWR _13175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_170_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24052_ _03384_ _03402_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_130_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21264_ _12740_ _13107_ VGND VGND VPWR VPWR _13108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23003_ top0.svm0.delta\[11\] VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__inv_2
X_20215_ _12062_ _12063_ VGND VGND VPWR VPWR _12064_ sky130_fd_sc_hd__and2b_1
XFILLER_0_40_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21195_ _13033_ _13038_ VGND VGND VPWR VPWR _13039_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20146_ net212 _11936_ _11978_ VGND VGND VPWR VPWR _12001_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24954_ _04212_ _04233_ _04304_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__a21o_1
X_20077_ net203 net187 VGND VGND VPWR VPWR _11938_ sky130_fd_sc_hd__xnor2_1
X_23905_ _03237_ _03242_ _03261_ _03262_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__a211o_1
X_24885_ _04170_ _04236_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__xnor2_2
X_26624_ clknet_leaf_29_clk_sys _00241_ net624 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_135_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23836_ _03192_ _03175_ _03176_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__nand3_2
XFILLER_0_197_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26555_ clknet_leaf_49_clk_sys _00178_ net675 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23767_ _03120_ _03121_ _03123_ _03124_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__and4_2
X_20979_ net225 net222 VGND VGND VPWR VPWR _12826_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25506_ top0.matmul0.matmul_stage_inst.mult1\[9\] _04470_ _04829_ VGND VGND VPWR
+ VPWR _04839_ sky130_fd_sc_hd__mux2_1
X_13520_ net1025 _05656_ _05639_ _05624_ net60 VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__a32o_1
X_22718_ _02257_ _02268_ VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__xnor2_1
X_26486_ clknet_leaf_62_clk_sys _00018_ net647 VGND VGND VPWR VPWR top0.pid_q.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_23698_ _03054_ _03055_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__or2_2
XFILLER_0_137_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_192_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25437_ _04776_ _04779_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__xor2_1
X_13451_ top0.matmul0.alpha_pass\[13\] _05435_ _05474_ _05464_ top0.c_out_calc\[13\]
+ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22649_ _02201_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__inv_2
XFILLER_0_192_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16170_ net456 net1029 VGND VGND VPWR VPWR _08262_ sky130_fd_sc_hd__nand2_2
X_25368_ _04406_ _04698_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__nor2_2
X_13382_ _05512_ _05516_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27107_ clknet_leaf_11_clk_sys _00724_ net601 VGND VGND VPWR VPWR top0.matmul0.op\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15121_ _07219_ VGND VGND VPWR VPWR _07220_ sky130_fd_sc_hd__clkbuf_2
X_24319_ _03664_ _03671_ _03675_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_23_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25299_ _04638_ _04644_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15052_ net528 net475 VGND VGND VPWR VPWR _07151_ sky130_fd_sc_hd__nand2_1
X_27038_ clknet_leaf_7_clk_sys _00655_ net593 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_181_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput4 net4 VGND VGND VPWR VPWR pwmA sky130_fd_sc_hd__clkbuf_4
X_14003_ _05567_ _05757_ net24 VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__o21bai_1
X_19860_ _11430_ _11736_ VGND VGND VPWR VPWR _11737_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18811_ _10786_ VGND VGND VPWR VPWR _10787_ sky130_fd_sc_hd__inv_2
X_19791_ net253 VGND VGND VPWR VPWR _11672_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15954_ net499 _08048_ VGND VGND VPWR VPWR _08049_ sky130_fd_sc_hd__nand2_4
X_18742_ net334 net338 net331 VGND VGND VPWR VPWR _10719_ sky130_fd_sc_hd__o21a_1
X_14905_ spi0.data_packed\[60\] top0.kpq\[12\] _07064_ VGND VGND VPWR VPWR _07073_
+ sky130_fd_sc_hd__mux2_1
X_18673_ _10550_ _10553_ _10650_ VGND VGND VPWR VPWR _10651_ sky130_fd_sc_hd__a21o_1
X_15885_ _07980_ _07880_ VGND VGND VPWR VPWR _07981_ sky130_fd_sc_hd__nand2_1
X_14836_ net824 _06279_ _07034_ _05465_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__a22o_1
X_17624_ net420 net426 _09610_ net1022 VGND VGND VPWR VPWR _09611_ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_176_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17555_ _09540_ _09541_ VGND VGND VPWR VPWR _09542_ sky130_fd_sc_hd__nor2_1
X_14767_ _06935_ _06968_ VGND VGND VPWR VPWR _06969_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16506_ _08312_ _08535_ VGND VGND VPWR VPWR _08594_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13718_ _05929_ _05930_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__xnor2_1
X_17486_ net408 net403 net343 net347 VGND VGND VPWR VPWR _09473_ sky130_fd_sc_hd__and4_1
X_14698_ _06870_ _06901_ VGND VGND VPWR VPWR _06902_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_184_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16437_ net498 _08447_ VGND VGND VPWR VPWR _08526_ sky130_fd_sc_hd__nand2_2
X_19225_ top0.pid_d.curr_error\[5\] VGND VGND VPWR VPWR _11173_ sky130_fd_sc_hd__inv_2
X_13649_ net66 _05605_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__nand2_1
XFILLER_0_171_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19156_ net374 _11095_ _11113_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__a21o_1
X_16368_ _08456_ _08457_ VGND VGND VPWR VPWR _08458_ sky130_fd_sc_hd__or2b_1
XFILLER_0_54_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_200_Left_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18107_ _09990_ _09999_ _09998_ VGND VGND VPWR VPWR _10091_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15319_ _07415_ _07417_ VGND VGND VPWR VPWR _07418_ sky130_fd_sc_hd__nand2_1
X_19087_ net311 _11057_ _11058_ VGND VGND VPWR VPWR _11059_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16299_ _08334_ _08389_ VGND VGND VPWR VPWR _08390_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18038_ _09909_ _09914_ _09907_ VGND VGND VPWR VPWR _10023_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout306 top0.cordic0.vec\[0\]\[0\] VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkbuf_4
X_20000_ _11852_ _11854_ _11866_ VGND VGND VPWR VPWR _11867_ sky130_fd_sc_hd__a21o_1
XFILLER_0_185_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout317 net318 VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__buf_2
Xfanout328 net329 VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_2
Xfanout339 top0.pid_d.mult0.b\[5\] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__buf_4
X_19989_ _11783_ VGND VGND VPWR VPWR _11857_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21951_ net166 _01123_ _01512_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20902_ _12711_ _12712_ VGND VGND VPWR VPWR _12750_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24670_ _04022_ _04023_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__xor2_1
XFILLER_0_55_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21882_ net156 _01440_ _01443_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23621_ net574 top0.matmul0.matmul_stage_inst.d\[8\] top0.matmul0.matmul_stage_inst.c\[8\]
+ net558 VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__a22o_2
X_20833_ net214 _12238_ VGND VGND VPWR VPWR _12682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26340_ spi0.data_packed\[68\] spi0.data_packed\[69\] net692 VGND VGND VPWR VPWR
+ _05402_ sky130_fd_sc_hd__mux2_1
X_23552_ _02942_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_194_Right_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20764_ _11438_ net292 VGND VGND VPWR VPWR _12613_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22503_ _02056_ _02058_ _01408_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__a21oi_1
X_26271_ _05367_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__clkbuf_1
X_20695_ _12531_ _12532_ _12515_ VGND VGND VPWR VPWR _12544_ sky130_fd_sc_hd__a21oi_1
X_23483_ _02906_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25222_ _04492_ _04504_ _04490_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_162_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22434_ _01990_ _01991_ _01896_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25153_ _04498_ _04500_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22365_ _01820_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__buf_4
XFILLER_0_143_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24104_ _03389_ _03390_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__xor2_2
X_21316_ _13112_ _13134_ _13036_ VGND VGND VPWR VPWR _13158_ sky130_fd_sc_hd__o21a_1
X_25084_ _04427_ _04432_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__xnor2_1
X_22296_ _01843_ _01855_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24035_ _03387_ _03392_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21247_ _12533_ _12665_ VGND VGND VPWR VPWR _13091_ sky130_fd_sc_hd__or2_1
X_21178_ _12134_ _12985_ _13019_ net252 _13021_ VGND VGND VPWR VPWR _13022_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20129_ net212 _11947_ VGND VGND VPWR VPWR _11985_ sky130_fd_sc_hd__nand2_1
X_25986_ net966 _05189_ _05165_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24937_ _03164_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15670_ _07366_ _07558_ _07559_ VGND VGND VPWR VPWR _07768_ sky130_fd_sc_hd__a21oi_1
X_24868_ _02985_ _02987_ _03741_ _03742_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__o22a_1
XFILLER_0_169_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14621_ _06768_ _06769_ _06825_ VGND VGND VPWR VPWR _06826_ sky130_fd_sc_hd__o21a_1
X_26607_ clknet_leaf_82_clk_sys _00002_ net637 VGND VGND VPWR VPWR top0.pid_d.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23819_ _02976_ _02977_ _03024_ _03025_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__o22a_2
X_24799_ _04141_ _04151_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_197_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17340_ _09323_ _09327_ _09328_ VGND VGND VPWR VPWR _09329_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14552_ _06753_ _06757_ VGND VGND VPWR VPWR _06758_ sky130_fd_sc_hd__xnor2_4
X_26538_ clknet_leaf_60_clk_sys _00161_ net653 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_161_Right_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13503_ _05649_ _05651_ _05715_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17271_ top0.matmul0.matmul_stage_inst.mult2\[3\] _09265_ _09269_ VGND VGND VPWR
+ VPWR _09270_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_138_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14483_ _06547_ _06550_ _06689_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__a21o_1
X_26469_ clknet_leaf_45_clk_sys _00100_ net681 VGND VGND VPWR VPWR top0.svm0.delta\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_138_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19010_ _10982_ _10983_ VGND VGND VPWR VPWR _10984_ sky130_fd_sc_hd__xnor2_1
X_16222_ _08311_ _08313_ VGND VGND VPWR VPWR _08314_ sky130_fd_sc_hd__xnor2_1
X_13434_ _05636_ _05646_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_68_clk_sys clknet_3_5__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_68_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_109_clk_sys clknet_3_2__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_109_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_16153_ _08243_ _08239_ _08244_ VGND VGND VPWR VPWR _08245_ sky130_fd_sc_hd__a21o_1
X_13365_ _05564_ _05570_ _05577_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15104_ _07156_ _07157_ _07202_ VGND VGND VPWR VPWR _07203_ sky130_fd_sc_hd__a21bo_1
X_16084_ _08123_ _08128_ _08049_ VGND VGND VPWR VPWR _08177_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13296_ _05482_ _05508_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19912_ net224 _11785_ VGND VGND VPWR VPWR _11786_ sky130_fd_sc_hd__nor2_1
X_15035_ top0.pid_d.prev_int\[5\] _07140_ _07144_ top0.pid_d.curr_int\[5\] VGND VGND
+ VPWR VPWR _00122_ sky130_fd_sc_hd__a22o_1
X_19843_ _11718_ _11720_ VGND VGND VPWR VPWR _11721_ sky130_fd_sc_hd__xnor2_2
X_19774_ net194 net190 VGND VGND VPWR VPWR _11656_ sky130_fd_sc_hd__or2_1
X_16986_ top0.matmul0.beta_pass\[12\] _09040_ VGND VGND VPWR VPWR _09041_ sky130_fd_sc_hd__xor2_1
X_18725_ _10456_ _10644_ VGND VGND VPWR VPWR _10702_ sky130_fd_sc_hd__and2b_1
X_15937_ _07938_ _07940_ _07939_ VGND VGND VPWR VPWR _08032_ sky130_fd_sc_hd__o21a_1
XFILLER_0_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire16 net17 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
X_18656_ _10537_ _10539_ _10538_ VGND VGND VPWR VPWR _10634_ sky130_fd_sc_hd__o21ai_1
X_15868_ _07928_ _07963_ VGND VGND VPWR VPWR _07964_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14819_ _07013_ _07018_ VGND VGND VPWR VPWR _07019_ sky130_fd_sc_hd__or2b_1
X_17607_ _09567_ _09593_ _09364_ _09559_ VGND VGND VPWR VPWR _09594_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18587_ net402 _10564_ _10565_ VGND VGND VPWR VPWR _10566_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15799_ net549 _07699_ _07895_ VGND VGND VPWR VPWR _07896_ sky130_fd_sc_hd__and3_1
XFILLER_0_171_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17538_ net418 net349 VGND VGND VPWR VPWR _09525_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_188_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17469_ _09427_ _09450_ _09452_ _09455_ VGND VGND VPWR VPWR _09456_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_50_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19208_ _11156_ _11157_ VGND VGND VPWR VPWR _11158_ sky130_fd_sc_hd__xnor2_1
X_20480_ _12059_ _12326_ _12328_ net287 VGND VGND VPWR VPWR _12329_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19139_ top0.kid\[4\] _11098_ _11100_ top0.kpd\[4\] VGND VGND VPWR VPWR _11105_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22150_ net99 _01223_ _01211_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21101_ _12875_ _12945_ _12946_ VGND VGND VPWR VPWR _12947_ sky130_fd_sc_hd__o21a_1
XFILLER_0_140_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22081_ _01066_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21032_ _12804_ _12805_ VGND VGND VPWR VPWR _12879_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout103 top0.cordic0.vec\[1\]\[13\] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout114 net116 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__buf_4
XFILLER_0_61_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout125 top0.cordic0.vec\[1\]\[8\] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__buf_2
Xfanout136 net137 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__buf_2
XFILLER_0_195_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout147 net148 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_4
X_25840_ net743 _05029_ _05031_ _05062_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__a22o_1
Xfanout158 top0.cordic0.vec\[1\]\[1\] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_4
Xfanout169 top0.svm0.counter\[10\] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25771_ net730 _00000_ _05006_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__o21a_1
X_22983_ top0.svm0.delta\[8\] VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__inv_2
X_24722_ _04073_ _04074_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__xnor2_1
X_21934_ net136 net153 VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24653_ _04000_ _04005_ _04006_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_106_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21865_ _01396_ _01426_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__xnor2_1
X_23604_ top0.matmul0.alpha_pass\[9\] _09302_ net559 VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20816_ _12463_ _12664_ VGND VGND VPWR VPWR _12665_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24584_ _03937_ _03938_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21796_ _01266_ net152 VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26323_ _05393_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23535_ _02933_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__clkbuf_1
X_20747_ _12590_ _12595_ net303 _12491_ VGND VGND VPWR VPWR _12596_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_64_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_190_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26254_ spi0.data_packed\[25\] spi0.data_packed\[26\] net698 VGND VGND VPWR VPWR
+ _05359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23466_ _02897_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20678_ net249 _12499_ _12526_ _12493_ VGND VGND VPWR VPWR _12527_ sky130_fd_sc_hd__o211ai_1
X_25205_ _04546_ _04551_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_110_clk_sys clknet_3_2__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_110_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22417_ net80 _01923_ _01925_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__or3b_1
X_26185_ _05320_ VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__clkbuf_1
X_23397_ _11513_ _02836_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25136_ _03200_ _04288_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_115_Left_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22348_ _11674_ _01845_ net87 VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25067_ _04252_ _04258_ _04415_ _04039_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__a31o_1
X_22279_ _01835_ _01838_ _01408_ VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__mux2_2
X_24018_ _03372_ _03374_ _03375_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__a21bo_1
Xhold190 _00319_ VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__dlygate4sd3_1
X_16840_ _08900_ _08904_ top0.currT_r\[2\] VGND VGND VPWR VPWR _08905_ sky130_fd_sc_hd__o21ai_1
Xfanout670 net673 VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__clkbuf_4
Xfanout681 net686 VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__clkbuf_4
X_16771_ _07698_ _08853_ VGND VGND VPWR VPWR _08854_ sky130_fd_sc_hd__nor2_4
Xfanout692 net693 VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__buf_2
X_13983_ _06191_ _06195_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__xnor2_1
X_25969_ top0.matmul0.beta_pass\[2\] _05169_ _05176_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__a21o_1
XFILLER_0_176_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18510_ _10464_ _10489_ VGND VGND VPWR VPWR _10490_ sky130_fd_sc_hd__xnor2_2
X_15722_ _07719_ _07720_ _07818_ VGND VGND VPWR VPWR _07819_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_124_Left_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19490_ top0.pid_d.curr_int\[12\] top0.pid_d.prev_int\[12\] _11379_ VGND VGND VPWR
+ VPWR _11383_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18441_ _10420_ _10421_ VGND VGND VPWR VPWR _10422_ sky130_fd_sc_hd__and2b_1
X_15653_ net540 net446 VGND VGND VPWR VPWR _07751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14604_ _06740_ _06742_ VGND VGND VPWR VPWR _06809_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18372_ net401 net312 VGND VGND VPWR VPWR _10353_ sky130_fd_sc_hd__nand2_1
X_15584_ _07589_ _07592_ _07546_ _07547_ VGND VGND VPWR VPWR _07683_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_0_68_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17323_ top0.matmul0.beta_pass\[11\] _09314_ net562 VGND VGND VPWR VPWR _09315_ sky130_fd_sc_hd__mux2_1
X_14535_ _06656_ _06657_ _06741_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_83_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17254_ top0.matmul0.beta_pass\[1\] _09255_ net563 VGND VGND VPWR VPWR _09256_ sky130_fd_sc_hd__mux2_1
X_14466_ _06553_ _06556_ VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_181_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16205_ _08207_ _08209_ _08205_ VGND VGND VPWR VPWR _08297_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_52_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13417_ _05629_ _05623_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__nor2_1
X_17185_ top0.pid_q.curr_int\[8\] top0.pid_q.prev_int\[8\] VGND VGND VPWR VPWR _09196_
+ sky130_fd_sc_hd__xnor2_1
X_14397_ _06536_ _06530_ _06604_ _06605_ _06540_ VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__a311o_1
XFILLER_0_148_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_133_Left_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16136_ _08227_ _08228_ VGND VGND VPWR VPWR _08229_ sky130_fd_sc_hd__xnor2_1
X_13348_ net50 _05520_ _05521_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16067_ _08160_ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__clkbuf_1
X_13279_ net40 _05489_ _05491_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15018_ _07134_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__clkbuf_1
X_19826_ _11703_ _11704_ VGND VGND VPWR VPWR _11705_ sky130_fd_sc_hd__or2_1
X_19757_ net83 _11631_ _11639_ net180 VGND VGND VPWR VPWR _11640_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_155_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_142_Left_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16969_ top0.pid_q.curr_error\[10\] VGND VGND VPWR VPWR _09025_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18708_ _10671_ _10673_ _10670_ VGND VGND VPWR VPWR _10685_ sky130_fd_sc_hd__o21a_1
X_19688_ net194 _11572_ VGND VGND VPWR VPWR _11574_ sky130_fd_sc_hd__nor2_1
XFILLER_0_182_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_188_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18639_ net387 net311 VGND VGND VPWR VPWR _10617_ sky130_fd_sc_hd__nand2_1
X_21650_ net114 _01211_ _01111_ VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20601_ net298 _12449_ VGND VGND VPWR VPWR _12450_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21581_ net119 net116 VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_191_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23320_ _11649_ _02765_ _11954_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__a21o_1
X_20532_ _12378_ _12379_ _12380_ VGND VGND VPWR VPWR _12381_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_151_Left_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20463_ _12284_ _12301_ _12307_ _12311_ net280 VGND VGND VPWR VPWR _12312_ sky130_fd_sc_hd__a311o_1
X_23251_ _11511_ _02660_ _02677_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_162_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22202_ _01759_ _01760_ _01761_ _01762_ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__a211o_1
X_23182_ _02646_ _06275_ _02649_ net729 VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__a22o_1
X_20394_ _12196_ _12242_ VGND VGND VPWR VPWR _12243_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22133_ _01685_ _01694_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__xor2_2
XFILLER_0_3_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26941_ clknet_leaf_9_clk_sys _00558_ net594 VGND VGND VPWR VPWR top0.matmul0.a\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_22064_ _01557_ _01623_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__nand2_1
XFILLER_0_199_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21015_ _12775_ _12780_ _12760_ VGND VGND VPWR VPWR _12862_ sky130_fd_sc_hd__o21a_1
X_26872_ clknet_leaf_37_clk_sys _00489_ net679 VGND VGND VPWR VPWR top0.svm0.tA\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_160_Left_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25823_ _05046_ _05047_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_16_clk_sys clknet_3_2__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_16_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_8_clk_sys clknet_3_2__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_8_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_25754_ net70 top0.matmul0.cos\[5\] _05458_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__and3_1
X_22966_ _02324_ _02476_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__nor2_1
X_24705_ _03965_ _04058_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__and2b_1
XFILLER_0_167_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21917_ net166 _01471_ _01473_ _01474_ _01478_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__o221a_1
X_25685_ _04913_ _04953_ net841 _00000_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__o2bb2a_1
X_22897_ _02332_ top0.svm0.tC\[4\] _02414_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24636_ _03980_ _03989_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_38_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21848_ net122 net141 VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__and2b_1
XFILLER_0_194_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24567_ _03919_ _03920_ _03915_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__o21ai_2
X_21779_ net130 net129 net121 net113 VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__and4_1
XFILLER_0_33_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14320_ _06510_ _06529_ VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__xnor2_4
X_26306_ spi0.data_packed\[51\] spi0.data_packed\[52\] net697 VGND VGND VPWR VPWR
+ _05385_ sky130_fd_sc_hd__mux2_1
X_23518_ _02924_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27286_ clknet_3_2__leaf_clk_mosi _00900_ VGND VGND VPWR VPWR spi0.data_packed\[72\]
+ sky130_fd_sc_hd__dfxtp_1
X_24498_ _03751_ _03847_ _03848_ _03752_ _03853_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__o221a_1
XFILLER_0_111_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14251_ _06459_ _06460_ _06461_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26237_ _05350_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23449_ net88 _02883_ _02884_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__a21bo_1
X_13202_ top0.pid_d.state\[0\] _05427_ net16 net433 VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14182_ _06344_ _06391_ _06392_ VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26168_ spi0.data_packed\[5\] spi0.data_packed\[6\] _05299_ net18 VGND VGND VPWR
+ VPWR _05307_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25119_ _04405_ _04408_ _04465_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18990_ net374 net371 _10495_ VGND VGND VPWR VPWR _10964_ sky130_fd_sc_hd__and3_1
X_26099_ _12017_ _12019_ _12012_ _12009_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__o22a_2
XFILLER_0_108_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17941_ _09834_ _09835_ _09926_ VGND VGND VPWR VPWR _09927_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_195_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17872_ _09788_ _09805_ _09804_ VGND VGND VPWR VPWR _09859_ sky130_fd_sc_hd__a21oi_1
X_19611_ top0.cordic0.slte0.opA\[10\] _11499_ _11475_ VGND VGND VPWR VPWR _11500_
+ sky130_fd_sc_hd__a21oi_1
X_16823_ _08882_ _08885_ _08887_ _08888_ _08889_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__o311a_1
X_19542_ _11424_ _11431_ net174 VGND VGND VPWR VPWR _11432_ sky130_fd_sc_hd__o21ai_1
X_13966_ _06171_ _06172_ _06174_ _06170_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__o22ai_4
X_16754_ _08806_ _08837_ VGND VGND VPWR VPWR _08838_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15705_ top0.pid_q.out\[0\] top0.pid_q.curr_int\[0\] top0.pid_q.curr_int\[1\] top0.pid_q.out\[1\]
+ VGND VGND VPWR VPWR _07802_ sky130_fd_sc_hd__a22o_1
X_16685_ _08700_ _08705_ _08698_ VGND VGND VPWR VPWR _08770_ sky130_fd_sc_hd__a21o_1
X_19473_ _11366_ _11359_ _11367_ VGND VGND VPWR VPWR _11368_ sky130_fd_sc_hd__o21a_1
X_13897_ _05756_ _05757_ _05758_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_159_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18424_ net310 _10263_ _10403_ VGND VGND VPWR VPWR _10405_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15636_ _07642_ _07646_ _07733_ VGND VGND VPWR VPWR _07734_ sky130_fd_sc_hd__a21o_1
XFILLER_0_185_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_186_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18355_ _10336_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__clkbuf_1
X_15567_ net484 _07274_ _07276_ VGND VGND VPWR VPWR _07666_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14518_ _06622_ _06627_ _06724_ VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__o21a_1
X_17306_ _09298_ _09294_ _09299_ VGND VGND VPWR VPWR _09300_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18286_ _10192_ _10194_ _10267_ VGND VGND VPWR VPWR _10268_ sky130_fd_sc_hd__o21a_1
X_15498_ net517 _07257_ VGND VGND VPWR VPWR _07597_ sky130_fd_sc_hd__nor2_1
X_14449_ net49 _06135_ VGND VGND VPWR VPWR _06657_ sky130_fd_sc_hd__and2_1
X_17237_ top0.pid_q.curr_int\[14\] _09236_ _09241_ net554 VGND VGND VPWR VPWR _09242_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17168_ _09178_ _09179_ VGND VGND VPWR VPWR _09181_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16119_ _08200_ _08211_ VGND VGND VPWR VPWR _08212_ sky130_fd_sc_hd__xor2_1
XFILLER_0_122_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17099_ top0.pid_q.curr_error\[8\] _08860_ _09117_ VGND VGND VPWR VPWR _09126_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19809_ net250 VGND VGND VPWR VPWR _11689_ sky130_fd_sc_hd__clkinv_4
X_22820_ _02339_ top0.svm0.tA\[3\] VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22751_ net549 _07704_ _05443_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__o21a_2
XFILLER_0_79_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21702_ _01151_ _01263_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__xnor2_2
X_25470_ _04717_ _04812_ _04810_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22682_ _02224_ _02233_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24421_ _03775_ _03776_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21633_ _01184_ _01190_ _01194_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27140_ clknet_leaf_14_clk_sys _00754_ net618 VGND VGND VPWR VPWR top0.b_in_matmul\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_24352_ _02989_ _02991_ _03054_ _03055_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__o22a_1
XFILLER_0_142_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21564_ net124 _01089_ _01124_ _01125_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_51_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23303_ net138 _02748_ _02749_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__a21bo_1
X_27071_ clknet_leaf_2_clk_sys _00688_ net582 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.c\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_20515_ _12266_ _12362_ _12363_ VGND VGND VPWR VPWR _12364_ sky130_fd_sc_hd__o21a_1
XFILLER_0_160_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24283_ _03301_ _03640_ VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__xnor2_4
X_21495_ _01057_ _01058_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_166_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26022_ net994 _05217_ _05196_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23234_ _02683_ _02660_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__nand2_1
X_20446_ net264 _12250_ _12294_ _11593_ _12090_ VGND VGND VPWR VPWR _12295_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23165_ _02641_ _06546_ _02645_ net811 VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__a22o_1
X_20377_ net276 _12131_ _12224_ _12225_ VGND VGND VPWR VPWR _12226_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_30_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22116_ _01672_ _01673_ _01676_ _01677_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__or4_1
X_23096_ net555 _02483_ _02596_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22047_ _01318_ _01608_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__nor2_1
X_26924_ clknet_leaf_4_clk_sys _00541_ net580 VGND VGND VPWR VPWR top0.matmul0.cos\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_26855_ clknet_leaf_46_clk_sys _00472_ net680 VGND VGND VPWR VPWR top0.svm0.delta\[15\]
+ sky130_fd_sc_hd__dfrtp_2
X_13820_ net58 _05683_ _06031_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_199_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25806_ top0.matmul0.alpha_pass\[1\] top0.matmul0.beta_pass\[1\] VGND VGND VPWR VPWR
+ _05033_ sky130_fd_sc_hd__or2_1
X_26786_ clknet_leaf_1_clk_sys _00403_ net582 VGND VGND VPWR VPWR top0.cordic0.sin\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23998_ _02976_ _02977_ _03057_ _03058_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__o22a_1
XFILLER_0_187_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13751_ net62 _05517_ _05961_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__and3_1
X_25737_ net73 _04954_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__nand2_1
X_22949_ _02458_ _02461_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16470_ _08554_ _08557_ VGND VGND VPWR VPWR _08558_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_168_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13682_ net47 _05682_ _05894_ net50 VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__a22o_1
X_25668_ net791 _04904_ _04936_ _04940_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15421_ _07332_ _07519_ VGND VGND VPWR VPWR _07520_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_167_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24619_ _03027_ _03028_ _03155_ _03156_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__o211ai_2
X_25599_ net73 _04886_ _04890_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__a21o_2
XFILLER_0_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18140_ _10121_ _10123_ VGND VGND VPWR VPWR _10124_ sky130_fd_sc_hd__xnor2_1
X_15352_ _07233_ _07404_ _07446_ _07447_ VGND VGND VPWR VPWR _07451_ sky130_fd_sc_hd__or4_1
XFILLER_0_110_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14303_ _06440_ _06511_ _06512_ VGND VGND VPWR VPWR _06513_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_124_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18071_ _09960_ _09969_ _10055_ VGND VGND VPWR VPWR _10056_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15283_ net525 _07374_ net479 VGND VGND VPWR VPWR _07382_ sky130_fd_sc_hd__o21ai_1
X_27269_ clknet_3_6__leaf_clk_mosi _00883_ VGND VGND VPWR VPWR spi0.data_packed\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17022_ top0.pid_q.prev_error\[14\] top0.pid_q.curr_error\[14\] VGND VGND VPWR VPWR
+ _09075_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14234_ _06442_ _06443_ _06440_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14165_ _06260_ _06267_ _06270_ _06271_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_42_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14096_ _05504_ _05543_ _05545_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__or3_1
X_18973_ net360 net316 VGND VGND VPWR VPWR _10947_ sky130_fd_sc_hd__or2_1
X_17924_ net1022 net404 VGND VGND VPWR VPWR _09910_ sky130_fd_sc_hd__nand2_2
XFILLER_0_79_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17855_ _09782_ _09786_ _09780_ VGND VGND VPWR VPWR _09842_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_191_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16806_ net506 _08855_ _08858_ net710 _08876_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__a221o_1
X_17786_ _09518_ _09771_ _09772_ VGND VGND VPWR VPWR _09773_ sky130_fd_sc_hd__and3_1
X_14998_ spi0.data_packed\[5\] top0.periodTop\[5\] _07108_ VGND VGND VPWR VPWR _07124_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19525_ net108 net103 net98 net94 net199 net193 VGND VGND VPWR VPWR _11415_ sky130_fd_sc_hd__mux4_2
X_16737_ _08287_ _07781_ net444 VGND VGND VPWR VPWR _08821_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13949_ _06123_ _06128_ _06138_ _06161_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19456_ _11351_ _11345_ _11352_ VGND VGND VPWR VPWR _11353_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16668_ _08751_ _08752_ net497 VGND VGND VPWR VPWR _08753_ sky130_fd_sc_hd__o21a_1
XFILLER_0_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18407_ net364 _10387_ VGND VGND VPWR VPWR _10388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_201_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15619_ _07636_ _07658_ _07637_ VGND VGND VPWR VPWR _07717_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_9_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19387_ _11292_ VGND VGND VPWR VPWR _11293_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16599_ _07701_ _08685_ VGND VGND VPWR VPWR _08686_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18338_ _10225_ _10230_ _10141_ VGND VGND VPWR VPWR _10320_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_45_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18269_ _10167_ _10241_ VGND VGND VPWR VPWR _10251_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20300_ _12146_ _12147_ _12137_ VGND VGND VPWR VPWR _12149_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21280_ _12699_ _13122_ net257 VGND VGND VPWR VPWR _13123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout5 _11517_ VGND VGND VPWR VPWR net1016 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20231_ net253 _12042_ VGND VGND VPWR VPWR _12080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_188_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20162_ _12013_ VGND VGND VPWR VPWR _12014_ sky130_fd_sc_hd__buf_2
XFILLER_0_200_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24970_ _04235_ _04318_ _04320_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20093_ _11857_ _11952_ VGND VGND VPWR VPWR _11953_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23921_ _03238_ _03277_ _03278_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26640_ clknet_leaf_80_clk_sys _00257_ net633 VGND VGND VPWR VPWR top0.pid_d.out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23852_ _02998_ _03000_ _03054_ _03055_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22803_ top0.svm0.tA\[5\] VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26571_ clknet_leaf_54_clk_sys _00194_ net667 VGND VGND VPWR VPWR top0.pid_q.curr_error\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_23783_ _03035_ _03138_ _03140_ _03085_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__a211o_1
XFILLER_0_200_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20995_ _12837_ _12841_ _11653_ _12778_ VGND VGND VPWR VPWR _12842_ sky130_fd_sc_hd__a211oi_1
X_25522_ _04847_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__clkbuf_1
X_22734_ net915 _11431_ net178 VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25453_ _04780_ _04795_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__xnor2_1
X_22665_ net99 net90 VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24404_ _02985_ _02987_ _03018_ _03019_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21616_ net146 VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__inv_2
X_25384_ _04670_ _04671_ _04727_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22596_ net103 _01980_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27123_ clknet_leaf_30_clk_sys _00737_ net623 VGND VGND VPWR VPWR top0.c_out_calc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_24335_ _03688_ _03691_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_145_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21547_ _01104_ _01108_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27054_ clknet_leaf_17_clk_sys _00671_ net609 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.d\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_24266_ net8 _03447_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__nand2_2
XFILLER_0_121_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21478_ top0.cordic0.cos\[11\] _12004_ _12036_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__and3_1
X_26005_ net430 _05203_ _05204_ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__a21o_1
X_23217_ net179 net215 VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__nand2_1
X_20429_ net291 _12277_ VGND VGND VPWR VPWR _12278_ sky130_fd_sc_hd__xnor2_4
X_24197_ _03547_ _03554_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23148_ _02635_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23079_ _02339_ _02538_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__xnor2_1
X_15970_ _07969_ _07973_ _07967_ VGND VGND VPWR VPWR _08065_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14921_ _07081_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__clkbuf_1
X_26907_ clknet_leaf_5_clk_sys _00524_ net590 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold50 top0.matmul0.matmul_stage_inst.d\[2\] VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 top0.cordic0.cos\[12\] VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 top0.pid_q.curr_int\[15\] VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__dlygate4sd3_1
X_17640_ _09468_ _09625_ _09626_ VGND VGND VPWR VPWR _09627_ sky130_fd_sc_hd__o21a_1
Xhold83 top0.svm0.tA\[2\] VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__dlygate4sd3_1
X_26838_ clknet_leaf_36_clk_sys _00455_ net676 VGND VGND VPWR VPWR top0.svm0.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_14852_ _07045_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold94 top0.cordic0.cos\[10\] VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_202_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13803_ _06003_ _06009_ _06014_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__a21o_1
X_14783_ _06960_ _06963_ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__and2_1
X_17571_ _09555_ _09554_ VGND VGND VPWR VPWR _09558_ sky130_fd_sc_hd__or2_1
XFILLER_0_187_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26769_ clknet_leaf_5_clk_sys _00386_ net590 VGND VGND VPWR VPWR top0.cordic0.cos\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_202_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19310_ _11249_ _11250_ VGND VGND VPWR VPWR _11251_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13734_ _05928_ _05943_ _05946_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16522_ _07701_ _08609_ VGND VGND VPWR VPWR _08610_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19241_ _11185_ _11186_ VGND VGND VPWR VPWR _11188_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13665_ _05830_ _05877_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__xnor2_4
X_16453_ _08492_ _08541_ VGND VGND VPWR VPWR _08542_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_151_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15404_ _07456_ _07457_ VGND VGND VPWR VPWR _07503_ sky130_fd_sc_hd__or2b_1
X_16384_ _08467_ _08473_ VGND VGND VPWR VPWR _08474_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19172_ _11123_ VGND VGND VPWR VPWR _11125_ sky130_fd_sc_hd__clkbuf_4
X_13596_ _05621_ _05804_ _05807_ _05808_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__a2bb2oi_4
XFILLER_0_5_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18123_ net1023 net403 VGND VGND VPWR VPWR _10107_ sky130_fd_sc_hd__nand2_1
X_15335_ _07414_ _07433_ VGND VGND VPWR VPWR _07434_ sky130_fd_sc_hd__and2_1
XFILLER_0_182_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18054_ _10007_ _10038_ VGND VGND VPWR VPWR _10039_ sky130_fd_sc_hd__xnor2_2
X_15266_ _07354_ _07364_ VGND VGND VPWR VPWR _07365_ sky130_fd_sc_hd__nand2b_2
XANTENNA_3 _02352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14217_ _06330_ _06426_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__nor2_2
X_17005_ _08899_ _09056_ _09058_ VGND VGND VPWR VPWR _09059_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15197_ _07194_ _07294_ _07295_ VGND VGND VPWR VPWR _07296_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_46_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14148_ _06124_ _06125_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14079_ _05565_ _05637_ _05638_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__or3_1
X_18956_ _10847_ _10928_ _10929_ VGND VGND VPWR VPWR _10930_ sky130_fd_sc_hd__o21ai_2
X_17907_ net439 _09339_ _09892_ _09893_ VGND VGND VPWR VPWR _09894_ sky130_fd_sc_hd__and4_1
X_18887_ _09395_ _10778_ _09356_ VGND VGND VPWR VPWR _10862_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_175_Right_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17838_ _09812_ _09815_ VGND VGND VPWR VPWR _09825_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17769_ _09754_ _09755_ VGND VGND VPWR VPWR _09756_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19508_ top0.pid_d.curr_int\[14\] top0.pid_d.prev_int\[14\] VGND VGND VPWR VPWR _11399_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20780_ net299 _12156_ _12611_ VGND VGND VPWR VPWR _12629_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_190_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19439_ _11336_ _11337_ VGND VGND VPWR VPWR _11338_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_174_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22450_ _01986_ _02005_ _02006_ _01985_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__a31o_2
XFILLER_0_18_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21401_ _00944_ _00945_ _00967_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22381_ _01936_ _01939_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_199_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24120_ _03456_ _03471_ _03477_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_26_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21332_ _11727_ net231 VGND VGND VPWR VPWR _13174_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24051_ _03400_ _03407_ _03408_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_41_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21263_ _13015_ _13106_ VGND VGND VPWR VPWR _13107_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_124_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23002_ _02345_ _02297_ _02505_ _02507_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__a31o_1
XFILLER_0_163_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20214_ _11550_ _12061_ VGND VGND VPWR VPWR _12063_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21194_ _13036_ _13037_ VGND VGND VPWR VPWR _13038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_198_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20145_ net180 _11974_ net212 VGND VGND VPWR VPWR _12000_ sky130_fd_sc_hd__or3b_1
X_24953_ _04212_ _04233_ _04214_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__o21ba_1
X_20076_ _11428_ _11936_ VGND VGND VPWR VPWR _11937_ sky130_fd_sc_hd__nand2_1
X_23904_ _03257_ _03258_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__xor2_2
XFILLER_0_100_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24884_ _04179_ _04235_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26623_ clknet_leaf_29_clk_sys _00240_ net623 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_23835_ _03175_ _03176_ _03192_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__a21o_1
XFILLER_0_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26554_ clknet_leaf_52_clk_sys _00177_ net670 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_23766_ _03093_ _03094_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__or2_2
XFILLER_0_135_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20978_ net227 _12822_ _12823_ _12824_ VGND VGND VPWR VPWR _12825_ sky130_fd_sc_hd__a22o_1
X_25505_ _04838_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__clkbuf_1
X_22717_ _01877_ _02267_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__or2_1
X_26485_ clknet_leaf_89_clk_sys _00116_ net603 VGND VGND VPWR VPWR top0.periodTop\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_23697_ net566 net560 top0.matmul0.matmul_stage_inst.e\[7\] VGND VGND VPWR VPWR _03055_
+ sky130_fd_sc_hd__o21a_4
XFILLER_0_32_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25436_ _04777_ _04778_ _04728_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__mux2_1
X_13450_ _05662_ _05601_ _05470_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__or3b_1
XFILLER_0_94_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22648_ _02199_ _02200_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__xor2_1
XFILLER_0_152_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25367_ _04711_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__clkbuf_1
X_13381_ _05582_ _05593_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__xnor2_2
X_22579_ net769 _12813_ _02133_ _12963_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15120_ _07196_ _07217_ _07218_ VGND VGND VPWR VPWR _07219_ sky130_fd_sc_hd__and3_1
X_24318_ _03673_ _03674_ _03666_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__mux2_1
X_27106_ clknet_leaf_21_clk_sys _00723_ net610 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.a\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_25298_ _04639_ _04643_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_181_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_27037_ clknet_leaf_8_clk_sys _00654_ net592 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_15051_ net531 net471 VGND VGND VPWR VPWR _07150_ sky130_fd_sc_hd__nand2_1
X_24249_ _03548_ _03547_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__and2b_1
X_14002_ net32 _06213_ _06214_ net1030 VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__o22a_1
Xoutput5 net5 VGND VGND VPWR VPWR pwmB sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18810_ _10769_ _10785_ VGND VGND VPWR VPWR _10786_ sky130_fd_sc_hd__xnor2_4
X_19790_ _11653_ _11670_ _11671_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__a21oi_1
X_18741_ _10635_ _10640_ _10717_ VGND VGND VPWR VPWR _10718_ sky130_fd_sc_hd__a21o_1
X_15953_ net488 _07914_ VGND VGND VPWR VPWR _08048_ sky130_fd_sc_hd__xor2_4
X_14904_ _07072_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__clkbuf_1
X_18672_ _10550_ _10553_ _10549_ VGND VGND VPWR VPWR _10650_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_105_clk_sys clknet_3_0__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_105_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_64_clk_sys clknet_3_5__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_64_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_15884_ _07869_ VGND VGND VPWR VPWR _07980_ sky130_fd_sc_hd__inv_2
X_17623_ net1023 net427 VGND VGND VPWR VPWR _09610_ sky130_fd_sc_hd__and2_1
X_14835_ _07032_ _07033_ VGND VGND VPWR VPWR _07034_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17554_ _09521_ _09527_ VGND VGND VPWR VPWR _09541_ sky130_fd_sc_hd__xnor2_2
X_14766_ _06951_ _06967_ VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16505_ _08532_ _08537_ _08538_ VGND VGND VPWR VPWR _08593_ sky130_fd_sc_hd__o21a_1
XFILLER_0_156_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13717_ _05910_ _05911_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__xor2_1
X_14697_ _06899_ _06900_ VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__and2_1
X_17485_ _09468_ _09471_ VGND VGND VPWR VPWR _09472_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_184_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19224_ net339 _11117_ _11170_ _11172_ _08889_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__o221a_1
XFILLER_0_160_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16436_ _08436_ _08438_ _08524_ VGND VGND VPWR VPWR _08525_ sky130_fd_sc_hd__o21a_1
X_13648_ top0.periodTop_r\[1\] _05640_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19155_ top0.kid\[12\] _11097_ _11099_ top0.kpd\[12\] VGND VGND VPWR VPWR _11113_
+ sky130_fd_sc_hd__a22o_1
X_13579_ _05653_ _05655_ _05791_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__a21o_1
X_16367_ _08444_ _08455_ VGND VGND VPWR VPWR _08457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18106_ _10031_ _10033_ _10089_ VGND VGND VPWR VPWR _10090_ sky130_fd_sc_hd__o21ai_1
X_15318_ _07355_ _07416_ VGND VGND VPWR VPWR _07417_ sky130_fd_sc_hd__xnor2_1
X_16298_ _08307_ _08388_ VGND VGND VPWR VPWR _08389_ sky130_fd_sc_hd__xnor2_1
X_19086_ net311 _10384_ net308 _09965_ VGND VGND VPWR VPWR _11058_ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18037_ _10013_ _10021_ VGND VGND VPWR VPWR _10022_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15249_ _07344_ _07345_ _07346_ _07347_ VGND VGND VPWR VPWR _07348_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_22_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout307 top0.pid_d.mult0.b\[15\] VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout318 net319 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__buf_1
X_19988_ net10 _11855_ VGND VGND VPWR VPWR _11856_ sky130_fd_sc_hd__xnor2_1
Xfanout329 top0.pid_d.mult0.b\[8\] VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__buf_4
X_18939_ top0.pid_d.out\[11\] top0.pid_d.curr_int\[11\] VGND VGND VPWR VPWR _10914_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21950_ net161 net137 VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_19_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_179_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20901_ _12238_ _12747_ _12748_ VGND VGND VPWR VPWR _12749_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21881_ _01281_ _01442_ _01437_ net156 VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_178_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23620_ _02976_ _02977_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__nor2_2
X_20832_ _12209_ _12680_ _12204_ VGND VGND VPWR VPWR _12681_ sky130_fd_sc_hd__o21ai_2
X_23551_ top0.a_in_matmul\[15\] top0.matmul0.a\[15\] _02937_ VGND VGND VPWR VPWR _02942_
+ sky130_fd_sc_hd__mux2_1
X_20763_ net300 _11550_ VGND VGND VPWR VPWR _12612_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22502_ _02057_ _01224_ _01312_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26270_ net958 net944 net688 VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23482_ net928 top0.matmul0.sin\[10\] _02904_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__mux2_1
X_20694_ _12359_ _12384_ _12536_ _12542_ VGND VGND VPWR VPWR _12543_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25221_ _04553_ _04567_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__xor2_2
X_22433_ _01885_ _01941_ _01898_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_190_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_28_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_190_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_25152_ _04437_ _04439_ _04499_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22364_ _01779_ _01922_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24103_ _03457_ _03460_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__xnor2_2
X_21315_ _13138_ _13136_ _13156_ VGND VGND VPWR VPWR _13157_ sky130_fd_sc_hd__o21a_1
X_25083_ _04428_ _04431_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22295_ _01845_ _01854_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24034_ _03388_ _03389_ _03391_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__o21ai_2
X_21246_ _13058_ _13089_ _12546_ VGND VGND VPWR VPWR _13090_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_130_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21177_ _12983_ _13020_ _12985_ VGND VGND VPWR VPWR _13021_ sky130_fd_sc_hd__o21ba_1
X_20128_ _11978_ VGND VGND VPWR VPWR _11984_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25985_ top0.matmul0.beta_pass\[6\] _05169_ _05188_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_37_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24936_ _04187_ _04193_ _04286_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__o21a_1
X_20059_ _11526_ _11921_ net178 VGND VGND VPWR VPWR _11922_ sky130_fd_sc_hd__o21a_1
X_24867_ _02994_ _02996_ _03162_ _03163_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__o22a_1
X_14620_ net41 _06824_ _06768_ _06769_ VGND VGND VPWR VPWR _06825_ sky130_fd_sc_hd__a22o_1
X_26606_ clknet_leaf_86_clk_sys _00017_ net641 VGND VGND VPWR VPWR top0.pid_d.state\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_197_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23818_ _03174_ _03170_ _03171_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__nand3_1
X_24798_ _04146_ _04148_ _04150_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14551_ _06755_ _06756_ VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_184_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23749_ _03093_ _03094_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__nor2_1
X_26537_ clknet_leaf_60_clk_sys _00160_ net652 VGND VGND VPWR VPWR top0.pid_q.mult0.a\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13502_ _05649_ _05651_ _05714_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__a21bo_1
X_14482_ _06557_ _06686_ _06688_ _06610_ VGND VGND VPWR VPWR _06689_ sky130_fd_sc_hd__o2bb2a_1
X_17270_ top0.matmul0.matmul_stage_inst.mult2\[3\] _09265_ top0.matmul0.matmul_stage_inst.mult1\[3\]
+ VGND VGND VPWR VPWR _09269_ sky130_fd_sc_hd__a21o_1
X_26468_ clknet_leaf_16_clk_sys net570 net611 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13433_ _05643_ _05645_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__xnor2_1
X_16221_ _08312_ _08222_ VGND VGND VPWR VPWR _08313_ sky130_fd_sc_hd__and2_1
X_25419_ _04762_ _04664_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26399_ clknet_leaf_98_clk_sys _00040_ net588 VGND VGND VPWR VPWR top0.kpd\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16152_ _08243_ _08239_ top0.pid_q.out\[6\] VGND VGND VPWR VPWR _08244_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13364_ _05564_ _05570_ _05576_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15103_ _07156_ _07157_ _07155_ VGND VGND VPWR VPWR _07202_ sky130_fd_sc_hd__o21ai_1
X_16083_ _08115_ _08117_ _08175_ VGND VGND VPWR VPWR _08176_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13295_ _05499_ _05507_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__xnor2_1
X_15034_ net964 _07140_ _07144_ top0.pid_d.curr_int\[4\] VGND VGND VPWR VPWR _00121_
+ sky130_fd_sc_hd__a22o_1
X_19911_ _11784_ VGND VGND VPWR VPWR _11785_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19842_ _11514_ _11719_ VGND VGND VPWR VPWR _11720_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19773_ _11415_ _11416_ _11654_ VGND VGND VPWR VPWR _11655_ sky130_fd_sc_hd__mux2_1
X_16985_ top0.matmul0.beta_pass\[11\] _09038_ _09039_ VGND VGND VPWR VPWR _09040_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_78_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18724_ _10458_ _10644_ net341 VGND VGND VPWR VPWR _10701_ sky130_fd_sc_hd__o21a_1
X_15936_ _08027_ _08030_ VGND VGND VPWR VPWR _08031_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18655_ net362 _10632_ VGND VGND VPWR VPWR _10633_ sky130_fd_sc_hd__nand2_4
X_15867_ _07930_ _07962_ VGND VGND VPWR VPWR _07963_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17606_ net423 VGND VGND VPWR VPWR _09593_ sky130_fd_sc_hd__inv_2
X_14818_ _07014_ _07015_ _07017_ VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__a21oi_1
X_18586_ net309 _10452_ _10563_ _09353_ VGND VGND VPWR VPWR _10565_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15798_ _07810_ _07894_ VGND VGND VPWR VPWR _07895_ sky130_fd_sc_hd__xor2_2
XFILLER_0_176_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17537_ net423 net343 net425 VGND VGND VPWR VPWR _09524_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14749_ _06896_ _06916_ _06950_ VGND VGND VPWR VPWR _06951_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_19_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17468_ _09439_ _09453_ _09454_ _09437_ VGND VGND VPWR VPWR _09455_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19207_ top0.pid_d.prev_error\[4\] top0.pid_d.curr_error\[4\] VGND VGND VPWR VPWR
+ _11157_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_172_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16419_ _08420_ _08425_ _08415_ VGND VGND VPWR VPWR _08508_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_61_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17399_ _09376_ _09385_ VGND VGND VPWR VPWR _09386_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19138_ net415 _11096_ _11104_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19069_ _11016_ _11040_ _11014_ VGND VGND VPWR VPWR _11041_ sky130_fd_sc_hd__or3b_1
XFILLER_0_140_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_196_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21100_ _12749_ _12802_ VGND VGND VPWR VPWR _12946_ sky130_fd_sc_hd__and2b_1
X_22080_ net115 net102 net97 _01641_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21031_ _12875_ _12877_ VGND VGND VPWR VPWR _12878_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout104 net105 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_196_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout115 net116 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_4
Xfanout126 net128 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout137 top0.cordic0.vec\[1\]\[5\] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_2
Xfanout148 net149 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_4
Xfanout159 top0.cordic0.vec\[1\]\[1\] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_201_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22982_ top0.svm0.counter\[8\] _02489_ _02490_ _02488_ VGND VGND VPWR VPWR _00450_
+ sky130_fd_sc_hd__a22o_1
X_25770_ _04886_ top0.matmul0.cos\[13\] _04878_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24721_ _02985_ _02987_ _03162_ _03163_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__o22a_1
X_21933_ net163 _01123_ _01280_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_179_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24652_ _04003_ _04004_ _04001_ _04002_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_139_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21864_ _01391_ _01425_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_194_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23603_ _02968_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20815_ _12475_ _12486_ VGND VGND VPWR VPWR _12664_ sky130_fd_sc_hd__xnor2_1
X_24583_ _03824_ _03935_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__nand2_1
X_21795_ net158 _01356_ _01179_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__mux2_1
X_26322_ spi0.data_packed\[59\] spi0.data_packed\[60\] net699 VGND VGND VPWR VPWR
+ _05393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23534_ top0.a_in_matmul\[7\] top0.matmul0.a\[7\] _02926_ VGND VGND VPWR VPWR _02933_
+ sky130_fd_sc_hd__mux2_1
X_20746_ _12264_ _12551_ VGND VGND VPWR VPWR _12595_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26253_ _05358_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__clkbuf_1
X_23465_ top0.cordic0.sin\[2\] top0.matmul0.sin\[2\] _05461_ VGND VGND VPWR VPWR _02897_
+ sky130_fd_sc_hd__mux2_1
X_20677_ net263 _12490_ VGND VGND VPWR VPWR _12526_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_4_clk_sys clknet_3_0__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_4_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_169_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_12_clk_sys clknet_3_3__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_12_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25204_ _04547_ _04550_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_150_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22416_ net97 _01230_ _01779_ _01922_ _11674_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__a221o_1
XFILLER_0_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26184_ _05319_ top0.cordic0.slte0.opB\[12\] _12003_ VGND VGND VPWR VPWR _05320_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23396_ _02824_ _02825_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_25135_ _04422_ _04481_ _04482_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22347_ net79 net87 _01902_ _01905_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25066_ _03234_ _03502_ _04131_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22278_ net144 net126 _01836_ _01837_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__a31o_1
XFILLER_0_130_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24017_ _03359_ _03362_ _03371_ VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__nand3_1
X_21229_ _12622_ _13072_ VGND VGND VPWR VPWR _13073_ sky130_fd_sc_hd__nand2_1
Xhold180 top0.pid_d.prev_error\[7\] VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 top0.matmul0.matmul_stage_inst.b\[11\] VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout660 net661 VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__clkbuf_4
Xfanout671 net673 VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__clkbuf_4
Xfanout682 net685 VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__clkbuf_4
X_16770_ top0.pid_q.state\[0\] net544 VGND VGND VPWR VPWR _08853_ sky130_fd_sc_hd__or2_2
XFILLER_0_176_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13982_ _06193_ _06194_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__xor2_1
Xfanout693 net700 VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__buf_2
X_25968_ top0.pid_q.out\[2\] _12032_ _05014_ spi0.data_packed\[50\] VGND VGND VPWR
+ VPWR _05176_ sky130_fd_sc_hd__a22o_1
X_15721_ _07719_ _07720_ _07721_ VGND VGND VPWR VPWR _07818_ sky130_fd_sc_hd__o21ai_1
X_24919_ _04198_ _04210_ _04269_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_38_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25899_ _05437_ _05104_ _05102_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_77_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18440_ _10323_ _10419_ _10418_ VGND VGND VPWR VPWR _10421_ sky130_fd_sc_hd__a21o_1
X_15652_ _07649_ _07654_ VGND VGND VPWR VPWR _07750_ sky130_fd_sc_hd__nor2_1
X_14603_ _06685_ _06744_ VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18371_ net319 _10350_ _10351_ _10208_ VGND VGND VPWR VPWR _10352_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15583_ _07546_ _07547_ VGND VGND VPWR VPWR _07682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17322_ _09312_ _09313_ VGND VGND VPWR VPWR _09314_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14534_ _06656_ _06657_ _06654_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17253_ _09253_ _09254_ VGND VGND VPWR VPWR _09255_ sky130_fd_sc_hd__xnor2_1
X_14465_ _06553_ _06556_ VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__nor2_2
XFILLER_0_37_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16204_ _08286_ _08295_ VGND VGND VPWR VPWR _08296_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13416_ _05608_ _05609_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__or2_2
XFILLER_0_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14396_ _06535_ _06530_ _06604_ VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__nor3_1
XFILLER_0_52_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17184_ _09193_ _09187_ _09194_ VGND VGND VPWR VPWR _09195_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13347_ net52 _05517_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__nand2_1
X_16135_ _08143_ _08145_ VGND VGND VPWR VPWR _08228_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_183_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13278_ _05490_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__buf_2
X_16066_ _07800_ _08159_ VGND VGND VPWR VPWR _08160_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15017_ spi0.data_packed\[14\] top0.periodTop\[14\] _07125_ VGND VGND VPWR VPWR _07134_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19825_ _11514_ _11702_ _11700_ VGND VGND VPWR VPWR _11704_ sky130_fd_sc_hd__and3_1
XFILLER_0_166_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_194_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19756_ _11612_ net187 _11634_ _11638_ VGND VGND VPWR VPWR _11639_ sky130_fd_sc_hd__o31a_1
X_16968_ _08882_ _09016_ _09023_ _09024_ _07800_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__o311a_1
X_18707_ _10606_ _10677_ _10683_ VGND VGND VPWR VPWR _10684_ sky130_fd_sc_hd__o21ai_2
X_15919_ net451 net526 VGND VGND VPWR VPWR _08014_ sky130_fd_sc_hd__nand2_1
X_19687_ _11572_ VGND VGND VPWR VPWR _11573_ sky130_fd_sc_hd__clkbuf_4
X_16899_ top0.matmul0.done_pass top0.matmul0.state\[1\] top0.matmul0.beta_pass\[6\]
+ VGND VGND VPWR VPWR _08960_ sky130_fd_sc_hd__and3_1
XFILLER_0_155_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18638_ net381 net314 VGND VGND VPWR VPWR _10616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_176_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18569_ _10543_ _10547_ VGND VGND VPWR VPWR _10548_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_192_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20600_ net287 _12059_ net302 VGND VGND VPWR VPWR _12449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21580_ _01134_ _01141_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__xor2_2
XFILLER_0_129_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20531_ _12316_ _12320_ _12319_ VGND VGND VPWR VPWR _12380_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23250_ _02699_ VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20462_ _11527_ _12308_ _12309_ _12310_ VGND VGND VPWR VPWR _12311_ sky130_fd_sc_hd__a31o_1
XFILLER_0_144_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22201_ net100 net95 VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_23181_ _02648_ VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20393_ _12230_ _12241_ VGND VGND VPWR VPWR _12242_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22132_ _01686_ _01689_ _01690_ _01693_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__o31a_1
XFILLER_0_101_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22063_ _01557_ _01558_ _01621_ _01552_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__a211o_1
X_26940_ clknet_leaf_9_clk_sys _00557_ net594 VGND VGND VPWR VPWR top0.matmul0.a\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_21014_ _12843_ _12860_ VGND VGND VPWR VPWR _12861_ sky130_fd_sc_hd__xnor2_2
X_26871_ clknet_leaf_37_clk_sys _00488_ net678 VGND VGND VPWR VPWR top0.svm0.tA\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25822_ top0.matmul0.alpha_pass\[3\] top0.matmul0.beta_pass\[3\] VGND VGND VPWR VPWR
+ _05047_ sky130_fd_sc_hd__xor2_2
X_22965_ _06277_ _02475_ net172 VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__o21a_1
X_25753_ net717 _04925_ _04997_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__a21o_1
X_24704_ _04049_ _04057_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__xnor2_1
X_21916_ _01472_ _01476_ _01477_ _01320_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__o22a_1
X_22896_ _02332_ top0.svm0.tC\[4\] _02412_ top0.svm0.tC\[3\] _02413_ VGND VGND VPWR
+ VPWR _02414_ sky130_fd_sc_hd__o221a_1
X_25684_ top0.matmul0.sin\[12\] _04952_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24635_ _03983_ _03988_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__xnor2_1
X_21847_ net135 net121 VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_194_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24566_ _03915_ _03919_ _03920_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__or3_2
XFILLER_0_194_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_21778_ net135 _01299_ _01336_ _01339_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_93_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26305_ _05384_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__clkbuf_1
X_20729_ _12577_ VGND VGND VPWR VPWR _12578_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23517_ top0.cordic0.cos\[13\] top0.matmul0.cos\[13\] _02915_ VGND VGND VPWR VPWR
+ _02924_ sky130_fd_sc_hd__mux2_1
X_24497_ _03851_ _03852_ _03658_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27285_ clknet_3_2__leaf_clk_mosi _00899_ VGND VGND VPWR VPWR spi0.data_packed\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14250_ _06303_ _06341_ _06342_ VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_108_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23448_ net88 _11783_ _02882_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__or3_1
X_26236_ spi0.data_packed\[16\] spi0.data_packed\[17\] net697 VGND VGND VPWR VPWR
+ _05350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13201_ top0.pid_q.state\[0\] _05427_ net16 net544 VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__a211o_1
X_14181_ _06344_ _06391_ _06346_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__o21a_1
X_23379_ net116 _11857_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__nor2_1
X_26167_ _05306_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25118_ _04466_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26098_ _05275_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__buf_2
XFILLER_0_143_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25049_ _04391_ _04398_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__xor2_2
X_17940_ _09834_ _09835_ _09836_ VGND VGND VPWR VPWR _09926_ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_178_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17871_ _09840_ _09857_ VGND VGND VPWR VPWR _09858_ sky130_fd_sc_hd__xnor2_2
X_19610_ top0.cordic0.slte0.opB\[10\] VGND VGND VPWR VPWR _11499_ sky130_fd_sc_hd__inv_2
X_16822_ net1019 VGND VGND VPWR VPWR _08889_ sky130_fd_sc_hd__buf_4
XFILLER_0_40_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout490 net492 VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__dlymetal6s2s_1
X_19541_ _11430_ VGND VGND VPWR VPWR _11431_ sky130_fd_sc_hd__buf_4
X_16753_ _08831_ _08836_ VGND VGND VPWR VPWR _08837_ sky130_fd_sc_hd__xnor2_1
X_13965_ _05858_ _06082_ _06177_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__a21o_2
X_15704_ top0.pid_q.out\[2\] _07703_ VGND VGND VPWR VPWR _07801_ sky130_fd_sc_hd__nor2_1
X_19472_ _11366_ _11359_ _10834_ VGND VGND VPWR VPWR _11367_ sky130_fd_sc_hd__a21o_1
X_16684_ _08762_ _08768_ VGND VGND VPWR VPWR _08769_ sky130_fd_sc_hd__xnor2_2
X_13896_ _06104_ _06108_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__xnor2_4
X_18423_ net307 _10403_ VGND VGND VPWR VPWR _10404_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15635_ _07642_ _07646_ _07644_ VGND VGND VPWR VPWR _07733_ sky130_fd_sc_hd__o21a_1
XFILLER_0_152_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18354_ net1018 _10335_ VGND VGND VPWR VPWR _10336_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15566_ _07557_ _07558_ _07664_ VGND VGND VPWR VPWR _07665_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_173_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17305_ _09298_ _09294_ top0.matmul0.matmul_stage_inst.mult1\[8\] VGND VGND VPWR
+ VPWR _09299_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_51_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14517_ _06622_ _06627_ _06619_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_185_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18285_ _10192_ _10194_ _10190_ VGND VGND VPWR VPWR _10267_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_56_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15497_ _07594_ _07595_ VGND VGND VPWR VPWR _07596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17236_ top0.pid_q.curr_int\[14\] _09237_ _09240_ VGND VGND VPWR VPWR _09241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14448_ _06562_ _06563_ _06655_ VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__o21a_1
XFILLER_0_181_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17167_ _09178_ _09179_ VGND VGND VPWR VPWR _09180_ sky130_fd_sc_hd__nand2_1
X_14379_ _06517_ _06519_ _06518_ VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16118_ _08205_ _08210_ VGND VGND VPWR VPWR _08211_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17098_ net818 _09115_ _09125_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__a21o_1
XFILLER_0_177_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16049_ net483 _08141_ _08003_ _08142_ VGND VGND VPWR VPWR _08143_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19808_ net175 _11673_ _11687_ _11688_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__a31o_1
X_19739_ net286 _11619_ VGND VGND VPWR VPWR _11623_ sky130_fd_sc_hd__nand2_1
XFILLER_0_193_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22750_ _11785_ _12034_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__nand2_1
X_21701_ net122 net106 VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__xnor2_2
X_22681_ _02180_ _02184_ _02209_ _02230_ _02232_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__o32a_1
XFILLER_0_47_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24420_ _03686_ _03692_ _03684_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21632_ _01184_ _01190_ _01193_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_47_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_24351_ _03705_ _03706_ _03703_ _03704_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21563_ net127 net124 VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__nor2_1
X_23302_ net138 _11784_ _02747_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__or3_1
X_27070_ clknet_leaf_2_clk_sys _00687_ net584 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.c\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_20514_ _12280_ _12360_ VGND VGND VPWR VPWR _12363_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24282_ _03634_ _03636_ _03637_ _03639_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__and4_2
XFILLER_0_117_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21494_ _01014_ _00994_ _01040_ _12744_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__a31o_1
XFILLER_0_117_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26021_ net428 _05203_ _05216_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__a21o_1
X_23233_ _01320_ _01267_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__nor2_1
X_20445_ _12250_ _12293_ VGND VGND VPWR VPWR _12294_ sky130_fd_sc_hd__or2b_1
XFILLER_0_127_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23164_ _02641_ _06473_ _02645_ net783 VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__a22o_1
X_20376_ net276 _12127_ _12131_ VGND VGND VPWR VPWR _12225_ sky130_fd_sc_hd__nor3_1
XFILLER_0_28_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_189_Right_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22115_ _01637_ _01675_ _01612_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__a21oi_1
X_23095_ _02595_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__buf_2
X_22046_ _01606_ _01348_ _01353_ _01607_ _01362_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__a32o_1
X_26923_ clknet_leaf_4_clk_sys _00540_ net581 VGND VGND VPWR VPWR top0.matmul0.cos\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_26854_ clknet_leaf_46_clk_sys _00471_ net680 VGND VGND VPWR VPWR top0.svm0.delta\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_199_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25805_ net833 _05029_ _05031_ _05032_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__a22o_1
X_26785_ clknet_leaf_3_clk_sys _00402_ net582 VGND VGND VPWR VPWR top0.cordic0.sin\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_23997_ _03040_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_202_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13750_ _05960_ _05961_ _05962_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__o21a_1
X_25736_ net813 _04890_ _04913_ _04988_ VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__a22o_1
X_22948_ top0.svm0.delta\[3\] _02453_ _02460_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_58_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13681_ _05893_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__buf_2
XFILLER_0_97_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_25667_ top0.matmul0.sin\[8\] _04939_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__xor2_1
X_22879_ net169 _02381_ _02397_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_195_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15420_ _07330_ _07349_ VGND VGND VPWR VPWR _07519_ sky130_fd_sc_hd__xor2_1
X_24618_ _03155_ _03156_ _03027_ _03028_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25598_ _05456_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__buf_2
XFILLER_0_54_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15351_ _07415_ _07417_ VGND VGND VPWR VPWR _07450_ sky130_fd_sc_hd__xnor2_1
X_24549_ _03902_ _03903_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14302_ _06433_ _06434_ _06511_ _06440_ VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__o22a_1
XFILLER_0_109_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18070_ _09960_ _09969_ _09961_ VGND VGND VPWR VPWR _10055_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15282_ _07378_ _07379_ _07333_ VGND VGND VPWR VPWR _07381_ sky130_fd_sc_hd__a21o_1
X_27268_ clknet_3_6__leaf_clk_mosi _00882_ VGND VGND VPWR VPWR spi0.data_packed\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_202_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17021_ top0.pid_q.prev_error\[14\] top0.pid_q.curr_error\[14\] VGND VGND VPWR VPWR
+ _09074_ sky130_fd_sc_hd__and2_1
XFILLER_0_184_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14233_ _06440_ _06442_ _06443_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__nand3_2
XFILLER_0_124_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26219_ _05341_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__clkbuf_1
X_27199_ clknet_leaf_91_clk_sys _00813_ net599 VGND VGND VPWR VPWR top0.cordic0.slte0.opB\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14164_ _06255_ _06373_ _06375_ _06178_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__o22a_1
XFILLER_0_132_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14095_ _06094_ _05538_ _05539_ VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__or3_1
X_18972_ net360 _10384_ _10945_ VGND VGND VPWR VPWR _10946_ sky130_fd_sc_hd__a21o_1
X_17923_ _09827_ _09828_ _09908_ VGND VGND VPWR VPWR _09909_ sky130_fd_sc_hd__a21bo_1
X_17854_ _09782_ _09786_ VGND VGND VPWR VPWR _09841_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16805_ top0.kiq\[12\] _05448_ _08866_ VGND VGND VPWR VPWR _08876_ sky130_fd_sc_hd__and3_1
X_17785_ net378 _09636_ VGND VGND VPWR VPWR _09772_ sky130_fd_sc_hd__xor2_1
X_14997_ _07123_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19524_ net83 net88 _11413_ VGND VGND VPWR VPWR _11414_ sky130_fd_sc_hd__mux2_1
X_16736_ _08817_ _08819_ VGND VGND VPWR VPWR _08820_ sky130_fd_sc_hd__xnor2_1
X_13948_ _06155_ _06160_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__xor2_2
XFILLER_0_191_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19455_ _11351_ _11345_ _10594_ VGND VGND VPWR VPWR _11352_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16667_ _08654_ _08711_ VGND VGND VPWR VPWR _08752_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13879_ _06088_ _06089_ _06090_ _06091_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_201_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18406_ net341 net344 net348 VGND VGND VPWR VPWR _10387_ sky130_fd_sc_hd__or3_1
XFILLER_0_147_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15618_ _07714_ _07686_ _07715_ VGND VGND VPWR VPWR _07716_ sky130_fd_sc_hd__a21oi_1
X_19386_ _11289_ _11291_ VGND VGND VPWR VPWR _11292_ sky130_fd_sc_hd__nor2_2
X_16598_ _08682_ _08683_ _08684_ VGND VGND VPWR VPWR _08685_ sky130_fd_sc_hd__mux2_2
XFILLER_0_189_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18337_ _10222_ _10234_ _10233_ VGND VGND VPWR VPWR _10319_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15549_ _07642_ _07647_ VGND VGND VPWR VPWR _07648_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18268_ _10167_ _10241_ VGND VGND VPWR VPWR _10250_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17219_ top0.pid_q.curr_int\[12\] top0.pid_q.prev_int\[12\] VGND VGND VPWR VPWR _09226_
+ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_59_clk_sys clknet_3_4__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_59_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_18199_ _10180_ _10181_ VGND VGND VPWR VPWR _10182_ sky130_fd_sc_hd__or2b_1
XFILLER_0_141_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20230_ _12044_ _12046_ _12051_ VGND VGND VPWR VPWR _12079_ sky130_fd_sc_hd__a21bo_1
Xfanout6 _03020_ VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__buf_4
XFILLER_0_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20161_ top0.state\[1\] _12012_ VGND VGND VPWR VPWR _12013_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_196_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20092_ _11949_ _11951_ VGND VGND VPWR VPWR _11952_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23920_ _03239_ _03240_ VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23851_ _03207_ _03208_ _03061_ _03062_ VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22802_ top0.svm0.tA\[4\] VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__inv_2
X_26570_ clknet_leaf_52_clk_sys _00193_ net673 VGND VGND VPWR VPWR top0.pid_q.curr_error\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_23782_ _03042_ _03052_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__nor2_1
X_20994_ net267 _12135_ VGND VGND VPWR VPWR _12841_ sky130_fd_sc_hd__nand2_1
XFILLER_0_196_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25521_ top0.matmul0.b\[0\] top0.matmul0.matmul_stage_inst.f\[0\] _04846_ VGND VGND
+ VPWR VPWR _04847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_22733_ net740 _12813_ _02281_ _12742_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25452_ _04786_ _04794_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22664_ net101 net90 net86 VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24403_ _03502_ _03758_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21615_ net146 net154 VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_180_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25383_ _04670_ _04671_ _04669_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__a21bo_1
X_22595_ _01074_ _01769_ _02146_ net100 _02148_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_27122_ clknet_leaf_33_clk_sys _00736_ net665 VGND VGND VPWR VPWR top0.c_out_calc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_24334_ _03689_ _03690_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_118_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21546_ _01106_ _01107_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24265_ _03620_ _03622_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27053_ clknet_leaf_20_clk_sys _00670_ net609 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.d\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_21477_ _01040_ _01041_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_26004_ top0.pid_q.out\[10\] _05198_ _05199_ spi0.data_packed\[58\] VGND VGND VPWR
+ VPWR _05204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23216_ _02663_ _02664_ _02665_ _02666_ _11572_ _11576_ VGND VGND VPWR VPWR _02667_
+ sky130_fd_sc_hd__mux4_1
X_20428_ net300 net297 VGND VGND VPWR VPWR _12277_ sky130_fd_sc_hd__nor2b_2
X_24196_ _03548_ _03553_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23147_ _02633_ _02634_ top0.svm0.delta\[14\] VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__mux2_1
X_20359_ net234 _12207_ VGND VGND VPWR VPWR _12208_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_140_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23078_ _02577_ _02578_ _02298_ net65 VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__a211o_1
XFILLER_0_140_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_22029_ _01590_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__inv_2
X_14920_ spi0.data_packed\[35\] top0.kid\[3\] _07075_ VGND VGND VPWR VPWR _07081_
+ sky130_fd_sc_hd__mux2_1
X_26906_ clknet_leaf_5_clk_sys _00523_ net581 VGND VGND VPWR VPWR top0.cordic0.vec\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold40 top0.cordic0.sin\[13\] VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 top0.kpq\[4\] VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold62 top0.cordic0.cos\[5\] VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__dlygate4sd3_1
X_26837_ clknet_leaf_36_clk_sys _00454_ net676 VGND VGND VPWR VPWR top0.svm0.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold73 _00434_ VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ spi0.data_packed\[66\] top0.kpd\[2\] _07042_ VGND VGND VPWR VPWR _07045_
+ sky130_fd_sc_hd__mux2_1
Xhold84 top0.matmul0.matmul_stage_inst.b\[4\] VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 top0.svm0.tA\[1\] VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ _06003_ _06009_ _06014_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__nand3_1
XFILLER_0_187_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17570_ _09555_ _09556_ VGND VGND VPWR VPWR _09557_ sky130_fd_sc_hd__or2_1
X_14782_ _06960_ _06963_ VGND VGND VPWR VPWR _06983_ sky130_fd_sc_hd__nor2_1
X_26768_ clknet_leaf_4_clk_sys _00385_ net580 VGND VGND VPWR VPWR top0.cordic0.cos\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_16521_ _08602_ _08608_ VGND VGND VPWR VPWR _08609_ sky130_fd_sc_hd__xnor2_2
X_13733_ _05928_ _05943_ _05945_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__a21o_1
X_25719_ net74 _04931_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26699_ clknet_leaf_63_clk_sys _00316_ net648 VGND VGND VPWR VPWR top0.pid_d.prev_error\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_19240_ _11185_ _11186_ VGND VGND VPWR VPWR _11187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16452_ _08493_ _08540_ VGND VGND VPWR VPWR _08541_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_168_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13664_ _05848_ _05876_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_195_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15403_ _07489_ _07490_ _07501_ VGND VGND VPWR VPWR _07502_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19171_ net361 _11117_ _11124_ _10067_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__o211a_1
X_16383_ _08468_ _08469_ _08471_ _08312_ _08472_ VGND VGND VPWR VPWR _08473_ sky130_fd_sc_hd__o221a_1
XFILLER_0_112_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13595_ net66 _05626_ _05621_ _05640_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18122_ net328 net394 VGND VGND VPWR VPWR _10106_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15334_ net539 net472 VGND VGND VPWR VPWR _07433_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_60_clk_sys clknet_3_4__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_60_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_101_clk_sys clknet_3_0__leaf_clk_sys VGND VGND VPWR VPWR clknet_leaf_101_clk_sys
+ sky130_fd_sc_hd__clkbuf_16
X_18053_ _10009_ _10037_ VGND VGND VPWR VPWR _10038_ sky130_fd_sc_hd__xor2_1
X_15265_ _07355_ _07360_ _07363_ VGND VGND VPWR VPWR _07364_ sky130_fd_sc_hd__a21o_1
XANTENNA_4 _02367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17004_ _09057_ _09038_ top0.currT_r\[12\] _09039_ VGND VGND VPWR VPWR _09058_ sky130_fd_sc_hd__o2bb2a_1
X_14216_ _06330_ _06426_ _06329_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_151_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15196_ _07193_ _07191_ VGND VGND VPWR VPWR _07295_ sky130_fd_sc_hd__and2_1
X_14147_ _06244_ _06245_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__or2b_1
XFILLER_0_22_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14078_ _05530_ _05608_ _05609_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__or3_1
X_18955_ _10890_ _10857_ VGND VGND VPWR VPWR _10929_ sky130_fd_sc_hd__or2b_1
XFILLER_0_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17906_ _09823_ _09891_ VGND VGND VPWR VPWR _09893_ sky130_fd_sc_hd__or2_2
X_18886_ _10777_ _10783_ _10860_ _10255_ VGND VGND VPWR VPWR _10861_ sky130_fd_sc_hd__a2bb2o_2
X_17837_ _09812_ _09815_ VGND VGND VPWR VPWR _09824_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17768_ _09662_ _09682_ _09669_ VGND VGND VPWR VPWR _09755_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16719_ _08754_ _08777_ _08802_ _08750_ VGND VGND VPWR VPWR _08803_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19507_ _11037_ _11397_ _11080_ VGND VGND VPWR VPWR _11398_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17699_ _09635_ _09685_ VGND VGND VPWR VPWR _09686_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_202_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19438_ top0.pid_d.curr_int\[7\] top0.pid_d.prev_int\[7\] VGND VGND VPWR VPWR _11337_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19369_ net892 _11285_ _11288_ top0.pid_d.curr_error\[2\] VGND VGND VPWR VPWR _00312_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21400_ _00944_ _00945_ _00940_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__o21a_1
XFILLER_0_199_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22380_ _11674_ _01938_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21331_ _13171_ _13172_ VGND VGND VPWR VPWR _13173_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24050_ _03393_ _03397_ _03406_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21262_ _13016_ _13105_ VGND VGND VPWR VPWR _13106_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_23001_ _02345_ _02506_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20213_ _11550_ _12061_ VGND VGND VPWR VPWR _12062_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21193_ net213 _13035_ VGND VGND VPWR VPWR _13037_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20144_ _11983_ _11515_ _11997_ top0.cordic0.slte0.opA\[17\] _11649_ VGND VGND VPWR
+ VPWR _11999_ sky130_fd_sc_hd__a32o_1
X_24952_ _04268_ _04302_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__xnor2_4
X_20075_ net181 _11519_ VGND VGND VPWR VPWR _11936_ sky130_fd_sc_hd__nor2_2
X_23903_ _03249_ _03253_ _03255_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__a21o_1
X_24883_ _04212_ _04234_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_135_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26622_ clknet_leaf_25_clk_sys _00239_ net627 VGND VGND VPWR VPWR top0.matmul0.beta_pass\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_197_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_23834_ _03181_ _03191_ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_169_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26553_ clknet_leaf_49_clk_sys _00176_ net675 VGND VGND VPWR VPWR top0.pid_q.mult0.b\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_23765_ _03122_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__buf_6
X_20977_ net227 net219 VGND VGND VPWR VPWR _12824_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25504_ top0.matmul0.matmul_stage_inst.mult1\[8\] _04401_ _04829_ VGND VGND VPWR
+ VPWR _04838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22716_ _02262_ _02266_ _02180_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__a21oi_1
X_26484_ clknet_leaf_89_clk_sys _00115_ net604 VGND VGND VPWR VPWR top0.periodTop\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_23696_ net571 net574 top0.matmul0.matmul_stage_inst.f\[7\] VGND VGND VPWR VPWR _03054_
+ sky130_fd_sc_hd__o21a_4
XFILLER_0_48_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_25435_ _04726_ _04730_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_22647_ _02161_ _02160_ _02153_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_180_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13380_ _05584_ _05592_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__xnor2_1
X_25366_ top0.matmul0.matmul_stage_inst.mult2\[13\] _04710_ _03146_ VGND VGND VPWR
+ VPWR _04711_ sky130_fd_sc_hd__mux2_1
X_22578_ _02127_ _02132_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27105_ clknet_leaf_22_clk_sys _00722_ net608 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.a\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_24317_ _03132_ _03664_ _03133_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_69_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21529_ net143 net146 VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__or2b_1
X_25297_ _04510_ _04642_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__xor2_2
XFILLER_0_181_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15050_ _07145_ _07148_ VGND VGND VPWR VPWR _07149_ sky130_fd_sc_hd__xnor2_2
X_27036_ clknet_leaf_9_clk_sys _00653_ net594 VGND VGND VPWR VPWR top0.matmul0.matmul_stage_inst.e\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_24248_ _03540_ _03546_ _03548_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_160_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14001_ _05683_ _05894_ net24 VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__o21a_1
Xoutput6 net6 VGND VGND VPWR VPWR pwmC sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_24179_ _03478_ _03533_ _03489_ VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18740_ _10635_ _10640_ _10633_ VGND VGND VPWR VPWR _10717_ sky130_fd_sc_hd__o21a_1
X_15952_ _07907_ _07908_ _08046_ VGND VGND VPWR VPWR _08047_ sky130_fd_sc_hd__a21bo_1
X_14903_ spi0.data_packed\[59\] top0.kpq\[11\] _07064_ VGND VGND VPWR VPWR _07072_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18671_ _10631_ _10648_ VGND VGND VPWR VPWR _10649_ sky130_fd_sc_hd__xnor2_1
X_15883_ _07964_ _07978_ VGND VGND VPWR VPWR _07979_ sky130_fd_sc_hd__xnor2_1
X_17622_ net325 net424 VGND VGND VPWR VPWR _09609_ sky130_fd_sc_hd__nand2_2
X_14834_ _07008_ _07025_ _07026_ VGND VGND VPWR VPWR _07033_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17553_ net337 net425 VGND VGND VPWR VPWR _09540_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14765_ _06952_ _06966_ VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16504_ _08587_ _08591_ VGND VGND VPWR VPWR _08592_ sky130_fd_sc_hd__xnor2_2
X_13716_ net59 _05472_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__nand2_1
X_17484_ _09469_ _09470_ VGND VGND VPWR VPWR _09471_ sky130_fd_sc_hd__xor2_1
X_14696_ _06879_ _06898_ VGND VGND VPWR VPWR _06900_ sky130_fd_sc_hd__or2_1
X_19223_ _11121_ _11171_ _11125_ VGND VGND VPWR VPWR _11172_ sky130_fd_sc_hd__a21o_1
XFILLER_0_195_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16435_ _08436_ _08438_ _08434_ VGND VGND VPWR VPWR _08524_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_6_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13647_ _05803_ _05859_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_186_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19154_ net380 _11095_ _11112_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__a21o_1
X_16366_ _08444_ _08455_ VGND VGND VPWR VPWR _08456_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13578_ _05653_ _05655_ _05674_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__o21ba_1
X_18105_ _10031_ _10033_ _10029_ VGND VGND VPWR VPWR _10089_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_81_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15317_ _07362_ _07360_ VGND VGND VPWR VPWR _07416_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19085_ net371 _11056_ _11053_ _09965_ VGND VGND VPWR VPWR _11057_ sky130_fd_sc_hd__a22o_1
X_16297_ _08381_ _08387_ VGND VGND VPWR VPWR _08388_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18036_ _10015_ _10020_ VGND VGND VPWR VPWR _10021_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15248_ _07304_ _07319_ _07342_ VGND VGND VPWR VPWR _07347_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15179_ _07274_ _07277_ VGND VGND VPWR VPWR _07278_ sky130_fd_sc_hd__xnor2_2
Xfanout308 net309 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__buf_2
Xfanout319 top0.pid_d.mult0.b\[11\] VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19987_ _11852_ _11854_ VGND VGND VPWR VPWR _11855_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_197_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18938_ top0.pid_d.out\[11\] top0.pid_d.curr_int\[11\] VGND VGND VPWR VPWR _10913_
+ sky130_fd_sc_hd__nor2_1
.ends

