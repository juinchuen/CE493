module top (clk,
    pid_d_wen,
    pid_q_wen,
    pwmA_out,
    pwmB_out,
    pwmC_out,
    ready,
    rstb,
    valid,
    angle_in,
    currA_in,
    currB_in,
    currC_in,
    currT_in,
    periodTop,
    pid_d_addr,
    pid_d_data,
    pid_q_addr,
    pid_q_data);
 input clk;
 input pid_d_wen;
 input pid_q_wen;
 output pwmA_out;
 output pwmB_out;
 output pwmC_out;
 output ready;
 input rstb;
 input valid;
 input [15:0] angle_in;
 input [15:0] currA_in;
 input [15:0] currB_in;
 input [15:0] currC_in;
 input [15:0] currT_in;
 input [15:0] periodTop;
 input [15:0] pid_d_addr;
 input [15:0] pid_d_data;
 input [15:0] pid_q_addr;
 input [15:0] pid_q_data;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire clarke_done;
 wire \cordic0.cos[0] ;
 wire \cordic0.cos[10] ;
 wire \cordic0.cos[11] ;
 wire \cordic0.cos[12] ;
 wire \cordic0.cos[13] ;
 wire \cordic0.cos[1] ;
 wire \cordic0.cos[2] ;
 wire \cordic0.cos[3] ;
 wire \cordic0.cos[4] ;
 wire \cordic0.cos[5] ;
 wire \cordic0.cos[6] ;
 wire \cordic0.cos[7] ;
 wire \cordic0.cos[8] ;
 wire \cordic0.cos[9] ;
 wire \cordic0.domain[0] ;
 wire \cordic0.domain[1] ;
 wire \cordic0.gm0.iter[0] ;
 wire \cordic0.gm0.iter[1] ;
 wire \cordic0.gm0.iter[2] ;
 wire \cordic0.gm0.iter[3] ;
 wire \cordic0.gm0.iter[4] ;
 wire \cordic0.in_valid ;
 wire \cordic0.out_valid ;
 wire \cordic0.sin[0] ;
 wire \cordic0.sin[10] ;
 wire \cordic0.sin[11] ;
 wire \cordic0.sin[12] ;
 wire \cordic0.sin[13] ;
 wire \cordic0.sin[1] ;
 wire \cordic0.sin[2] ;
 wire \cordic0.sin[3] ;
 wire \cordic0.sin[4] ;
 wire \cordic0.sin[5] ;
 wire \cordic0.sin[6] ;
 wire \cordic0.sin[7] ;
 wire \cordic0.sin[8] ;
 wire \cordic0.sin[9] ;
 wire \cordic0.slte0.opA[0] ;
 wire \cordic0.slte0.opA[10] ;
 wire \cordic0.slte0.opA[11] ;
 wire \cordic0.slte0.opA[12] ;
 wire \cordic0.slte0.opA[13] ;
 wire \cordic0.slte0.opA[14] ;
 wire \cordic0.slte0.opA[15] ;
 wire \cordic0.slte0.opA[16] ;
 wire \cordic0.slte0.opA[17] ;
 wire \cordic0.slte0.opA[1] ;
 wire \cordic0.slte0.opA[2] ;
 wire \cordic0.slte0.opA[3] ;
 wire \cordic0.slte0.opA[4] ;
 wire \cordic0.slte0.opA[5] ;
 wire \cordic0.slte0.opA[6] ;
 wire \cordic0.slte0.opA[7] ;
 wire \cordic0.slte0.opA[8] ;
 wire \cordic0.slte0.opA[9] ;
 wire \cordic0.slte0.opB[10] ;
 wire \cordic0.slte0.opB[11] ;
 wire \cordic0.slte0.opB[12] ;
 wire \cordic0.slte0.opB[13] ;
 wire \cordic0.slte0.opB[14] ;
 wire \cordic0.slte0.opB[15] ;
 wire \cordic0.slte0.opB[2] ;
 wire \cordic0.slte0.opB[3] ;
 wire \cordic0.slte0.opB[4] ;
 wire \cordic0.slte0.opB[5] ;
 wire \cordic0.slte0.opB[6] ;
 wire \cordic0.slte0.opB[7] ;
 wire \cordic0.slte0.opB[8] ;
 wire \cordic0.slte0.opB[9] ;
 wire \cordic0.state[0] ;
 wire \cordic0.vec[0][0] ;
 wire \cordic0.vec[0][10] ;
 wire \cordic0.vec[0][11] ;
 wire \cordic0.vec[0][12] ;
 wire \cordic0.vec[0][13] ;
 wire \cordic0.vec[0][14] ;
 wire \cordic0.vec[0][15] ;
 wire \cordic0.vec[0][16] ;
 wire \cordic0.vec[0][17] ;
 wire \cordic0.vec[0][1] ;
 wire \cordic0.vec[0][2] ;
 wire \cordic0.vec[0][3] ;
 wire \cordic0.vec[0][4] ;
 wire \cordic0.vec[0][5] ;
 wire \cordic0.vec[0][6] ;
 wire \cordic0.vec[0][7] ;
 wire \cordic0.vec[0][8] ;
 wire \cordic0.vec[0][9] ;
 wire \cordic0.vec[1][0] ;
 wire \cordic0.vec[1][10] ;
 wire \cordic0.vec[1][11] ;
 wire \cordic0.vec[1][12] ;
 wire \cordic0.vec[1][13] ;
 wire \cordic0.vec[1][14] ;
 wire \cordic0.vec[1][15] ;
 wire \cordic0.vec[1][16] ;
 wire \cordic0.vec[1][17] ;
 wire \cordic0.vec[1][1] ;
 wire \cordic0.vec[1][2] ;
 wire \cordic0.vec[1][3] ;
 wire \cordic0.vec[1][4] ;
 wire \cordic0.vec[1][5] ;
 wire \cordic0.vec[1][6] ;
 wire \cordic0.vec[1][7] ;
 wire \cordic0.vec[1][8] ;
 wire \cordic0.vec[1][9] ;
 wire cordic_done;
 wire \matmul0.a[0] ;
 wire \matmul0.a[10] ;
 wire \matmul0.a[11] ;
 wire \matmul0.a[12] ;
 wire \matmul0.a[13] ;
 wire \matmul0.a[14] ;
 wire \matmul0.a[15] ;
 wire \matmul0.a[1] ;
 wire \matmul0.a[2] ;
 wire \matmul0.a[3] ;
 wire \matmul0.a[4] ;
 wire \matmul0.a[5] ;
 wire \matmul0.a[6] ;
 wire \matmul0.a[7] ;
 wire \matmul0.a[8] ;
 wire \matmul0.a[9] ;
 wire \matmul0.a_in[0] ;
 wire \matmul0.a_in[10] ;
 wire \matmul0.a_in[11] ;
 wire \matmul0.a_in[12] ;
 wire \matmul0.a_in[13] ;
 wire \matmul0.a_in[14] ;
 wire \matmul0.a_in[15] ;
 wire \matmul0.a_in[1] ;
 wire \matmul0.a_in[2] ;
 wire \matmul0.a_in[3] ;
 wire \matmul0.a_in[4] ;
 wire \matmul0.a_in[5] ;
 wire \matmul0.a_in[6] ;
 wire \matmul0.a_in[7] ;
 wire \matmul0.a_in[8] ;
 wire \matmul0.a_in[9] ;
 wire \matmul0.alpha_pass[0] ;
 wire \matmul0.alpha_pass[10] ;
 wire \matmul0.alpha_pass[11] ;
 wire \matmul0.alpha_pass[12] ;
 wire \matmul0.alpha_pass[13] ;
 wire \matmul0.alpha_pass[14] ;
 wire \matmul0.alpha_pass[15] ;
 wire \matmul0.alpha_pass[1] ;
 wire \matmul0.alpha_pass[2] ;
 wire \matmul0.alpha_pass[3] ;
 wire \matmul0.alpha_pass[4] ;
 wire \matmul0.alpha_pass[5] ;
 wire \matmul0.alpha_pass[6] ;
 wire \matmul0.alpha_pass[7] ;
 wire \matmul0.alpha_pass[8] ;
 wire \matmul0.alpha_pass[9] ;
 wire \matmul0.b[0] ;
 wire \matmul0.b[10] ;
 wire \matmul0.b[11] ;
 wire \matmul0.b[12] ;
 wire \matmul0.b[13] ;
 wire \matmul0.b[14] ;
 wire \matmul0.b[15] ;
 wire \matmul0.b[1] ;
 wire \matmul0.b[2] ;
 wire \matmul0.b[3] ;
 wire \matmul0.b[4] ;
 wire \matmul0.b[5] ;
 wire \matmul0.b[6] ;
 wire \matmul0.b[7] ;
 wire \matmul0.b[8] ;
 wire \matmul0.b[9] ;
 wire \matmul0.b_in[0] ;
 wire \matmul0.b_in[10] ;
 wire \matmul0.b_in[11] ;
 wire \matmul0.b_in[12] ;
 wire \matmul0.b_in[13] ;
 wire \matmul0.b_in[14] ;
 wire \matmul0.b_in[15] ;
 wire \matmul0.b_in[1] ;
 wire \matmul0.b_in[2] ;
 wire \matmul0.b_in[3] ;
 wire \matmul0.b_in[4] ;
 wire \matmul0.b_in[5] ;
 wire \matmul0.b_in[6] ;
 wire \matmul0.b_in[7] ;
 wire \matmul0.b_in[8] ;
 wire \matmul0.b_in[9] ;
 wire \matmul0.beta_pass[0] ;
 wire \matmul0.beta_pass[10] ;
 wire \matmul0.beta_pass[11] ;
 wire \matmul0.beta_pass[12] ;
 wire \matmul0.beta_pass[13] ;
 wire \matmul0.beta_pass[14] ;
 wire \matmul0.beta_pass[15] ;
 wire \matmul0.beta_pass[1] ;
 wire \matmul0.beta_pass[2] ;
 wire \matmul0.beta_pass[3] ;
 wire \matmul0.beta_pass[4] ;
 wire \matmul0.beta_pass[5] ;
 wire \matmul0.beta_pass[6] ;
 wire \matmul0.beta_pass[7] ;
 wire \matmul0.beta_pass[8] ;
 wire \matmul0.beta_pass[9] ;
 wire \matmul0.cos[0] ;
 wire \matmul0.cos[10] ;
 wire \matmul0.cos[11] ;
 wire \matmul0.cos[12] ;
 wire \matmul0.cos[13] ;
 wire \matmul0.cos[1] ;
 wire \matmul0.cos[2] ;
 wire \matmul0.cos[3] ;
 wire \matmul0.cos[4] ;
 wire \matmul0.cos[5] ;
 wire \matmul0.cos[6] ;
 wire \matmul0.cos[7] ;
 wire \matmul0.cos[8] ;
 wire \matmul0.cos[9] ;
 wire \matmul0.done_pass ;
 wire \matmul0.matmul_stage_inst.a[0] ;
 wire \matmul0.matmul_stage_inst.a[10] ;
 wire \matmul0.matmul_stage_inst.a[11] ;
 wire \matmul0.matmul_stage_inst.a[12] ;
 wire \matmul0.matmul_stage_inst.a[13] ;
 wire \matmul0.matmul_stage_inst.a[14] ;
 wire \matmul0.matmul_stage_inst.a[1] ;
 wire \matmul0.matmul_stage_inst.a[2] ;
 wire \matmul0.matmul_stage_inst.a[3] ;
 wire \matmul0.matmul_stage_inst.a[4] ;
 wire \matmul0.matmul_stage_inst.a[5] ;
 wire \matmul0.matmul_stage_inst.a[6] ;
 wire \matmul0.matmul_stage_inst.a[7] ;
 wire \matmul0.matmul_stage_inst.a[8] ;
 wire \matmul0.matmul_stage_inst.a[9] ;
 wire \matmul0.matmul_stage_inst.b[0] ;
 wire \matmul0.matmul_stage_inst.b[10] ;
 wire \matmul0.matmul_stage_inst.b[11] ;
 wire \matmul0.matmul_stage_inst.b[12] ;
 wire \matmul0.matmul_stage_inst.b[13] ;
 wire \matmul0.matmul_stage_inst.b[14] ;
 wire \matmul0.matmul_stage_inst.b[15] ;
 wire \matmul0.matmul_stage_inst.b[1] ;
 wire \matmul0.matmul_stage_inst.b[2] ;
 wire \matmul0.matmul_stage_inst.b[3] ;
 wire \matmul0.matmul_stage_inst.b[4] ;
 wire \matmul0.matmul_stage_inst.b[5] ;
 wire \matmul0.matmul_stage_inst.b[6] ;
 wire \matmul0.matmul_stage_inst.b[7] ;
 wire \matmul0.matmul_stage_inst.b[8] ;
 wire \matmul0.matmul_stage_inst.b[9] ;
 wire \matmul0.matmul_stage_inst.c[10] ;
 wire \matmul0.matmul_stage_inst.c[11] ;
 wire \matmul0.matmul_stage_inst.c[12] ;
 wire \matmul0.matmul_stage_inst.c[13] ;
 wire \matmul0.matmul_stage_inst.c[14] ;
 wire \matmul0.matmul_stage_inst.c[15] ;
 wire \matmul0.matmul_stage_inst.c[1] ;
 wire \matmul0.matmul_stage_inst.c[2] ;
 wire \matmul0.matmul_stage_inst.c[3] ;
 wire \matmul0.matmul_stage_inst.c[4] ;
 wire \matmul0.matmul_stage_inst.c[5] ;
 wire \matmul0.matmul_stage_inst.c[6] ;
 wire \matmul0.matmul_stage_inst.c[7] ;
 wire \matmul0.matmul_stage_inst.c[8] ;
 wire \matmul0.matmul_stage_inst.c[9] ;
 wire \matmul0.matmul_stage_inst.d[0] ;
 wire \matmul0.matmul_stage_inst.d[10] ;
 wire \matmul0.matmul_stage_inst.d[11] ;
 wire \matmul0.matmul_stage_inst.d[12] ;
 wire \matmul0.matmul_stage_inst.d[13] ;
 wire \matmul0.matmul_stage_inst.d[1] ;
 wire \matmul0.matmul_stage_inst.d[2] ;
 wire \matmul0.matmul_stage_inst.d[4] ;
 wire \matmul0.matmul_stage_inst.d[5] ;
 wire \matmul0.matmul_stage_inst.d[6] ;
 wire \matmul0.matmul_stage_inst.d[7] ;
 wire \matmul0.matmul_stage_inst.d[8] ;
 wire \matmul0.matmul_stage_inst.d[9] ;
 wire \matmul0.matmul_stage_inst.e[0] ;
 wire \matmul0.matmul_stage_inst.e[10] ;
 wire \matmul0.matmul_stage_inst.e[11] ;
 wire \matmul0.matmul_stage_inst.e[12] ;
 wire \matmul0.matmul_stage_inst.e[13] ;
 wire \matmul0.matmul_stage_inst.e[14] ;
 wire \matmul0.matmul_stage_inst.e[15] ;
 wire \matmul0.matmul_stage_inst.e[1] ;
 wire \matmul0.matmul_stage_inst.e[2] ;
 wire \matmul0.matmul_stage_inst.e[3] ;
 wire \matmul0.matmul_stage_inst.e[4] ;
 wire \matmul0.matmul_stage_inst.e[5] ;
 wire \matmul0.matmul_stage_inst.e[6] ;
 wire \matmul0.matmul_stage_inst.e[7] ;
 wire \matmul0.matmul_stage_inst.e[8] ;
 wire \matmul0.matmul_stage_inst.e[9] ;
 wire \matmul0.matmul_stage_inst.f[0] ;
 wire \matmul0.matmul_stage_inst.f[10] ;
 wire \matmul0.matmul_stage_inst.f[11] ;
 wire \matmul0.matmul_stage_inst.f[12] ;
 wire \matmul0.matmul_stage_inst.f[13] ;
 wire \matmul0.matmul_stage_inst.f[14] ;
 wire \matmul0.matmul_stage_inst.f[15] ;
 wire \matmul0.matmul_stage_inst.f[1] ;
 wire \matmul0.matmul_stage_inst.f[2] ;
 wire \matmul0.matmul_stage_inst.f[3] ;
 wire \matmul0.matmul_stage_inst.f[4] ;
 wire \matmul0.matmul_stage_inst.f[5] ;
 wire \matmul0.matmul_stage_inst.f[6] ;
 wire \matmul0.matmul_stage_inst.f[7] ;
 wire \matmul0.matmul_stage_inst.f[8] ;
 wire \matmul0.matmul_stage_inst.f[9] ;
 wire \matmul0.matmul_stage_inst.mult1[0] ;
 wire \matmul0.matmul_stage_inst.mult1[10] ;
 wire \matmul0.matmul_stage_inst.mult1[11] ;
 wire \matmul0.matmul_stage_inst.mult1[12] ;
 wire \matmul0.matmul_stage_inst.mult1[13] ;
 wire \matmul0.matmul_stage_inst.mult1[14] ;
 wire \matmul0.matmul_stage_inst.mult1[15] ;
 wire \matmul0.matmul_stage_inst.mult1[1] ;
 wire \matmul0.matmul_stage_inst.mult1[2] ;
 wire \matmul0.matmul_stage_inst.mult1[3] ;
 wire \matmul0.matmul_stage_inst.mult1[4] ;
 wire \matmul0.matmul_stage_inst.mult1[5] ;
 wire \matmul0.matmul_stage_inst.mult1[6] ;
 wire \matmul0.matmul_stage_inst.mult1[7] ;
 wire \matmul0.matmul_stage_inst.mult1[8] ;
 wire \matmul0.matmul_stage_inst.mult1[9] ;
 wire \matmul0.matmul_stage_inst.mult2[0] ;
 wire \matmul0.matmul_stage_inst.mult2[10] ;
 wire \matmul0.matmul_stage_inst.mult2[11] ;
 wire \matmul0.matmul_stage_inst.mult2[12] ;
 wire \matmul0.matmul_stage_inst.mult2[13] ;
 wire \matmul0.matmul_stage_inst.mult2[14] ;
 wire \matmul0.matmul_stage_inst.mult2[15] ;
 wire \matmul0.matmul_stage_inst.mult2[1] ;
 wire \matmul0.matmul_stage_inst.mult2[2] ;
 wire \matmul0.matmul_stage_inst.mult2[3] ;
 wire \matmul0.matmul_stage_inst.mult2[4] ;
 wire \matmul0.matmul_stage_inst.mult2[5] ;
 wire \matmul0.matmul_stage_inst.mult2[6] ;
 wire \matmul0.matmul_stage_inst.mult2[7] ;
 wire \matmul0.matmul_stage_inst.mult2[8] ;
 wire \matmul0.matmul_stage_inst.mult2[9] ;
 wire \matmul0.matmul_stage_inst.start ;
 wire \matmul0.matmul_stage_inst.state[0] ;
 wire \matmul0.matmul_stage_inst.state[1] ;
 wire \matmul0.matmul_stage_inst.state[2] ;
 wire \matmul0.matmul_stage_inst.state[4] ;
 wire \matmul0.matmul_stage_inst.state[5] ;
 wire \matmul0.matmul_stage_inst.state[6] ;
 wire \matmul0.op[0] ;
 wire \matmul0.op[1] ;
 wire \matmul0.op_in[0] ;
 wire \matmul0.op_in[1] ;
 wire \matmul0.sin[0] ;
 wire \matmul0.sin[10] ;
 wire \matmul0.sin[11] ;
 wire \matmul0.sin[12] ;
 wire \matmul0.sin[13] ;
 wire \matmul0.sin[1] ;
 wire \matmul0.sin[2] ;
 wire \matmul0.sin[3] ;
 wire \matmul0.sin[4] ;
 wire \matmul0.sin[5] ;
 wire \matmul0.sin[6] ;
 wire \matmul0.sin[7] ;
 wire \matmul0.sin[8] ;
 wire \matmul0.sin[9] ;
 wire \matmul0.start ;
 wire \matmul0.state[0] ;
 wire \matmul0.state[1] ;
 wire \pid_d.curr_error[0] ;
 wire \pid_d.curr_error[10] ;
 wire \pid_d.curr_error[11] ;
 wire \pid_d.curr_error[12] ;
 wire \pid_d.curr_error[13] ;
 wire \pid_d.curr_error[14] ;
 wire \pid_d.curr_error[15] ;
 wire \pid_d.curr_error[1] ;
 wire \pid_d.curr_error[2] ;
 wire \pid_d.curr_error[3] ;
 wire \pid_d.curr_error[4] ;
 wire \pid_d.curr_error[5] ;
 wire \pid_d.curr_error[6] ;
 wire \pid_d.curr_error[7] ;
 wire \pid_d.curr_error[8] ;
 wire \pid_d.curr_error[9] ;
 wire \pid_d.curr_int[0] ;
 wire \pid_d.curr_int[10] ;
 wire \pid_d.curr_int[11] ;
 wire \pid_d.curr_int[12] ;
 wire \pid_d.curr_int[13] ;
 wire \pid_d.curr_int[14] ;
 wire \pid_d.curr_int[15] ;
 wire \pid_d.curr_int[1] ;
 wire \pid_d.curr_int[2] ;
 wire \pid_d.curr_int[3] ;
 wire \pid_d.curr_int[4] ;
 wire \pid_d.curr_int[5] ;
 wire \pid_d.curr_int[6] ;
 wire \pid_d.curr_int[7] ;
 wire \pid_d.curr_int[8] ;
 wire \pid_d.curr_int[9] ;
 wire \pid_d.iterate_enable ;
 wire \pid_d.ki[0] ;
 wire \pid_d.ki[10] ;
 wire \pid_d.ki[11] ;
 wire \pid_d.ki[12] ;
 wire \pid_d.ki[13] ;
 wire \pid_d.ki[14] ;
 wire \pid_d.ki[15] ;
 wire \pid_d.ki[1] ;
 wire \pid_d.ki[2] ;
 wire \pid_d.ki[3] ;
 wire \pid_d.ki[4] ;
 wire \pid_d.ki[5] ;
 wire \pid_d.ki[6] ;
 wire \pid_d.ki[7] ;
 wire \pid_d.ki[8] ;
 wire \pid_d.ki[9] ;
 wire \pid_d.kp[0] ;
 wire \pid_d.kp[10] ;
 wire \pid_d.kp[11] ;
 wire \pid_d.kp[12] ;
 wire \pid_d.kp[13] ;
 wire \pid_d.kp[14] ;
 wire \pid_d.kp[15] ;
 wire \pid_d.kp[1] ;
 wire \pid_d.kp[2] ;
 wire \pid_d.kp[3] ;
 wire \pid_d.kp[4] ;
 wire \pid_d.kp[5] ;
 wire \pid_d.kp[6] ;
 wire \pid_d.kp[7] ;
 wire \pid_d.kp[8] ;
 wire \pid_d.kp[9] ;
 wire \pid_d.mult0.a[0] ;
 wire \pid_d.mult0.a[10] ;
 wire \pid_d.mult0.a[11] ;
 wire \pid_d.mult0.a[12] ;
 wire \pid_d.mult0.a[13] ;
 wire \pid_d.mult0.a[14] ;
 wire \pid_d.mult0.a[15] ;
 wire \pid_d.mult0.a[1] ;
 wire \pid_d.mult0.a[2] ;
 wire \pid_d.mult0.a[3] ;
 wire \pid_d.mult0.a[4] ;
 wire \pid_d.mult0.a[5] ;
 wire \pid_d.mult0.a[6] ;
 wire \pid_d.mult0.a[7] ;
 wire \pid_d.mult0.a[8] ;
 wire \pid_d.mult0.a[9] ;
 wire \pid_d.mult0.b[0] ;
 wire \pid_d.mult0.b[10] ;
 wire \pid_d.mult0.b[11] ;
 wire \pid_d.mult0.b[12] ;
 wire \pid_d.mult0.b[13] ;
 wire \pid_d.mult0.b[14] ;
 wire \pid_d.mult0.b[15] ;
 wire \pid_d.mult0.b[1] ;
 wire \pid_d.mult0.b[2] ;
 wire \pid_d.mult0.b[3] ;
 wire \pid_d.mult0.b[4] ;
 wire \pid_d.mult0.b[5] ;
 wire \pid_d.mult0.b[6] ;
 wire \pid_d.mult0.b[7] ;
 wire \pid_d.mult0.b[8] ;
 wire \pid_d.mult0.b[9] ;
 wire \pid_d.out[0] ;
 wire \pid_d.out[10] ;
 wire \pid_d.out[11] ;
 wire \pid_d.out[12] ;
 wire \pid_d.out[13] ;
 wire \pid_d.out[14] ;
 wire \pid_d.out[15] ;
 wire \pid_d.out[1] ;
 wire \pid_d.out[2] ;
 wire \pid_d.out[3] ;
 wire \pid_d.out[4] ;
 wire \pid_d.out[5] ;
 wire \pid_d.out[6] ;
 wire \pid_d.out[7] ;
 wire \pid_d.out[8] ;
 wire \pid_d.out[9] ;
 wire \pid_d.out_valid ;
 wire \pid_d.prev_error[0] ;
 wire \pid_d.prev_error[10] ;
 wire \pid_d.prev_error[11] ;
 wire \pid_d.prev_error[12] ;
 wire \pid_d.prev_error[13] ;
 wire \pid_d.prev_error[14] ;
 wire \pid_d.prev_error[15] ;
 wire \pid_d.prev_error[1] ;
 wire \pid_d.prev_error[2] ;
 wire \pid_d.prev_error[3] ;
 wire \pid_d.prev_error[4] ;
 wire \pid_d.prev_error[5] ;
 wire \pid_d.prev_error[6] ;
 wire \pid_d.prev_error[7] ;
 wire \pid_d.prev_error[8] ;
 wire \pid_d.prev_error[9] ;
 wire \pid_d.prev_int[0] ;
 wire \pid_d.prev_int[10] ;
 wire \pid_d.prev_int[11] ;
 wire \pid_d.prev_int[12] ;
 wire \pid_d.prev_int[13] ;
 wire \pid_d.prev_int[14] ;
 wire \pid_d.prev_int[15] ;
 wire \pid_d.prev_int[1] ;
 wire \pid_d.prev_int[2] ;
 wire \pid_d.prev_int[3] ;
 wire \pid_d.prev_int[4] ;
 wire \pid_d.prev_int[5] ;
 wire \pid_d.prev_int[6] ;
 wire \pid_d.prev_int[7] ;
 wire \pid_d.prev_int[8] ;
 wire \pid_d.prev_int[9] ;
 wire \pid_d.state[0] ;
 wire \pid_d.state[1] ;
 wire \pid_d.state[2] ;
 wire \pid_d.state[3] ;
 wire \pid_d.state[4] ;
 wire \pid_d.state[5] ;
 wire \pid_q.curr_error[0] ;
 wire \pid_q.curr_error[10] ;
 wire \pid_q.curr_error[11] ;
 wire \pid_q.curr_error[12] ;
 wire \pid_q.curr_error[13] ;
 wire \pid_q.curr_error[14] ;
 wire \pid_q.curr_error[15] ;
 wire \pid_q.curr_error[1] ;
 wire \pid_q.curr_error[2] ;
 wire \pid_q.curr_error[3] ;
 wire \pid_q.curr_error[4] ;
 wire \pid_q.curr_error[5] ;
 wire \pid_q.curr_error[6] ;
 wire \pid_q.curr_error[7] ;
 wire \pid_q.curr_error[8] ;
 wire \pid_q.curr_error[9] ;
 wire \pid_q.curr_int[0] ;
 wire \pid_q.curr_int[10] ;
 wire \pid_q.curr_int[11] ;
 wire \pid_q.curr_int[12] ;
 wire \pid_q.curr_int[13] ;
 wire \pid_q.curr_int[14] ;
 wire \pid_q.curr_int[15] ;
 wire \pid_q.curr_int[1] ;
 wire \pid_q.curr_int[2] ;
 wire \pid_q.curr_int[3] ;
 wire \pid_q.curr_int[4] ;
 wire \pid_q.curr_int[5] ;
 wire \pid_q.curr_int[6] ;
 wire \pid_q.curr_int[7] ;
 wire \pid_q.curr_int[8] ;
 wire \pid_q.curr_int[9] ;
 wire \pid_q.ki[0] ;
 wire \pid_q.ki[10] ;
 wire \pid_q.ki[11] ;
 wire \pid_q.ki[12] ;
 wire \pid_q.ki[13] ;
 wire \pid_q.ki[14] ;
 wire \pid_q.ki[15] ;
 wire \pid_q.ki[1] ;
 wire \pid_q.ki[2] ;
 wire \pid_q.ki[3] ;
 wire \pid_q.ki[4] ;
 wire \pid_q.ki[5] ;
 wire \pid_q.ki[6] ;
 wire \pid_q.ki[7] ;
 wire \pid_q.ki[8] ;
 wire \pid_q.ki[9] ;
 wire \pid_q.kp[0] ;
 wire \pid_q.kp[10] ;
 wire \pid_q.kp[11] ;
 wire \pid_q.kp[12] ;
 wire \pid_q.kp[13] ;
 wire \pid_q.kp[14] ;
 wire \pid_q.kp[15] ;
 wire \pid_q.kp[1] ;
 wire \pid_q.kp[2] ;
 wire \pid_q.kp[3] ;
 wire \pid_q.kp[4] ;
 wire \pid_q.kp[5] ;
 wire \pid_q.kp[6] ;
 wire \pid_q.kp[7] ;
 wire \pid_q.kp[8] ;
 wire \pid_q.kp[9] ;
 wire \pid_q.mult0.a[0] ;
 wire \pid_q.mult0.a[10] ;
 wire \pid_q.mult0.a[11] ;
 wire \pid_q.mult0.a[12] ;
 wire \pid_q.mult0.a[13] ;
 wire \pid_q.mult0.a[14] ;
 wire \pid_q.mult0.a[15] ;
 wire \pid_q.mult0.a[1] ;
 wire \pid_q.mult0.a[2] ;
 wire \pid_q.mult0.a[3] ;
 wire \pid_q.mult0.a[4] ;
 wire \pid_q.mult0.a[5] ;
 wire \pid_q.mult0.a[6] ;
 wire \pid_q.mult0.a[7] ;
 wire \pid_q.mult0.a[8] ;
 wire \pid_q.mult0.a[9] ;
 wire \pid_q.mult0.b[0] ;
 wire \pid_q.mult0.b[10] ;
 wire \pid_q.mult0.b[11] ;
 wire \pid_q.mult0.b[12] ;
 wire \pid_q.mult0.b[13] ;
 wire \pid_q.mult0.b[14] ;
 wire \pid_q.mult0.b[15] ;
 wire \pid_q.mult0.b[1] ;
 wire \pid_q.mult0.b[2] ;
 wire \pid_q.mult0.b[3] ;
 wire \pid_q.mult0.b[4] ;
 wire \pid_q.mult0.b[5] ;
 wire \pid_q.mult0.b[6] ;
 wire \pid_q.mult0.b[7] ;
 wire \pid_q.mult0.b[8] ;
 wire \pid_q.mult0.b[9] ;
 wire \pid_q.out[0] ;
 wire \pid_q.out[10] ;
 wire \pid_q.out[11] ;
 wire \pid_q.out[12] ;
 wire \pid_q.out[13] ;
 wire \pid_q.out[14] ;
 wire \pid_q.out[15] ;
 wire \pid_q.out[1] ;
 wire \pid_q.out[2] ;
 wire \pid_q.out[3] ;
 wire \pid_q.out[4] ;
 wire \pid_q.out[5] ;
 wire \pid_q.out[6] ;
 wire \pid_q.out[7] ;
 wire \pid_q.out[8] ;
 wire \pid_q.out[9] ;
 wire \pid_q.prev_error[0] ;
 wire \pid_q.prev_error[10] ;
 wire \pid_q.prev_error[11] ;
 wire \pid_q.prev_error[12] ;
 wire \pid_q.prev_error[13] ;
 wire \pid_q.prev_error[14] ;
 wire \pid_q.prev_error[15] ;
 wire \pid_q.prev_error[1] ;
 wire \pid_q.prev_error[2] ;
 wire \pid_q.prev_error[3] ;
 wire \pid_q.prev_error[4] ;
 wire \pid_q.prev_error[5] ;
 wire \pid_q.prev_error[6] ;
 wire \pid_q.prev_error[7] ;
 wire \pid_q.prev_error[8] ;
 wire \pid_q.prev_error[9] ;
 wire \pid_q.prev_int[0] ;
 wire \pid_q.prev_int[10] ;
 wire \pid_q.prev_int[11] ;
 wire \pid_q.prev_int[12] ;
 wire \pid_q.prev_int[13] ;
 wire \pid_q.prev_int[14] ;
 wire \pid_q.prev_int[15] ;
 wire \pid_q.prev_int[1] ;
 wire \pid_q.prev_int[2] ;
 wire \pid_q.prev_int[3] ;
 wire \pid_q.prev_int[4] ;
 wire \pid_q.prev_int[5] ;
 wire \pid_q.prev_int[6] ;
 wire \pid_q.prev_int[7] ;
 wire \pid_q.prev_int[8] ;
 wire \pid_q.prev_int[9] ;
 wire \pid_q.state[0] ;
 wire \pid_q.state[1] ;
 wire \pid_q.state[2] ;
 wire \pid_q.state[3] ;
 wire \pid_q.state[4] ;
 wire \pid_q.state[5] ;
 wire \pid_q.target[0] ;
 wire \pid_q.target[10] ;
 wire \pid_q.target[11] ;
 wire \pid_q.target[12] ;
 wire \pid_q.target[13] ;
 wire \pid_q.target[14] ;
 wire \pid_q.target[15] ;
 wire \pid_q.target[1] ;
 wire \pid_q.target[2] ;
 wire \pid_q.target[3] ;
 wire \pid_q.target[4] ;
 wire \pid_q.target[5] ;
 wire \pid_q.target[6] ;
 wire \pid_q.target[7] ;
 wire \pid_q.target[8] ;
 wire \pid_q.target[9] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \svm0.calc_ready ;
 wire \svm0.counter[0] ;
 wire \svm0.counter[10] ;
 wire \svm0.counter[11] ;
 wire \svm0.counter[12] ;
 wire \svm0.counter[13] ;
 wire \svm0.counter[14] ;
 wire \svm0.counter[15] ;
 wire \svm0.counter[1] ;
 wire \svm0.counter[2] ;
 wire \svm0.counter[3] ;
 wire \svm0.counter[4] ;
 wire \svm0.counter[5] ;
 wire \svm0.counter[6] ;
 wire \svm0.counter[7] ;
 wire \svm0.counter[8] ;
 wire \svm0.counter[9] ;
 wire \svm0.delta[0] ;
 wire \svm0.delta[10] ;
 wire \svm0.delta[11] ;
 wire \svm0.delta[12] ;
 wire \svm0.delta[13] ;
 wire \svm0.delta[14] ;
 wire \svm0.delta[15] ;
 wire \svm0.delta[1] ;
 wire \svm0.delta[2] ;
 wire \svm0.delta[3] ;
 wire \svm0.delta[4] ;
 wire \svm0.delta[5] ;
 wire \svm0.delta[6] ;
 wire \svm0.delta[7] ;
 wire \svm0.delta[8] ;
 wire \svm0.delta[9] ;
 wire \svm0.in_valid ;
 wire \svm0.periodTop[0] ;
 wire \svm0.periodTop[10] ;
 wire \svm0.periodTop[11] ;
 wire \svm0.periodTop[12] ;
 wire \svm0.periodTop[13] ;
 wire \svm0.periodTop[14] ;
 wire \svm0.periodTop[15] ;
 wire \svm0.periodTop[1] ;
 wire \svm0.periodTop[2] ;
 wire \svm0.periodTop[3] ;
 wire \svm0.periodTop[4] ;
 wire \svm0.periodTop[5] ;
 wire \svm0.periodTop[6] ;
 wire \svm0.periodTop[7] ;
 wire \svm0.periodTop[8] ;
 wire \svm0.periodTop[9] ;
 wire \svm0.ready ;
 wire \svm0.rising ;
 wire \svm0.state[0] ;
 wire \svm0.state[1] ;
 wire \svm0.state[2] ;
 wire \svm0.tA[0] ;
 wire \svm0.tA[10] ;
 wire \svm0.tA[11] ;
 wire \svm0.tA[12] ;
 wire \svm0.tA[13] ;
 wire \svm0.tA[14] ;
 wire \svm0.tA[15] ;
 wire \svm0.tA[1] ;
 wire \svm0.tA[2] ;
 wire \svm0.tA[3] ;
 wire \svm0.tA[4] ;
 wire \svm0.tA[5] ;
 wire \svm0.tA[6] ;
 wire \svm0.tA[7] ;
 wire \svm0.tA[8] ;
 wire \svm0.tA[9] ;
 wire \svm0.tB[0] ;
 wire \svm0.tB[10] ;
 wire \svm0.tB[11] ;
 wire \svm0.tB[12] ;
 wire \svm0.tB[13] ;
 wire \svm0.tB[14] ;
 wire \svm0.tB[15] ;
 wire \svm0.tB[1] ;
 wire \svm0.tB[2] ;
 wire \svm0.tB[3] ;
 wire \svm0.tB[4] ;
 wire \svm0.tB[5] ;
 wire \svm0.tB[6] ;
 wire \svm0.tB[7] ;
 wire \svm0.tB[8] ;
 wire \svm0.tB[9] ;
 wire \svm0.tC[0] ;
 wire \svm0.tC[10] ;
 wire \svm0.tC[11] ;
 wire \svm0.tC[12] ;
 wire \svm0.tC[13] ;
 wire \svm0.tC[14] ;
 wire \svm0.tC[15] ;
 wire \svm0.tC[1] ;
 wire \svm0.tC[2] ;
 wire \svm0.tC[3] ;
 wire \svm0.tC[4] ;
 wire \svm0.tC[5] ;
 wire \svm0.tC[6] ;
 wire \svm0.tC[7] ;
 wire \svm0.tC[8] ;
 wire \svm0.tC[9] ;
 wire \svm0.vC[0] ;
 wire \svm0.vC[10] ;
 wire \svm0.vC[11] ;
 wire \svm0.vC[12] ;
 wire \svm0.vC[13] ;
 wire \svm0.vC[14] ;
 wire \svm0.vC[15] ;
 wire \svm0.vC[1] ;
 wire \svm0.vC[2] ;
 wire \svm0.vC[3] ;
 wire \svm0.vC[4] ;
 wire \svm0.vC[5] ;
 wire \svm0.vC[6] ;
 wire \svm0.vC[7] ;
 wire \svm0.vC[8] ;
 wire \svm0.vC[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4363;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4409;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net4440;
 wire net4441;
 wire net4442;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net4540;
 wire net4541;
 wire net4542;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net5349;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;
 wire net5389;
 wire net5390;
 wire net5391;
 wire net5392;
 wire net5393;
 wire net5394;
 wire net5395;
 wire net5396;
 wire net5397;
 wire net5398;
 wire net5399;
 wire net5400;
 wire net5401;
 wire net5402;
 wire net5403;
 wire net5404;
 wire net5405;
 wire net5406;
 wire net5407;
 wire net5408;
 wire net5409;
 wire net5410;
 wire net5411;
 wire net5412;
 wire net5413;
 wire net5414;
 wire net5415;
 wire net5416;
 wire net5417;
 wire net5418;
 wire net5419;
 wire net5420;
 wire net5421;
 wire net5422;
 wire net5423;
 wire net5424;
 wire net5425;
 wire net5426;
 wire net5427;
 wire net5428;
 wire net5429;
 wire net5430;
 wire net5431;
 wire net5432;
 wire net5433;
 wire net5434;
 wire net5435;
 wire net5436;
 wire net5437;
 wire net5438;
 wire net5439;
 wire net5440;
 wire net5441;
 wire net5442;
 wire net5443;
 wire net5444;
 wire net5445;
 wire net5446;
 wire net5447;
 wire net5448;
 wire net5449;
 wire net5450;
 wire net5451;
 wire net5452;
 wire net5453;
 wire net5454;
 wire net5455;
 wire net5456;
 wire net5457;
 wire net5458;
 wire net5459;
 wire net5460;
 wire net5461;
 wire net5462;
 wire net5463;
 wire net5464;
 wire net5465;
 wire net5466;
 wire net5467;
 wire net5468;
 wire net5469;
 wire net5470;
 wire net5471;
 wire net5472;
 wire net5473;
 wire net5474;
 wire net5475;
 wire net5476;
 wire net5477;
 wire net5478;
 wire net5479;
 wire net5480;
 wire net5481;
 wire net5482;
 wire net5483;
 wire net5484;
 wire net5485;
 wire net5486;
 wire net5487;
 wire net5488;
 wire net5489;
 wire net5490;
 wire net5491;
 wire net5492;
 wire net5493;
 wire net5494;
 wire net5495;
 wire net5496;
 wire net5497;
 wire net5498;
 wire net5499;
 wire net5500;
 wire net5501;
 wire net5502;
 wire net5503;
 wire net5504;
 wire net5505;
 wire net5506;
 wire net5507;
 wire net5508;
 wire net5509;
 wire net5510;
 wire net5511;
 wire net5512;
 wire net5513;
 wire net5514;
 wire net5515;
 wire net5516;
 wire net5517;
 wire net5518;
 wire net5519;
 wire net5520;
 wire net5521;
 wire net5522;
 wire net5523;
 wire net5524;
 wire net5525;
 wire net5526;
 wire net5527;
 wire net5528;
 wire net5529;
 wire net5530;
 wire net5531;
 wire net5532;
 wire net5533;
 wire net5534;
 wire net5535;
 wire net5536;
 wire net5537;
 wire net5538;
 wire net5539;
 wire net5540;
 wire net5541;
 wire net5542;
 wire net5543;
 wire net5544;
 wire net5545;
 wire net5546;
 wire net5547;
 wire net5548;
 wire net5549;
 wire net5550;
 wire net5551;
 wire net5552;
 wire net5553;
 wire net5554;
 wire net5555;
 wire net5556;
 wire net5557;
 wire net5558;
 wire net5559;
 wire net5560;
 wire net5561;
 wire net5562;
 wire net5563;
 wire net5564;
 wire net5565;
 wire net5566;
 wire net5567;
 wire net5568;
 wire net5569;
 wire net5570;
 wire net5571;
 wire net5572;
 wire net5573;
 wire net5574;
 wire net5575;
 wire net5576;
 wire net5577;
 wire net5578;
 wire net5579;
 wire net5580;
 wire net5581;
 wire net5582;
 wire net5583;
 wire net5584;
 wire net5585;
 wire net5586;
 wire net5587;
 wire net5588;
 wire net5589;
 wire net5590;
 wire net5591;
 wire net5592;
 wire net5593;
 wire net5594;
 wire net5595;
 wire net5596;
 wire net5597;
 wire net5598;
 wire net5599;
 wire net5600;
 wire net5601;
 wire net5602;
 wire net5603;
 wire net5604;
 wire net5605;
 wire net5606;
 wire net5607;
 wire net5608;
 wire net5609;
 wire net5610;
 wire net5611;
 wire net5612;
 wire net5613;
 wire net5614;
 wire net5615;
 wire net5616;
 wire net5617;
 wire net5618;
 wire net5619;
 wire net5620;
 wire net5621;
 wire net5622;
 wire net5623;
 wire net5624;
 wire net5625;
 wire net5626;
 wire net5627;
 wire net5628;
 wire net5629;
 wire net5630;
 wire net5631;
 wire net5632;
 wire net5633;
 wire net5634;
 wire net5635;
 wire net5636;
 wire net5637;
 wire net5638;
 wire net5639;
 wire net5640;
 wire net5641;
 wire net5642;
 wire net5643;
 wire net5644;
 wire net5645;
 wire net5646;
 wire net5647;
 wire net5648;
 wire net5649;
 wire net5650;
 wire net5651;
 wire net5652;
 wire net5653;
 wire net5654;
 wire net5655;
 wire net5656;
 wire net5657;
 wire net5658;
 wire net5659;
 wire net5660;
 wire net5661;
 wire net5662;
 wire net5663;
 wire net5664;
 wire net5665;
 wire net5666;
 wire net5667;
 wire net5668;
 wire net5669;
 wire net5670;
 wire net5671;
 wire net5672;
 wire net5673;
 wire net5674;
 wire net5675;
 wire net5676;
 wire net5677;
 wire net5678;
 wire net5679;
 wire net5680;
 wire net5681;
 wire net5682;
 wire net5683;
 wire net5684;
 wire net5685;
 wire net5686;
 wire net5687;
 wire net5688;
 wire net5689;
 wire net5690;
 wire net5691;
 wire net5692;
 wire net5693;
 wire net5694;
 wire net5695;
 wire net5696;
 wire net5697;
 wire net5698;
 wire net5699;
 wire net5700;
 wire net5701;
 wire net5702;
 wire net5703;
 wire net5704;
 wire net5705;
 wire net5706;
 wire net5707;
 wire net5708;
 wire net5709;
 wire net5710;
 wire net5711;
 wire net5712;
 wire net5713;
 wire net5714;
 wire net5715;
 wire net5716;
 wire net5717;
 wire net5718;
 wire net5719;
 wire net5720;
 wire net5721;
 wire net5722;
 wire net5723;
 wire net5724;
 wire net5725;
 wire net5726;
 wire net5727;
 wire net5728;
 wire net5729;
 wire net5730;
 wire net5731;
 wire net5732;
 wire net5733;
 wire net5734;
 wire net5735;
 wire net5736;
 wire net5737;
 wire net5738;
 wire net5739;
 wire net5740;
 wire net5741;
 wire net5742;
 wire net5743;
 wire net5744;
 wire net5745;
 wire net5746;
 wire net5747;
 wire net5748;
 wire net5749;
 wire net5750;
 wire net5751;
 wire net5752;
 wire net5753;
 wire net5754;
 wire net5755;
 wire net5756;
 wire net5757;
 wire net5758;
 wire net5759;
 wire net5760;
 wire net5761;
 wire net5762;
 wire net5763;
 wire net5764;
 wire net5765;
 wire net5766;
 wire net5767;
 wire net5768;
 wire net5769;
 wire net5770;
 wire net5771;
 wire net5772;
 wire net5773;
 wire net5774;
 wire net5775;
 wire net5776;
 wire net5777;
 wire net5778;
 wire net5779;
 wire net5780;
 wire net5781;
 wire net5782;
 wire net5783;
 wire net5784;
 wire net5785;
 wire net5786;
 wire net5787;
 wire net5788;
 wire net5789;
 wire net5790;
 wire net5791;
 wire net5792;
 wire net5793;
 wire net5794;
 wire net5795;
 wire net5796;
 wire net5797;
 wire net5798;
 wire net5799;
 wire net5800;
 wire net5801;
 wire net5802;
 wire net5803;
 wire net5804;
 wire net5805;
 wire net5806;
 wire net5807;
 wire net5808;
 wire net5809;
 wire net5810;
 wire net5811;
 wire net5812;
 wire net5813;
 wire net5814;
 wire net5815;
 wire net5816;
 wire net5817;
 wire net5818;
 wire net5819;
 wire net5820;
 wire net5821;
 wire net5822;
 wire net5823;
 wire net5824;
 wire net5825;
 wire net5826;
 wire net5827;
 wire net5828;
 wire net5829;
 wire net5830;
 wire net5831;
 wire net5832;
 wire net5833;
 wire net5834;
 wire net5835;
 wire net5836;
 wire net5837;
 wire net5838;
 wire net5839;
 wire net5840;
 wire net5841;
 wire net5842;
 wire net5843;
 wire net5844;
 wire net5845;
 wire net5846;
 wire net5847;
 wire net5848;
 wire net5849;
 wire net5850;
 wire net5851;
 wire net5852;
 wire net5853;
 wire net5854;
 wire net5855;
 wire net5856;
 wire net5857;
 wire net5858;
 wire net5859;
 wire net5860;
 wire net5861;
 wire net5862;
 wire net5863;
 wire net5864;
 wire net5865;
 wire net5866;
 wire net5867;
 wire net5868;
 wire net5869;
 wire net5870;
 wire net5871;
 wire net5872;
 wire net5873;
 wire net5874;
 wire net5875;
 wire net5876;
 wire net5877;
 wire net5878;
 wire net5879;
 wire net5880;
 wire net5881;
 wire net5882;
 wire net5883;
 wire net5884;
 wire net5885;
 wire net5886;
 wire net5887;
 wire net5888;
 wire net5889;
 wire net5890;
 wire net5891;
 wire net5892;
 wire net5893;
 wire net5894;
 wire net5895;
 wire net5896;
 wire net5897;
 wire net5898;
 wire net5899;
 wire net5900;
 wire net5901;
 wire net5902;
 wire net5903;
 wire net5904;
 wire net5905;
 wire net5906;
 wire net5907;
 wire net5908;
 wire net5909;
 wire net5910;
 wire net5911;
 wire net5912;
 wire net5913;
 wire net5914;
 wire net5915;
 wire net5916;
 wire net5917;
 wire net5918;
 wire net5919;
 wire net5920;
 wire net5921;
 wire net5922;
 wire net5923;
 wire net5924;
 wire net5925;
 wire net5926;
 wire net5927;
 wire net5928;
 wire net5929;
 wire net5930;
 wire net5931;
 wire net5932;
 wire net5933;
 wire net5934;
 wire net5935;
 wire net5936;
 wire net5937;
 wire net5938;
 wire net5939;
 wire net5940;
 wire net5941;
 wire net5942;
 wire net5943;
 wire net5944;
 wire net5945;
 wire net5946;
 wire net5947;
 wire net5948;
 wire net5949;
 wire net5950;
 wire net5951;
 wire net5952;
 wire net5953;
 wire net5954;
 wire net5955;
 wire net5956;
 wire net5957;
 wire net5958;
 wire net5959;
 wire net5960;
 wire net5961;
 wire net5962;
 wire net5963;
 wire net5964;
 wire net5965;
 wire net5966;
 wire net5967;
 wire net5968;
 wire net5969;
 wire net5970;
 wire net5971;
 wire net5972;
 wire net5973;
 wire net5974;
 wire net5975;
 wire net5976;
 wire net5977;
 wire net5978;
 wire net5979;
 wire net5980;
 wire net5981;
 wire net5982;
 wire net5983;
 wire net5984;
 wire net5985;
 wire net5986;
 wire net5987;
 wire net5988;
 wire net5989;
 wire net5990;
 wire net5991;
 wire net5992;
 wire net5993;
 wire net5994;
 wire net5995;
 wire net5996;
 wire net5997;
 wire net5998;
 wire net5999;
 wire net6000;
 wire net6001;
 wire net6002;
 wire net6003;
 wire net6004;
 wire net6005;
 wire net6006;
 wire net6007;
 wire net6008;
 wire net6009;
 wire net6010;
 wire net6011;
 wire net6012;
 wire net6013;
 wire net6014;
 wire net6015;
 wire net6016;
 wire net6017;
 wire net6018;
 wire net6019;
 wire net6020;
 wire net6021;
 wire net6022;
 wire net6023;
 wire net6024;
 wire net6025;
 wire net6026;
 wire net6027;
 wire net6028;
 wire net6029;
 wire net6030;
 wire net6031;
 wire net6032;
 wire net6033;
 wire net6034;
 wire net6035;
 wire net6036;
 wire net6037;
 wire net6038;
 wire net6039;
 wire net6040;
 wire net6041;
 wire net6042;
 wire net6043;
 wire net6044;
 wire net6045;
 wire net6046;
 wire net6047;
 wire net6048;
 wire net6049;
 wire net6050;
 wire net6051;
 wire net6052;
 wire net6053;
 wire net6054;
 wire net6055;
 wire net6056;
 wire net6057;
 wire net6058;
 wire net6059;
 wire net6060;
 wire net6061;
 wire net6062;
 wire net6063;
 wire net6064;
 wire net6065;
 wire net6066;
 wire net6067;
 wire net6068;
 wire net6069;
 wire net6070;
 wire net6071;
 wire net6072;
 wire net6073;
 wire net6074;
 wire net6075;
 wire net6076;
 wire net6077;
 wire net6078;
 wire net6079;
 wire net6080;
 wire net6081;
 wire net6082;
 wire net6083;
 wire net6084;
 wire net6085;
 wire net6086;
 wire net6087;
 wire net6088;
 wire net6089;
 wire net6090;
 wire net6091;
 wire net6092;
 wire net6093;
 wire net6094;
 wire net6095;
 wire net6096;
 wire net6097;
 wire net6098;
 wire net6099;
 wire net6100;
 wire net6101;
 wire net6102;
 wire net6103;
 wire net6104;
 wire net6105;
 wire net6106;
 wire net6107;
 wire net6108;
 wire net6109;
 wire net6110;
 wire net6111;
 wire net6112;
 wire net6113;
 wire net6114;
 wire net6115;
 wire net6116;
 wire net6117;
 wire net6118;
 wire net6119;
 wire net6120;
 wire net6121;
 wire net6122;
 wire net6123;
 wire net6124;
 wire net6125;
 wire net6126;
 wire net6127;
 wire net6128;
 wire net6129;
 wire net6130;
 wire net6131;
 wire net6132;
 wire net6133;
 wire net6134;
 wire net6135;
 wire net6136;
 wire net6137;
 wire net6138;
 wire net6139;
 wire net6140;
 wire net6141;
 wire net6142;
 wire net6143;
 wire net6144;
 wire net6145;
 wire net6146;
 wire net6147;
 wire net6148;
 wire net6149;
 wire net6150;
 wire net6151;
 wire net6152;
 wire net6153;
 wire net6154;
 wire net6155;
 wire net6156;
 wire net6157;
 wire net6158;
 wire net6159;
 wire net6160;
 wire net6161;
 wire net6162;
 wire net6163;
 wire net6164;
 wire net6165;
 wire net6166;
 wire net6167;
 wire net6168;
 wire net6169;
 wire net6170;
 wire net6171;
 wire net6172;
 wire net6173;
 wire net6174;
 wire net6175;
 wire net6176;
 wire net6177;
 wire net6178;
 wire net6179;
 wire net6180;
 wire net6181;
 wire net6182;
 wire net6183;
 wire net6184;
 wire net6185;
 wire net6186;
 wire net6187;
 wire net6188;
 wire net6189;
 wire net6190;
 wire net6191;
 wire net6192;
 wire net6193;
 wire net6194;
 wire net6195;
 wire net6196;
 wire net6197;
 wire net6198;
 wire net6199;
 wire net6200;
 wire net6201;
 wire net6202;
 wire net6203;
 wire net6204;
 wire net6205;
 wire net6206;
 wire net6207;
 wire net6208;
 wire net6209;
 wire net6210;
 wire net6211;
 wire net6212;
 wire net6213;
 wire net6214;
 wire net6215;
 wire net6216;
 wire net6217;
 wire net6218;
 wire net6219;
 wire net6220;
 wire net6221;
 wire net6222;
 wire net6223;
 wire net6224;
 wire net6225;
 wire net6226;
 wire net6227;
 wire net6228;
 wire net6229;
 wire net6230;
 wire net6231;
 wire net6232;
 wire net6233;
 wire net6234;
 wire net6235;
 wire net6236;
 wire net6237;
 wire net6238;
 wire net6239;
 wire net6240;
 wire net6241;
 wire net6242;
 wire net6243;
 wire net6244;
 wire net6245;
 wire net6246;
 wire net6247;
 wire net6248;
 wire net6249;
 wire net6250;
 wire net6251;
 wire net6252;
 wire net6253;
 wire net6254;
 wire net6255;
 wire net6256;
 wire net6257;
 wire net6258;
 wire net6259;
 wire net6260;
 wire net6261;
 wire net6262;
 wire net6263;
 wire net6264;
 wire net6265;
 wire net6266;
 wire net6267;
 wire net6268;
 wire net6269;
 wire net6270;
 wire net6271;
 wire net6272;
 wire net6273;
 wire net6274;
 wire net6275;
 wire net6276;
 wire net6277;
 wire net6278;
 wire net6279;
 wire net6280;
 wire net6281;
 wire net6282;
 wire net6283;
 wire net6284;
 wire net6285;
 wire net6286;
 wire net6287;
 wire net6288;
 wire net6289;
 wire net6290;
 wire net6291;
 wire net6292;
 wire net6293;
 wire net6294;
 wire net6295;
 wire net6296;
 wire net6297;
 wire net6298;
 wire net6299;
 wire net6300;
 wire net6301;
 wire net6302;
 wire net6303;
 wire net6304;
 wire net6305;
 wire net6306;
 wire net6307;
 wire net6308;
 wire net6309;
 wire net6310;
 wire net6311;
 wire net6312;
 wire net6313;
 wire net6314;
 wire net6315;
 wire net6316;
 wire net6317;
 wire net6318;
 wire net6319;
 wire net6320;
 wire net6321;
 wire net6322;
 wire net6323;
 wire net6324;
 wire net6325;
 wire net6326;
 wire net6327;
 wire net6328;
 wire net6329;
 wire net6330;
 wire net6331;
 wire net6332;
 wire net6333;
 wire net6334;
 wire net6335;
 wire net6336;
 wire net6337;
 wire net6338;
 wire net6339;
 wire net6340;
 wire net6341;
 wire net6342;
 wire net6343;
 wire net6344;
 wire net6345;
 wire net6346;
 wire net6347;
 wire net6348;
 wire net6349;
 wire net6350;
 wire net6351;
 wire net6352;
 wire net6353;
 wire net6354;
 wire net6355;
 wire net6356;
 wire net6357;
 wire net6358;
 wire net6359;
 wire net6360;
 wire net6361;
 wire net6362;
 wire net6363;
 wire net6364;
 wire net6365;
 wire net6366;
 wire net6367;
 wire net6368;
 wire net6369;
 wire net6370;
 wire net6371;
 wire net6372;
 wire net6373;
 wire net6374;
 wire net6375;
 wire net6376;
 wire net6377;
 wire net6378;
 wire net6379;
 wire net6380;
 wire net6381;
 wire net6382;
 wire net6383;
 wire net6384;
 wire net6385;
 wire net6386;
 wire net6387;
 wire net6388;
 wire net6389;
 wire net6390;
 wire net6391;
 wire net6392;
 wire net6393;
 wire net6394;
 wire net6395;
 wire net6396;
 wire net6397;
 wire net6398;
 wire net6399;
 wire net6400;
 wire net6401;
 wire net6402;
 wire net6403;
 wire net6404;
 wire net6405;
 wire net6406;
 wire net6407;
 wire net6408;
 wire net6409;
 wire net6410;
 wire net6411;
 wire net6412;
 wire net6413;
 wire net6414;
 wire net6415;
 wire net6416;
 wire net6417;
 wire net6418;
 wire net6419;
 wire net6420;
 wire net6421;
 wire net6422;
 wire net6423;
 wire net6424;
 wire net6425;
 wire net6426;
 wire net6427;
 wire net6428;
 wire net6429;
 wire net6430;
 wire net6431;
 wire net6432;
 wire net6433;
 wire net6434;
 wire net6435;
 wire net6436;
 wire net6437;
 wire net6438;
 wire net6439;
 wire net6440;
 wire net6441;
 wire net6442;
 wire net6443;
 wire net6444;
 wire net6445;
 wire net6446;
 wire net6447;
 wire net6448;
 wire net6449;
 wire net6450;
 wire net6451;
 wire net6452;
 wire net6453;
 wire net6454;
 wire net6455;
 wire net6456;
 wire net6457;
 wire net6458;
 wire net6459;
 wire net6460;
 wire net6461;
 wire net6462;
 wire net6463;
 wire net6464;
 wire net6465;
 wire net6466;
 wire net6467;
 wire net6468;
 wire net6469;
 wire net6470;
 wire net6471;
 wire net6472;
 wire net6473;
 wire net6474;
 wire net6475;
 wire net6476;
 wire net6477;
 wire net6478;
 wire net6479;
 wire net6480;
 wire net6481;
 wire net6482;
 wire net6483;
 wire net6484;
 wire net6485;
 wire net6486;
 wire net6487;
 wire net6488;
 wire net6489;
 wire net6490;
 wire net6491;
 wire net6492;
 wire net6493;
 wire net6494;
 wire net6495;
 wire net6496;
 wire net6497;
 wire net6498;
 wire net6499;
 wire net6500;
 wire net6501;
 wire net6502;
 wire net6503;
 wire net6504;
 wire net6505;
 wire net6506;
 wire net6507;
 wire net6508;
 wire net6509;
 wire net6510;
 wire net6511;
 wire net6512;
 wire net6513;
 wire net6514;
 wire net6515;
 wire net6516;
 wire net6517;
 wire net6518;
 wire net6519;
 wire net6520;
 wire net6521;
 wire net6522;
 wire net6523;
 wire net6524;
 wire net6525;
 wire net6526;
 wire net6527;
 wire net6528;
 wire net6529;
 wire net6530;
 wire net6531;
 wire net6532;
 wire net6533;
 wire net6534;
 wire net6535;
 wire net6536;
 wire net6537;
 wire net6538;
 wire net6539;
 wire net6540;
 wire net6541;
 wire net6542;
 wire net6543;
 wire net6544;
 wire net6545;
 wire net6546;
 wire net6547;
 wire net6548;
 wire net6549;
 wire net6550;
 wire net6551;
 wire net6552;
 wire net6553;
 wire net6554;
 wire net6555;
 wire net6556;
 wire net6557;
 wire net6558;
 wire net6559;
 wire net6560;
 wire net6561;
 wire net6562;
 wire net6563;
 wire net6564;
 wire net6565;
 wire net6566;
 wire net6567;
 wire net6568;
 wire net6569;
 wire net6570;
 wire net6571;
 wire net6572;
 wire net6573;
 wire net6574;
 wire net6575;
 wire net6576;
 wire net6577;
 wire net6578;
 wire net6579;
 wire net6580;
 wire net6581;
 wire net6582;
 wire net6583;
 wire net6584;
 wire net6585;
 wire net6586;
 wire net6587;
 wire net6588;
 wire net6589;
 wire net6590;
 wire net6591;
 wire net6592;
 wire net6593;
 wire net6594;
 wire net6595;
 wire net6596;
 wire net6597;
 wire net6598;
 wire net6599;
 wire net6600;
 wire net6601;
 wire net6602;
 wire net6603;
 wire net6604;
 wire net6605;
 wire net6606;
 wire net6607;
 wire net6608;
 wire net6609;
 wire net6610;
 wire net6611;
 wire net6612;
 wire net6613;
 wire net6614;
 wire net6615;
 wire net6616;
 wire net6617;
 wire net6618;
 wire net6619;
 wire net6620;
 wire net6621;
 wire net6622;
 wire net6623;
 wire net6624;
 wire net6625;
 wire net6626;
 wire net6627;
 wire net6628;
 wire net6629;
 wire net6630;
 wire net6631;
 wire net6632;
 wire net6633;
 wire net6634;
 wire net6635;
 wire net6636;
 wire net6637;
 wire net6638;
 wire net6639;
 wire net6640;
 wire net6641;
 wire net6642;
 wire net6643;
 wire net6644;
 wire net6645;
 wire net6646;
 wire net6647;
 wire net6648;
 wire net6649;
 wire net6650;
 wire net6651;
 wire net6652;
 wire net6653;
 wire net6654;
 wire net6655;
 wire net6656;
 wire net6657;
 wire net6658;
 wire net6659;
 wire net6660;
 wire net6661;
 wire net6662;
 wire net6663;
 wire net6664;
 wire net6665;
 wire net6666;
 wire net6667;
 wire net6668;
 wire net6669;
 wire net6670;
 wire net6671;
 wire net6672;
 wire net6673;
 wire net6674;
 wire net6675;
 wire net6676;
 wire net6677;
 wire net6678;
 wire net6679;
 wire net6680;
 wire net6681;
 wire net6682;
 wire net6683;
 wire net6684;
 wire net6685;
 wire net6686;
 wire net6687;
 wire net6688;
 wire net6689;
 wire net6690;
 wire net6691;
 wire net6692;
 wire net6693;
 wire net6694;
 wire net6695;
 wire net6696;
 wire net6697;
 wire net6698;
 wire net6699;
 wire net6700;
 wire net6701;
 wire net6702;
 wire net6703;
 wire net6704;
 wire net6705;
 wire net6706;
 wire net6707;
 wire net6708;
 wire net6709;
 wire net6710;
 wire net6711;
 wire net6712;
 wire net6713;
 wire net6714;
 wire net6715;
 wire net6716;
 wire net6717;
 wire net6718;
 wire net6719;
 wire net6720;
 wire net6721;
 wire net6722;
 wire net6723;
 wire net6724;
 wire net6725;
 wire net6726;
 wire net6727;
 wire net6728;
 wire net6729;
 wire net6730;
 wire net6731;
 wire net6732;
 wire net6733;
 wire net6734;
 wire net6735;
 wire net6736;
 wire net6737;
 wire net6738;
 wire net6739;
 wire net6740;
 wire net6741;
 wire net6742;
 wire net6743;
 wire net6744;
 wire net6745;
 wire net6746;
 wire net6747;
 wire net6748;
 wire net6749;
 wire net6750;
 wire net6751;
 wire net6752;
 wire net6753;
 wire net6754;
 wire net6755;
 wire net6756;
 wire net6757;
 wire net6758;
 wire net6759;
 wire net6760;
 wire net6761;
 wire net6762;
 wire net6763;
 wire net6764;
 wire net6765;
 wire net6766;
 wire net6767;
 wire net6768;
 wire net6769;
 wire net6770;
 wire net6771;
 wire net6772;
 wire net6773;
 wire net6774;
 wire net6775;
 wire net6776;
 wire net6777;
 wire net6778;
 wire net6779;
 wire net6780;
 wire net6781;
 wire net6782;
 wire net6783;
 wire net6784;
 wire net6785;
 wire net6786;
 wire net6787;
 wire net6788;
 wire net6789;
 wire net6790;
 wire net6791;
 wire net6792;
 wire net6793;
 wire net6794;
 wire net6795;
 wire net6796;
 wire net6797;
 wire net6798;
 wire net6799;
 wire net6800;
 wire net6801;
 wire net6802;
 wire net6803;
 wire net6804;
 wire net6805;
 wire net6806;
 wire net6807;
 wire net6808;
 wire net6809;
 wire net6810;
 wire net6811;
 wire net6812;
 wire net6813;
 wire net6814;
 wire net6815;
 wire net6816;
 wire net6817;
 wire net6818;
 wire net6819;
 wire net6820;
 wire net6821;
 wire net6822;
 wire net6823;
 wire net6824;
 wire net6825;
 wire net6826;
 wire net6827;
 wire net6828;
 wire net6829;
 wire net6830;
 wire net6831;
 wire net6832;
 wire net6833;
 wire net6834;
 wire net6835;
 wire net6836;
 wire net6837;
 wire net6838;
 wire net6839;
 wire net6840;
 wire net6841;
 wire net6842;
 wire net6843;
 wire net6844;
 wire net6845;
 wire net6846;
 wire net6847;
 wire net6848;
 wire net6849;
 wire net6850;
 wire net6851;
 wire net6852;
 wire net6853;
 wire net6854;
 wire net6855;
 wire net6856;
 wire net6857;
 wire net6858;
 wire net6859;
 wire net6860;
 wire net6861;
 wire net6862;
 wire net6863;
 wire net6864;
 wire net6865;
 wire net6866;
 wire net6867;
 wire net6868;
 wire net6869;
 wire net6870;
 wire net6871;
 wire net6872;
 wire net6873;
 wire net6874;
 wire net6875;
 wire net6876;
 wire net6877;
 wire net6878;
 wire net6879;
 wire net6880;
 wire net6881;
 wire net6882;
 wire net6883;
 wire net6884;
 wire net6885;
 wire net6886;
 wire net6887;
 wire net6888;
 wire net6889;
 wire net6890;
 wire net6891;
 wire net6892;
 wire net6893;
 wire net6894;
 wire net6895;
 wire net6896;
 wire net6897;
 wire net6898;
 wire net6899;
 wire net6900;
 wire net6901;
 wire net6902;
 wire net6903;
 wire net6904;
 wire net6905;
 wire net6906;
 wire net6907;
 wire net6908;
 wire net6909;
 wire net6910;
 wire net6911;
 wire net6912;
 wire net6913;
 wire net6914;
 wire net6915;
 wire net6916;
 wire net6917;
 wire net6918;
 wire net6919;
 wire net6920;
 wire net6921;
 wire net6922;
 wire net6923;
 wire net6924;
 wire net6925;
 wire net6926;
 wire net6927;
 wire net6928;
 wire net6929;
 wire net6930;
 wire net6931;
 wire net6932;
 wire net6933;
 wire net6934;
 wire net6935;
 wire net6936;
 wire net6937;
 wire net6938;
 wire net6939;
 wire net6940;
 wire net6941;
 wire net6942;
 wire net6943;
 wire net6944;
 wire net6945;
 wire net6946;
 wire net6947;
 wire net6948;
 wire net6949;
 wire net6950;
 wire net6951;
 wire net6952;
 wire net6953;
 wire net6954;
 wire net6955;
 wire net6956;
 wire net6957;
 wire net6958;
 wire net6959;
 wire net6960;
 wire net6961;
 wire net6962;
 wire net6963;
 wire net6964;
 wire net6965;
 wire net6966;
 wire net6967;
 wire net6968;
 wire net6969;
 wire net6970;
 wire net6971;
 wire net6972;
 wire net6973;
 wire net6974;
 wire net6975;
 wire net6976;
 wire net6977;
 wire net6978;
 wire net6979;
 wire net6980;
 wire net6981;
 wire net6982;
 wire net6983;
 wire net6984;
 wire net6985;
 wire net6986;
 wire net6987;
 wire net6988;
 wire net6989;
 wire net6990;
 wire net6991;
 wire net6992;
 wire net6993;
 wire net6994;
 wire net6995;
 wire net6996;
 wire net6997;
 wire net6998;
 wire net6999;
 wire net7000;
 wire net7001;
 wire net7002;
 wire net7003;
 wire net7004;
 wire net7005;
 wire net7006;
 wire net7007;
 wire net7008;
 wire net7009;
 wire net7010;
 wire net7011;
 wire net7012;
 wire net7013;
 wire net7014;
 wire net7015;
 wire net7016;
 wire net7017;
 wire net7018;
 wire net7019;
 wire net7020;
 wire net7021;
 wire net7022;
 wire net7023;
 wire net7024;
 wire net7025;
 wire net7026;
 wire net7027;
 wire net7028;
 wire net7029;
 wire net7030;
 wire net7031;
 wire net7032;
 wire net7033;
 wire net7034;
 wire net7035;
 wire net7036;
 wire net7037;
 wire net7038;
 wire net7039;
 wire net7040;
 wire net7041;
 wire net7042;
 wire net7043;
 wire net7044;
 wire net7045;
 wire net7046;
 wire net7047;
 wire net7048;
 wire net7049;
 wire net7050;
 wire net7051;
 wire net7052;
 wire net7053;
 wire net7054;
 wire net7055;
 wire net7056;
 wire net7057;
 wire net7058;
 wire net7059;
 wire net7060;
 wire net7061;
 wire net7062;
 wire net7063;
 wire net7064;
 wire net7065;
 wire net7066;
 wire net7067;
 wire net7068;
 wire net7069;
 wire net7070;
 wire net7071;
 wire net7072;
 wire net7073;
 wire net7074;
 wire net7075;
 wire net7076;
 wire net7077;
 wire net7078;
 wire net7079;
 wire net7080;
 wire net7081;
 wire net7082;
 wire net7083;
 wire net7084;
 wire net7085;
 wire net7086;
 wire net7087;
 wire net7088;
 wire net7089;
 wire net7090;
 wire net7091;
 wire net7092;
 wire net7093;
 wire net7094;
 wire net7095;
 wire net7096;
 wire net7097;
 wire net7098;
 wire net7099;
 wire net7100;
 wire net7101;
 wire net7102;
 wire net7103;
 wire net7104;
 wire net7105;
 wire net7106;
 wire net7107;
 wire net7108;
 wire net7109;
 wire net7110;
 wire net7111;
 wire net7112;
 wire net7113;
 wire net7114;
 wire net7115;
 wire net7116;
 wire net7117;
 wire net7118;
 wire net7119;
 wire net7120;
 wire net7121;
 wire net7122;
 wire net7123;
 wire net7124;
 wire net7125;
 wire net7126;
 wire net7127;
 wire net7128;
 wire net7129;
 wire net7130;
 wire net7131;
 wire net7132;
 wire net7133;
 wire net7134;
 wire net7135;
 wire net7136;
 wire net7137;
 wire net7138;
 wire net7139;
 wire net7140;
 wire net7141;
 wire net7142;
 wire net7143;
 wire net7144;
 wire net7145;
 wire net7146;
 wire net7147;
 wire net7148;
 wire net7149;
 wire net7150;
 wire net7151;
 wire net7152;
 wire net7153;
 wire net7154;
 wire net7155;
 wire net7156;
 wire net7157;
 wire net7158;
 wire net7159;
 wire net7160;
 wire net7161;
 wire net7162;
 wire net7163;
 wire net7164;
 wire net7165;
 wire net7166;
 wire net7167;
 wire net7168;
 wire net7169;
 wire net7170;
 wire net7171;
 wire net7172;
 wire net7173;
 wire net7174;
 wire net7175;
 wire net7176;
 wire net7177;
 wire net7178;
 wire net7179;
 wire net7180;
 wire net7181;
 wire net7182;
 wire net7183;
 wire net7184;
 wire net7185;
 wire net7186;
 wire net7187;
 wire net7188;
 wire net7189;
 wire net7190;
 wire net7191;
 wire net7192;
 wire net7193;
 wire net7194;
 wire net7195;
 wire net7196;
 wire net7197;
 wire net7198;
 wire net7199;
 wire net7200;
 wire net7201;
 wire net7202;
 wire net7203;
 wire net7204;
 wire net7205;
 wire net7206;
 wire net7207;
 wire net7208;
 wire net7209;
 wire net7210;
 wire net7211;
 wire net7212;
 wire net7213;
 wire net7214;
 wire net7215;
 wire net7216;
 wire net7217;
 wire net7218;
 wire net7219;
 wire net7220;
 wire net7221;
 wire net7222;
 wire net7223;
 wire net7224;
 wire net7225;
 wire net7226;
 wire net7227;
 wire net7228;
 wire net7229;
 wire net7230;
 wire net7231;
 wire net7232;
 wire net7233;
 wire net7234;
 wire net7235;
 wire net7236;
 wire net7237;
 wire net7238;
 wire net7239;
 wire net7240;
 wire net7241;
 wire net7242;
 wire net7243;
 wire net7244;
 wire net7245;
 wire net7246;
 wire net7247;
 wire net7248;
 wire net7249;
 wire net7250;
 wire net7251;
 wire net7252;
 wire net7253;
 wire net7254;
 wire net7255;
 wire net7256;
 wire net7257;
 wire net7258;
 wire net7259;
 wire net7260;
 wire net7261;
 wire net7262;
 wire net7263;
 wire net7264;
 wire net7265;
 wire net7266;
 wire net7267;
 wire net7268;
 wire net7269;
 wire net7270;
 wire net7271;
 wire net7272;
 wire net7273;
 wire net7274;
 wire net7275;
 wire net7276;
 wire net7277;
 wire net7278;
 wire net7279;
 wire net7280;
 wire net7281;
 wire net7282;
 wire net7283;
 wire net7284;
 wire net7285;
 wire net7286;
 wire net7287;
 wire net7288;
 wire net7289;
 wire net7290;
 wire net7291;
 wire net7292;
 wire net7293;
 wire net7294;
 wire net7295;
 wire net7296;
 wire net7297;
 wire net7298;
 wire net7299;
 wire net7300;
 wire net7301;
 wire net7302;
 wire net7303;
 wire net7304;
 wire net7305;
 wire net7306;
 wire net7307;
 wire net7308;
 wire net7309;
 wire net7310;
 wire net7311;
 wire net7312;
 wire net7313;
 wire net7314;
 wire net7315;
 wire net7316;
 wire net7317;
 wire net7318;
 wire net7319;
 wire net7320;
 wire net7321;
 wire net7322;
 wire net7323;
 wire net7324;
 wire net7325;
 wire net7326;
 wire net7327;
 wire net7328;
 wire net7329;
 wire net7330;
 wire net7331;
 wire net7332;
 wire net7333;
 wire net7334;
 wire net7335;
 wire net7336;
 wire net7337;
 wire net7338;
 wire net7339;
 wire net7340;
 wire net7341;
 wire net7342;
 wire net7343;
 wire net7344;
 wire net7345;
 wire net7346;
 wire net7347;
 wire net7348;
 wire net7349;
 wire net7350;
 wire net7351;
 wire net7352;
 wire net7353;
 wire net7354;
 wire net7355;
 wire net7356;
 wire net7357;
 wire net7358;
 wire net7359;
 wire net7360;
 wire net7361;
 wire net7362;
 wire net7363;
 wire net7364;
 wire net7365;
 wire net7366;
 wire net7367;
 wire net7368;
 wire net7369;
 wire net7370;
 wire net7371;
 wire net7372;
 wire net7373;
 wire net7374;
 wire net7375;
 wire net7376;
 wire net7377;
 wire net7378;
 wire net7379;
 wire net7380;
 wire net7381;
 wire net7382;
 wire net7383;
 wire net7384;
 wire net7385;
 wire net7386;
 wire net7387;
 wire net7388;
 wire net7389;
 wire net7390;
 wire net7391;
 wire net7392;
 wire net7393;
 wire net7394;
 wire net7395;
 wire net7396;
 wire net7397;
 wire net7398;
 wire net7399;
 wire net7400;
 wire net7401;
 wire net7402;
 wire net7403;
 wire net7404;
 wire net7405;
 wire net7406;
 wire net7407;
 wire net7408;
 wire net7409;
 wire net7410;
 wire net7411;
 wire net7412;
 wire net7413;
 wire net7414;
 wire net7415;
 wire net7416;
 wire net7417;
 wire net7418;
 wire net7419;
 wire net7420;
 wire net7421;
 wire net7422;
 wire net7423;
 wire net7424;
 wire net7425;
 wire net7426;
 wire net7427;
 wire net7428;
 wire net7429;
 wire net7430;
 wire net7431;
 wire net7432;
 wire net7433;
 wire net7434;
 wire net7435;
 wire net7436;
 wire net7437;
 wire net7438;
 wire net7439;
 wire net7440;
 wire net7441;
 wire net7442;
 wire net7443;
 wire net7444;
 wire net7445;
 wire net7446;
 wire net7447;
 wire net7448;
 wire net7449;
 wire net7450;
 wire net7451;
 wire net7452;
 wire net7453;
 wire net7454;
 wire net7455;
 wire net7456;
 wire net7457;
 wire net7458;
 wire net7459;
 wire net7460;
 wire net7461;
 wire net7462;
 wire net7463;
 wire net7464;
 wire net7465;
 wire net7466;
 wire net7467;
 wire net7468;
 wire net7469;
 wire net7470;
 wire net7471;
 wire net7472;
 wire net7473;
 wire net7474;
 wire net7475;
 wire net7476;
 wire net7477;
 wire net7478;
 wire net7479;
 wire net7480;
 wire net7481;
 wire net7482;
 wire net7483;
 wire net7484;
 wire net7485;
 wire net7486;
 wire net7487;
 wire net7488;
 wire net7489;
 wire net7490;
 wire net7491;
 wire net7492;
 wire net7493;
 wire net7494;
 wire net7495;
 wire net7496;
 wire net7497;
 wire net7498;
 wire net7499;
 wire net7500;
 wire net7501;
 wire net7502;
 wire net7503;
 wire net7504;
 wire net7505;
 wire net7506;
 wire net7507;
 wire net7508;
 wire net7509;
 wire net7510;
 wire net7511;
 wire net7512;
 wire net7513;
 wire net7514;
 wire net7515;
 wire net7516;
 wire net7517;
 wire net7518;
 wire net7519;
 wire net7520;
 wire net7521;
 wire net7522;
 wire net7523;
 wire net7524;
 wire net7525;
 wire net7526;
 wire net7527;
 wire net7528;
 wire net7529;
 wire net7530;
 wire net7531;
 wire net7532;
 wire net7533;
 wire net7534;
 wire net7535;
 wire net7536;
 wire net7537;
 wire net7538;
 wire net7539;
 wire net7540;
 wire net7541;
 wire net7542;
 wire net7543;
 wire net7544;
 wire net7545;
 wire net7546;
 wire net7547;
 wire net7548;
 wire net7549;
 wire net7550;
 wire net7551;
 wire net7552;
 wire net7553;
 wire net7554;
 wire net7555;
 wire net7556;
 wire net7557;
 wire net7558;
 wire net7559;
 wire net7560;
 wire net7561;
 wire net7562;
 wire net7563;
 wire net7564;
 wire net7565;
 wire net7566;
 wire net7567;
 wire net7568;
 wire net7569;
 wire net7570;
 wire net7571;
 wire net7572;
 wire net7573;
 wire net7574;
 wire net7575;
 wire net7576;
 wire net7577;
 wire net7578;
 wire net7579;
 wire net7580;
 wire net7581;
 wire net7582;
 wire net7583;
 wire net7584;
 wire net7585;
 wire net7586;
 wire net7587;
 wire net7588;
 wire net7589;
 wire net7590;
 wire net7591;
 wire net7592;
 wire net7593;
 wire net7594;
 wire net7595;
 wire net7596;
 wire net7597;
 wire net7598;
 wire net7599;
 wire net7600;
 wire net7601;
 wire net7602;
 wire net7603;
 wire net7604;
 wire net7605;
 wire net7606;
 wire net7607;
 wire net7608;
 wire net7609;
 wire net7610;
 wire net7611;
 wire net7612;
 wire net7613;
 wire net7614;
 wire net7615;
 wire net7616;
 wire net7617;
 wire net7618;
 wire net7619;
 wire net7620;
 wire net7621;
 wire net7622;
 wire net7623;
 wire net7624;
 wire net7625;
 wire net7626;
 wire net7627;
 wire net7628;
 wire net7629;
 wire net7630;
 wire net7631;
 wire net7632;
 wire net7633;
 wire net7634;
 wire net7635;
 wire net7636;
 wire net7637;
 wire net7638;
 wire net7639;
 wire net7640;
 wire net7641;
 wire net7642;
 wire net7643;
 wire net7644;
 wire net7645;
 wire net7646;
 wire net7647;
 wire net7648;
 wire net7649;
 wire net7650;
 wire net7651;
 wire net7652;
 wire net7653;
 wire net7654;
 wire net7655;
 wire net7656;
 wire net7657;
 wire net7658;
 wire net7659;
 wire net7660;
 wire net7661;
 wire net7662;
 wire net7663;
 wire net7664;
 wire net7665;
 wire net7666;
 wire net7667;
 wire net7668;
 wire net7669;
 wire net7670;
 wire net7671;
 wire net7672;
 wire net7673;
 wire net7674;
 wire net7675;
 wire net7676;
 wire net7677;
 wire net7678;
 wire net7679;
 wire net7680;
 wire net7681;
 wire net7682;
 wire net7683;
 wire net7684;
 wire net7685;
 wire net7686;
 wire net7687;
 wire net7688;
 wire net7689;
 wire net7690;
 wire net7691;
 wire net7692;
 wire net7693;
 wire net7694;
 wire net7695;
 wire net7696;
 wire net7697;
 wire net7698;
 wire net7699;
 wire net7700;
 wire net7701;
 wire net7702;
 wire net7703;
 wire net7704;
 wire net7705;
 wire net7706;
 wire net7707;
 wire net7708;
 wire net7709;
 wire net7710;
 wire net7711;
 wire net7712;
 wire net7713;
 wire net7714;
 wire net7715;
 wire net7716;
 wire net7717;
 wire net7718;
 wire net7719;
 wire net7720;
 wire net7721;
 wire net7722;
 wire net7723;
 wire net7724;
 wire net7725;
 wire net7726;
 wire net7727;
 wire net7728;
 wire net7729;
 wire net7730;
 wire net7731;
 wire net7732;
 wire net7733;
 wire net7734;
 wire net7735;
 wire net7736;
 wire net7737;
 wire net7738;
 wire net7739;
 wire net7740;
 wire net7741;
 wire net7742;
 wire net7743;
 wire net7744;
 wire net7745;
 wire net7746;
 wire net7747;
 wire net7748;
 wire net7749;
 wire net7750;
 wire net7751;
 wire net7752;
 wire net7753;
 wire net7754;
 wire net7755;
 wire net7756;
 wire net7757;
 wire net7758;
 wire net7759;
 wire net7760;
 wire net7761;
 wire net7762;
 wire net7763;
 wire net7764;
 wire net7765;
 wire net7766;
 wire net7767;
 wire net7768;
 wire net7769;
 wire net7770;
 wire net7771;
 wire net7772;
 wire net7773;
 wire net7774;
 wire net7775;
 wire net7776;
 wire net7777;
 wire net7778;
 wire net7779;
 wire net7780;
 wire net7781;
 wire net7782;
 wire net7783;
 wire net7784;
 wire net7785;
 wire net7786;
 wire net7787;
 wire net7788;
 wire net7789;
 wire net7790;
 wire net7791;
 wire net7792;
 wire net7793;
 wire net7794;
 wire net7795;
 wire net7796;
 wire net7797;
 wire net7798;
 wire net7799;
 wire net7800;
 wire net7801;
 wire net7802;
 wire net7803;
 wire net7804;
 wire net7805;
 wire net7806;
 wire net7807;
 wire net7808;
 wire net7809;
 wire net7810;
 wire net7811;
 wire net7812;
 wire net7813;
 wire net7814;
 wire net7815;
 wire net7816;
 wire net7817;
 wire net7818;
 wire net7819;
 wire net7820;
 wire net7821;
 wire net7822;
 wire net7823;
 wire net7824;
 wire net7825;
 wire net7826;
 wire net7827;
 wire net7828;
 wire net7829;
 wire net7830;
 wire net7831;
 wire net7832;
 wire net7833;
 wire net7834;
 wire net7835;
 wire net7836;
 wire net7837;
 wire net7838;
 wire net7839;
 wire net7840;
 wire net7841;
 wire net7842;
 wire net7843;
 wire net7844;
 wire net7845;
 wire net7846;
 wire net7847;
 wire net7848;
 wire net7849;
 wire net7850;
 wire net7851;
 wire net7852;
 wire net7853;
 wire net7854;
 wire net7855;
 wire net7856;
 wire net7857;
 wire net7858;
 wire net7859;
 wire net7860;
 wire net7861;
 wire net7862;
 wire net7863;
 wire net7864;
 wire net7865;
 wire net7866;
 wire net7867;
 wire net7868;
 wire net7869;
 wire net7870;
 wire net7871;
 wire net7872;
 wire net7873;
 wire net7874;
 wire net7875;
 wire net7876;
 wire net7877;
 wire net7878;
 wire net7879;
 wire net7880;
 wire net7881;
 wire net7882;
 wire net7883;
 wire net7884;
 wire net7885;
 wire net7886;
 wire net7887;
 wire net7888;
 wire net7889;
 wire net7890;
 wire net7891;
 wire net7892;
 wire net7893;
 wire net7894;
 wire net7895;
 wire net7896;
 wire net7897;
 wire net7898;
 wire net7899;
 wire net7900;
 wire net7901;
 wire net7902;
 wire net7903;
 wire net7904;
 wire net7905;
 wire net7906;
 wire net7907;
 wire net7908;
 wire net7909;
 wire net7910;
 wire net7911;
 wire net7912;
 wire net7913;
 wire net7914;
 wire net7915;
 wire net7916;
 wire net7917;
 wire net7918;
 wire net7919;
 wire net7920;
 wire net7921;
 wire net7922;
 wire net7923;
 wire net7924;
 wire net7925;
 wire net7926;
 wire net7927;
 wire net7928;
 wire net7929;
 wire net7930;
 wire net7931;
 wire net7932;
 wire net7933;
 wire net7934;
 wire net7935;
 wire net7936;
 wire net7937;
 wire net7938;
 wire net7939;
 wire net7940;
 wire net7941;
 wire net7942;
 wire net7943;
 wire net7944;
 wire net7945;
 wire net7946;
 wire net7947;
 wire net7948;
 wire net7949;
 wire net7950;
 wire net7951;
 wire net7952;
 wire net7953;
 wire net7954;
 wire net7955;
 wire net7956;
 wire net7957;
 wire net7958;
 wire net7959;
 wire net7960;
 wire net7961;
 wire net7962;
 wire net7963;
 wire net7964;
 wire net7965;
 wire net7966;
 wire net7967;
 wire net7968;
 wire net7969;
 wire net7970;
 wire net7971;
 wire net7972;
 wire net7973;
 wire net7974;
 wire net7975;
 wire net7976;
 wire net7977;
 wire net7978;
 wire net7979;
 wire net7980;
 wire net7981;
 wire net7982;
 wire net7983;
 wire net7984;
 wire net7985;
 wire net7986;
 wire net7987;
 wire net7988;
 wire net7989;
 wire net7990;
 wire net7991;
 wire net7992;
 wire net7993;
 wire net7994;
 wire net7995;
 wire net7996;
 wire net7997;
 wire net7998;
 wire net7999;
 wire net8000;
 wire net8001;
 wire net8002;
 wire net8003;
 wire net8004;
 wire net8005;
 wire net8006;
 wire net8007;
 wire net8008;
 wire net8009;
 wire net8010;
 wire net8011;
 wire net8012;
 wire net8013;
 wire net8014;
 wire net8015;
 wire net8016;
 wire net8017;
 wire net8018;
 wire net8019;
 wire net8020;
 wire net8021;
 wire net8022;
 wire net8023;
 wire net8024;
 wire net8025;
 wire net8026;
 wire net8027;
 wire net8028;
 wire net8029;
 wire net8030;
 wire net8031;
 wire net8032;
 wire net8033;
 wire net8034;
 wire net8035;
 wire net8036;
 wire net8037;
 wire net8038;
 wire net8039;
 wire net8040;
 wire net8041;
 wire net8042;
 wire net8043;
 wire net8044;
 wire net8045;
 wire net8046;
 wire net8047;
 wire net8048;
 wire net8049;
 wire net8050;
 wire net8051;
 wire net8052;
 wire net8053;
 wire net8054;
 wire net8055;
 wire net8056;
 wire net8057;
 wire net8058;
 wire net8059;
 wire net8060;
 wire net8061;
 wire net8062;
 wire net8063;
 wire net8064;
 wire net8065;
 wire net8066;
 wire net8067;
 wire net8068;
 wire net8069;
 wire net8070;
 wire net8071;
 wire net8072;
 wire net8073;
 wire net8074;
 wire net8075;
 wire net8076;
 wire net8077;
 wire net8078;
 wire net8079;
 wire net8080;
 wire net8081;
 wire net8082;
 wire net8083;
 wire net8084;
 wire net8085;
 wire net8086;
 wire net8087;
 wire net8088;
 wire net8089;
 wire net8090;
 wire net8091;
 wire net8092;
 wire net8093;
 wire net8094;
 wire net8095;
 wire net8096;
 wire net8097;
 wire net8098;
 wire net8099;
 wire net8100;
 wire net8101;
 wire net8102;
 wire net8103;
 wire net8104;
 wire net8105;
 wire net8106;
 wire net8107;
 wire net8108;
 wire net8109;
 wire net8110;
 wire net8111;
 wire net8112;
 wire net8113;
 wire net8114;
 wire net8115;
 wire net8116;
 wire net8117;
 wire net8118;
 wire net8119;
 wire net8120;
 wire net8121;
 wire net8122;
 wire net8123;
 wire net8124;
 wire net8125;
 wire net8126;
 wire net8127;
 wire net8128;
 wire net8129;
 wire net8130;
 wire net8131;
 wire net8132;
 wire net8133;
 wire net8134;
 wire net8135;
 wire net8136;
 wire net8137;
 wire net8138;
 wire net8139;
 wire net8140;
 wire net8141;
 wire net8142;
 wire net8143;
 wire net8144;
 wire net8145;
 wire net8146;
 wire net8147;
 wire net8148;
 wire net8149;
 wire net8150;
 wire net8151;
 wire net8152;
 wire net8153;
 wire net8154;
 wire net8155;
 wire net8156;
 wire net8157;
 wire net8158;
 wire net8159;
 wire net8160;
 wire net8161;
 wire net8162;
 wire net8163;
 wire net8164;
 wire net8165;
 wire net8166;
 wire net8167;
 wire net8168;
 wire net8169;
 wire net8170;
 wire net8171;
 wire net8172;
 wire net8173;
 wire net8174;
 wire net8175;
 wire net8176;
 wire net8177;
 wire net8178;
 wire net8179;
 wire net8180;
 wire net8181;
 wire net8182;
 wire net8183;
 wire net8184;
 wire net8185;
 wire net8186;
 wire net8187;
 wire net8188;
 wire net8189;
 wire net8190;
 wire net8191;
 wire net8192;
 wire net8193;
 wire net8194;
 wire net8195;
 wire net8196;
 wire net8197;
 wire net8198;
 wire net8199;
 wire net8200;
 wire net8201;
 wire net8202;
 wire net8203;
 wire net8204;
 wire net8205;
 wire net8206;
 wire net8207;
 wire net8208;
 wire net8209;
 wire net8210;
 wire net8211;
 wire net8212;
 wire net8213;
 wire net8214;
 wire net8215;
 wire net8216;
 wire net8217;
 wire net8218;
 wire net8219;
 wire net8220;
 wire net8221;
 wire net8222;
 wire net8223;
 wire net8224;
 wire net8225;
 wire net8226;
 wire net8227;
 wire net8228;
 wire net8229;
 wire net8230;
 wire net8231;
 wire net8232;
 wire net8233;
 wire net8234;
 wire net8235;
 wire net8236;
 wire net8237;
 wire net8238;
 wire net8239;
 wire net8240;
 wire net8241;
 wire net8242;
 wire net8243;
 wire net8244;
 wire net8245;
 wire net8246;
 wire net8247;
 wire net8248;
 wire net8249;
 wire net8250;
 wire net8251;
 wire net8252;
 wire net8253;
 wire net8254;
 wire net8255;
 wire net8256;
 wire net8257;
 wire net8258;
 wire net8259;
 wire net8260;
 wire net8261;
 wire net8262;
 wire net8263;
 wire net8264;
 wire net8265;
 wire net8266;
 wire net8267;
 wire net8268;
 wire net8269;
 wire net8270;
 wire net8271;
 wire net8272;
 wire net8273;
 wire net8274;
 wire net8275;
 wire net8276;
 wire net8277;
 wire net8278;
 wire net8279;
 wire net8280;
 wire net8281;
 wire net8282;
 wire net8283;
 wire net8284;
 wire net8285;
 wire net8286;
 wire net8287;
 wire net8288;
 wire net8289;
 wire net8290;
 wire net8291;
 wire net8292;
 wire net8293;
 wire net8294;
 wire net8295;
 wire net8296;
 wire net8297;
 wire net8298;
 wire net8299;
 wire net8300;
 wire net8301;
 wire net8302;
 wire net8303;
 wire net8304;
 wire net8305;
 wire net8306;
 wire net8307;
 wire net8308;
 wire net8309;
 wire net8310;
 wire net8311;
 wire net8312;
 wire net8313;
 wire net8314;
 wire net8315;
 wire net8316;
 wire net8317;
 wire net8318;
 wire net8319;
 wire net8320;
 wire net8321;
 wire net8322;
 wire net8323;
 wire net8324;
 wire net8325;
 wire net8326;
 wire net8327;
 wire net8328;
 wire net8329;
 wire net8330;
 wire net8331;
 wire net8332;
 wire net8333;
 wire net8334;
 wire net8335;
 wire net8336;
 wire net8337;
 wire net8338;
 wire net8339;
 wire net8340;
 wire net8341;
 wire net8342;
 wire net8343;
 wire net8344;
 wire net8345;
 wire net8346;
 wire net8347;
 wire net8348;
 wire net8349;
 wire net8350;
 wire net8351;
 wire net8352;
 wire net8353;
 wire net8354;
 wire net8355;
 wire net8356;
 wire net8357;
 wire net8358;
 wire net8359;
 wire net8360;
 wire net8361;
 wire net8362;
 wire net8363;
 wire net8364;
 wire net8365;
 wire net8366;
 wire net8367;
 wire net8368;
 wire net8369;
 wire net8370;
 wire net8371;
 wire net8372;
 wire net8373;
 wire net8374;
 wire net8375;
 wire net8376;
 wire net8377;
 wire net8378;
 wire net8379;
 wire net8380;
 wire net8381;
 wire net8382;
 wire net8383;
 wire net8384;
 wire net8385;
 wire net8386;
 wire net8387;
 wire net8388;
 wire net8389;
 wire net8390;
 wire net8391;
 wire net8392;
 wire net8393;
 wire net8394;
 wire net8395;
 wire net8396;
 wire net8397;
 wire net8398;
 wire net8399;
 wire net8400;
 wire net8401;
 wire net8402;
 wire net8403;
 wire net8404;
 wire net8405;
 wire net8406;
 wire net8407;
 wire net8408;
 wire net8409;
 wire net8410;
 wire net8411;
 wire net8412;
 wire net8413;
 wire net8414;
 wire net8415;
 wire net8416;
 wire net8417;
 wire net8418;
 wire net8419;
 wire net8420;
 wire net8421;
 wire net8422;
 wire net8423;
 wire net8424;
 wire net8425;
 wire net8426;
 wire net8427;
 wire net8428;
 wire net8429;
 wire net8430;
 wire net8431;
 wire net8432;
 wire net8433;
 wire net8434;
 wire net8435;
 wire net8436;
 wire net8437;
 wire net8438;
 wire net8439;
 wire net8440;
 wire net8441;
 wire net8442;
 wire net8443;
 wire net8444;
 wire net8445;
 wire net8446;
 wire net8447;
 wire net8448;
 wire net8449;
 wire net8450;
 wire net8451;
 wire net8452;
 wire net8453;
 wire net8454;
 wire net8455;
 wire net8456;
 wire net8457;
 wire net8458;
 wire net8459;
 wire net8460;
 wire net8461;
 wire net8462;
 wire net8463;
 wire net8464;
 wire net8465;
 wire net8466;
 wire net8467;
 wire net8468;
 wire net8469;
 wire net8470;
 wire net8471;
 wire net8472;
 wire net8473;
 wire net8474;
 wire net8475;
 wire net8476;
 wire net8477;
 wire net8478;
 wire net8479;
 wire net8480;
 wire net8481;
 wire net8482;
 wire net8483;
 wire net8484;
 wire net8485;
 wire net8486;
 wire net8487;
 wire net8488;
 wire net8489;
 wire net8490;
 wire net8491;
 wire net8492;
 wire net8493;
 wire net8494;
 wire net8495;
 wire net8496;
 wire net8497;
 wire net8498;
 wire net8499;
 wire net8500;
 wire net8501;
 wire net8502;
 wire net8503;
 wire net8504;
 wire net8505;
 wire net8506;
 wire net8507;
 wire net8508;
 wire net8509;
 wire net8510;
 wire net8511;
 wire net8512;
 wire net8513;
 wire net8514;
 wire net8515;
 wire net8516;
 wire net8517;
 wire net8518;
 wire net8519;
 wire net8520;
 wire net8521;
 wire net8522;
 wire net8523;
 wire net8524;
 wire net8525;
 wire net8526;
 wire net8527;
 wire net8528;
 wire net8529;
 wire net8530;
 wire net8531;
 wire net8532;
 wire net8533;
 wire net8534;
 wire net8535;
 wire net8536;
 wire net8537;
 wire net8538;
 wire net8539;
 wire net8540;
 wire net8541;
 wire net8542;
 wire net8543;
 wire net8544;
 wire net8545;
 wire net8546;
 wire net8547;
 wire net8548;
 wire net8549;
 wire net8550;
 wire net8551;
 wire net8552;
 wire net8553;
 wire net8554;
 wire net8555;
 wire net8556;
 wire net8557;
 wire net8558;
 wire net8559;
 wire net8560;
 wire net8561;
 wire net8562;
 wire net8563;
 wire net8564;
 wire net8565;
 wire net8566;
 wire net8567;
 wire net8568;
 wire net8569;
 wire net8570;
 wire net8571;
 wire net8572;
 wire net8573;
 wire net8574;
 wire net8575;
 wire net8576;
 wire net8577;
 wire net8578;
 wire net8579;
 wire net8580;
 wire net8581;
 wire net8582;
 wire net8583;
 wire net8584;
 wire net8585;
 wire net8586;
 wire net8587;
 wire net8588;
 wire net8589;
 wire net8590;
 wire net8591;
 wire net8592;
 wire net8593;
 wire net8594;
 wire net8595;
 wire net8596;
 wire net8597;
 wire net8598;
 wire net8599;
 wire net8600;
 wire net8601;
 wire net8602;
 wire net8603;
 wire net8604;
 wire net8605;
 wire net8606;
 wire net8607;
 wire net8608;
 wire net8609;
 wire net8610;
 wire net8611;
 wire net8612;
 wire net8613;
 wire net8614;
 wire net8615;
 wire net8616;
 wire net8617;
 wire net8618;
 wire net8619;
 wire net8620;
 wire net8621;
 wire net8622;
 wire net8623;
 wire net8624;
 wire net8625;
 wire net8626;
 wire net8627;
 wire net8628;
 wire net8629;
 wire net8630;
 wire net8631;
 wire net8632;
 wire net8633;
 wire net8634;
 wire net8635;
 wire net8636;
 wire net8637;
 wire net8638;
 wire net8639;
 wire net8640;
 wire net8641;
 wire net8642;
 wire net8643;
 wire net8644;
 wire net8645;
 wire net8646;
 wire net8647;
 wire net8648;
 wire net8649;
 wire net8650;
 wire net8651;
 wire net8652;
 wire net8653;
 wire net8654;
 wire net8655;
 wire net8656;
 wire net8657;
 wire net8658;
 wire net8659;
 wire net8660;
 wire net8661;
 wire net8662;
 wire net8663;
 wire net8664;
 wire net8665;
 wire net8666;
 wire net8667;
 wire net8668;
 wire net8669;
 wire net8670;
 wire net8671;
 wire net8672;
 wire net8673;
 wire net8674;
 wire net8675;
 wire net8676;
 wire net8677;
 wire net8678;
 wire net8679;
 wire net8680;
 wire net8681;
 wire net8682;
 wire net8683;
 wire net8684;
 wire net8685;
 wire net8686;
 wire net8687;
 wire net8688;
 wire net8689;
 wire net8690;
 wire net8691;
 wire net8692;
 wire net8693;
 wire net8694;
 wire net8695;
 wire net8696;
 wire net8697;
 wire net8698;
 wire net8699;
 wire net8700;
 wire net8701;
 wire net8702;
 wire net8703;
 wire net8704;
 wire net8705;
 wire net8706;
 wire net8707;
 wire net8708;
 wire net8709;
 wire net8710;
 wire net8711;
 wire net8712;
 wire net8713;
 wire net8714;
 wire net8715;
 wire net8716;
 wire net8717;
 wire net8718;
 wire net8719;
 wire net8720;
 wire net8721;
 wire net8722;
 wire net8723;
 wire net8724;
 wire net8725;
 wire net8726;
 wire net8727;
 wire net8728;
 wire net8729;
 wire net8730;
 wire net8731;
 wire net8732;
 wire net8733;
 wire net8734;
 wire net8735;
 wire net8736;
 wire net8737;
 wire net8738;
 wire net8739;
 wire net8740;
 wire net8741;
 wire net8742;
 wire net8743;
 wire net8744;
 wire net8745;
 wire net8746;
 wire net8747;
 wire net8748;
 wire net8749;
 wire net8750;
 wire net8751;
 wire net8752;
 wire net8753;
 wire net8754;
 wire net8755;
 wire net8756;
 wire net8757;
 wire net8758;
 wire net8759;
 wire net8760;
 wire net8761;
 wire net8762;
 wire net8763;
 wire net8764;
 wire net8765;
 wire net8766;
 wire net8767;
 wire net8768;
 wire net8769;
 wire net8770;
 wire net8771;
 wire net8772;
 wire net8773;
 wire net8774;
 wire net8775;
 wire net8776;
 wire net8777;
 wire net8778;
 wire net8779;
 wire net8780;
 wire net8781;
 wire net8782;
 wire net8783;
 wire net8784;
 wire net8785;
 wire net8786;
 wire net8787;
 wire net8788;
 wire net8789;
 wire net8790;
 wire net8791;
 wire net8792;
 wire net8793;
 wire net8794;
 wire net8795;
 wire net8796;
 wire net8797;
 wire net8798;
 wire net8799;
 wire net8800;
 wire net8801;
 wire net8802;
 wire net8803;
 wire net8804;
 wire net8805;
 wire net8806;
 wire net8807;
 wire net8808;
 wire net8809;
 wire net8810;
 wire net8811;
 wire net8812;
 wire net8813;
 wire net8814;
 wire net8815;
 wire net8816;
 wire net8817;
 wire net8818;
 wire net8819;
 wire net8820;
 wire net8821;
 wire net8822;
 wire net8823;
 wire net8824;
 wire net8825;
 wire net8826;
 wire net8827;
 wire net8828;
 wire net8829;
 wire net8830;
 wire net8831;
 wire net8832;
 wire net8833;
 wire net8834;
 wire net8835;
 wire net8836;
 wire net8837;
 wire net8838;
 wire net8839;
 wire net8840;
 wire net8841;
 wire net8842;
 wire net8843;
 wire net8844;
 wire net8845;
 wire net8846;
 wire net8847;
 wire net8848;
 wire net8849;
 wire net8850;
 wire net8851;
 wire net8852;
 wire net8853;
 wire net8854;
 wire net8855;
 wire net8856;
 wire net8857;
 wire net8858;
 wire net8859;
 wire net8860;
 wire net8861;
 wire net8862;
 wire net8863;
 wire net8864;
 wire net8865;
 wire net8866;
 wire net8867;
 wire net8868;
 wire net8869;
 wire net8870;
 wire net8871;
 wire net8872;
 wire net8873;
 wire net8874;
 wire net8875;
 wire net8876;
 wire net8877;
 wire net8878;
 wire net8879;
 wire net8880;
 wire net8881;
 wire net8882;
 wire net8883;
 wire net8884;
 wire net8885;
 wire net8886;
 wire net8887;
 wire net8888;
 wire net8889;
 wire net8890;
 wire net8891;
 wire net8892;
 wire net8893;
 wire net8894;
 wire net8895;
 wire net8896;
 wire net8897;
 wire net8898;
 wire net8899;
 wire net8900;
 wire net8901;
 wire net8902;
 wire net8903;
 wire net8904;
 wire net8905;
 wire net8906;
 wire net8907;
 wire net8908;
 wire net8909;
 wire net8910;
 wire net8911;
 wire net8912;
 wire net8913;
 wire net8914;
 wire net8915;
 wire net8916;
 wire net8917;
 wire net8918;
 wire net8919;
 wire net8920;
 wire net8921;
 wire net8922;
 wire net8923;
 wire net8924;
 wire net8925;
 wire net8926;
 wire net8927;
 wire net8928;
 wire net8929;
 wire net8930;
 wire net8931;
 wire net8932;
 wire net8933;
 wire net8934;
 wire net8935;
 wire net8936;
 wire net8937;
 wire net8938;
 wire net8939;
 wire net8940;
 wire net8941;
 wire net8942;
 wire net8943;
 wire net8944;
 wire net8945;
 wire net8946;
 wire net8947;
 wire net8948;
 wire net8949;
 wire net8950;
 wire net8951;
 wire net8952;
 wire net8953;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_4_0__leaf_clk;
 wire clknet_4_1__leaf_clk;
 wire clknet_4_2__leaf_clk;
 wire clknet_4_3__leaf_clk;
 wire clknet_4_4__leaf_clk;
 wire clknet_4_5__leaf_clk;
 wire clknet_4_6__leaf_clk;
 wire clknet_4_7__leaf_clk;
 wire clknet_4_8__leaf_clk;
 wire clknet_4_9__leaf_clk;
 wire clknet_4_10__leaf_clk;
 wire clknet_4_11__leaf_clk;
 wire clknet_4_12__leaf_clk;
 wire clknet_4_13__leaf_clk;
 wire clknet_4_14__leaf_clk;
 wire clknet_4_15__leaf_clk;
 wire net8954;
 wire net8955;
 wire net8956;
 wire net8957;
 wire net8958;
 wire net8959;
 wire net8960;
 wire net8961;
 wire net8962;
 wire net8963;
 wire net8964;
 wire net8965;
 wire net8966;
 wire net8967;
 wire net8968;
 wire net8969;
 wire net8970;
 wire net8971;
 wire net8972;
 wire net8973;
 wire net8974;
 wire net8975;
 wire net8976;
 wire net8977;
 wire net8978;
 wire net8979;
 wire net8980;
 wire net8981;
 wire net8982;
 wire net8983;
 wire net8984;
 wire net8985;
 wire net8986;
 wire net8987;
 wire net8988;
 wire net8989;
 wire net8990;
 wire net8991;
 wire net8992;
 wire net8993;
 wire net8994;
 wire net8995;
 wire net8996;
 wire net8997;
 wire net8998;
 wire net8999;
 wire net9000;
 wire net9001;
 wire net9002;
 wire net9003;
 wire net9004;
 wire net9005;
 wire net9006;
 wire net9007;
 wire net9008;
 wire net9009;
 wire net9010;
 wire net9011;
 wire net9012;
 wire net9013;
 wire net9014;
 wire net9015;
 wire net9016;
 wire net9017;
 wire net9018;
 wire net9019;
 wire net9020;
 wire net9021;
 wire net9022;
 wire net9023;
 wire net9024;
 wire net9025;
 wire net9026;
 wire net9027;
 wire net9028;
 wire net9029;
 wire net9030;
 wire net9031;
 wire net9032;
 wire net9033;
 wire net9034;
 wire net9035;
 wire net9036;
 wire net9037;
 wire net9038;
 wire net9039;
 wire net9040;
 wire net9041;
 wire net9042;
 wire net9043;
 wire net9044;
 wire net9045;
 wire net9046;
 wire net9047;
 wire net9048;
 wire net9049;
 wire net9050;
 wire net9051;
 wire net9052;
 wire net9053;
 wire net9054;
 wire net9055;
 wire net9056;
 wire net9057;
 wire net9058;
 wire net9059;
 wire net9060;
 wire net9061;
 wire net9062;
 wire net9063;
 wire net9064;
 wire net9065;
 wire net9066;
 wire net9067;
 wire net9068;
 wire net9069;
 wire net9070;
 wire net9071;
 wire net9072;
 wire net9073;
 wire net9074;
 wire net9075;
 wire net9076;
 wire net9077;
 wire net9078;
 wire net9079;
 wire net9080;
 wire net9081;
 wire net9082;
 wire net9083;
 wire net9084;
 wire net9085;
 wire net9086;
 wire net9087;
 wire net9088;
 wire net9089;
 wire net9090;
 wire net9091;
 wire net9092;
 wire net9093;
 wire net9094;
 wire net9095;
 wire net9096;
 wire net9097;
 wire net9098;
 wire net9099;
 wire net9100;
 wire net9101;
 wire net9102;
 wire net9103;
 wire net9104;
 wire net9105;
 wire net9106;
 wire net9107;
 wire net9108;
 wire net9109;
 wire net9110;
 wire net9111;
 wire net9112;
 wire net9113;
 wire net9114;
 wire net9115;
 wire net9116;
 wire net9117;
 wire net9118;
 wire net9119;
 wire net9120;
 wire net9121;
 wire net9122;
 wire net9123;
 wire net9124;
 wire net9125;
 wire net9126;
 wire net9127;
 wire net9128;
 wire net9129;
 wire net9130;
 wire net9131;
 wire net9132;
 wire net9133;
 wire net9134;
 wire net9135;
 wire net9136;
 wire net9137;
 wire net9138;
 wire net9139;
 wire net9140;
 wire net9141;
 wire net9142;
 wire net9143;
 wire net9144;
 wire net9145;
 wire net9146;
 wire net9147;
 wire net9148;
 wire net9149;
 wire net9150;
 wire net9151;
 wire net9152;
 wire net9153;
 wire net9154;
 wire net9155;
 wire net9156;
 wire net9157;
 wire net9158;
 wire net9159;
 wire net9160;
 wire net9161;
 wire net9162;
 wire net9163;
 wire net9164;
 wire net9165;
 wire net9166;
 wire net9167;
 wire net9168;
 wire net9169;
 wire net9170;
 wire net9171;
 wire net9172;
 wire net9173;
 wire net9174;
 wire net9175;
 wire net9176;
 wire net9177;
 wire net9178;
 wire net9179;
 wire net9180;
 wire net9181;
 wire net9182;
 wire net9183;
 wire net9184;
 wire net9185;
 wire net9186;
 wire net9187;
 wire net9188;
 wire net9189;
 wire net9190;
 wire net9191;
 wire net9192;
 wire net9193;
 wire net9194;
 wire net9195;
 wire net9196;
 wire net9197;
 wire net9198;
 wire net9199;
 wire net9200;
 wire net9201;
 wire net9202;
 wire net9203;
 wire net9204;
 wire net9205;
 wire net9206;
 wire net9207;
 wire net9208;
 wire net9209;
 wire net9210;
 wire net9211;
 wire net9212;
 wire net9213;
 wire net9214;
 wire net9215;
 wire net9216;
 wire net9217;
 wire net9218;
 wire net9219;
 wire net9220;
 wire net9221;
 wire net9222;
 wire net9223;
 wire net9224;
 wire net9225;
 wire net9226;
 wire net9227;
 wire net9228;
 wire net9229;
 wire net9230;
 wire net9231;
 wire net9232;
 wire net9233;
 wire net9234;
 wire net9235;
 wire net9236;
 wire net9237;
 wire net9238;
 wire net9239;
 wire net9240;
 wire net9241;
 wire net9242;
 wire net9243;
 wire net9244;
 wire net9245;
 wire net9246;
 wire net9247;
 wire net9248;

 sky130_fd_sc_hd__inv_2 _12564_ (.A(\matmul0.start ),
    .Y(_04854_));
 sky130_fd_sc_hd__and2_1 _12565_ (.A(net6748),
    .B(net6598),
    .X(_04855_));
 sky130_fd_sc_hd__buf_2 _12566_ (.A(_04855_),
    .X(_04856_));
 sky130_fd_sc_hd__buf_1 _12567_ (.A(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__clkbuf_1 _12568_ (.A(net3031),
    .X(_04858_));
 sky130_fd_sc_hd__buf_1 _12569_ (.A(net2388),
    .X(_04859_));
 sky130_fd_sc_hd__buf_1 _12570_ (.A(net1987),
    .X(_04860_));
 sky130_fd_sc_hd__a21o_1 _12571_ (.A1(net9150),
    .A2(_04854_),
    .B1(net1622),
    .X(_00013_));
 sky130_fd_sc_hd__inv_2 _12572_ (.A(net7531),
    .Y(_04861_));
 sky130_fd_sc_hd__or2b_1 _12573_ (.A(net7478),
    .B_N(net8863),
    .X(_04862_));
 sky130_fd_sc_hd__a21o_1 _12574_ (.A1(net4313),
    .A2(\pid_q.state[0] ),
    .B1(_04862_),
    .X(_00016_));
 sky130_fd_sc_hd__inv_2 _12575_ (.A(\matmul0.matmul_stage_inst.start ),
    .Y(_04863_));
 sky130_fd_sc_hd__a21o_1 _12576_ (.A1(net9148),
    .A2(_04863_),
    .B1(net6597),
    .X(_00012_));
 sky130_fd_sc_hd__inv_2 _12577_ (.A(net6597),
    .Y(_04864_));
 sky130_fd_sc_hd__a21o_1 _12578_ (.A1(\matmul0.state[1] ),
    .A2(_04864_),
    .B1(net8976),
    .X(_00014_));
 sky130_fd_sc_hd__inv_2 _12579_ (.A(net8906),
    .Y(_04865_));
 sky130_fd_sc_hd__clkbuf_1 _12580_ (.A(_04865_),
    .X(_04866_));
 sky130_fd_sc_hd__buf_1 _12581_ (.A(net4309),
    .X(_04867_));
 sky130_fd_sc_hd__a211o_1 _12582_ (.A1(net4311),
    .A2(\pid_d.state[0] ),
    .B1(net4327),
    .C1(_04867_),
    .X(_00015_));
 sky130_fd_sc_hd__and2_1 _12583_ (.A(net8863),
    .B(net7496),
    .X(_04868_));
 sky130_fd_sc_hd__buf_1 _12584_ (.A(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__clkbuf_1 _12585_ (.A(net3716),
    .X(_04870_));
 sky130_fd_sc_hd__buf_1 _12586_ (.A(net3019),
    .X(_00011_));
 sky130_fd_sc_hd__and2_1 _12587_ (.A(net8864),
    .B(net7521),
    .X(_04871_));
 sky130_fd_sc_hd__clkbuf_1 _12588_ (.A(_04871_),
    .X(_00010_));
 sky130_fd_sc_hd__inv_2 _12589_ (.A(net4365),
    .Y(_04872_));
 sky130_fd_sc_hd__nor2_1 _12590_ (.A(_04865_),
    .B(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__clkbuf_1 _12591_ (.A(net3709),
    .X(_04874_));
 sky130_fd_sc_hd__clkbuf_1 _12592_ (.A(net3016),
    .X(_00006_));
 sky130_fd_sc_hd__inv_2 _12593_ (.A(net4384),
    .Y(_04875_));
 sky130_fd_sc_hd__nor2_1 _12594_ (.A(_04865_),
    .B(net4293),
    .Y(_00005_));
 sky130_fd_sc_hd__nand2_1 _12595_ (.A(\matmul0.state[0] ),
    .B(\matmul0.start ),
    .Y(_04876_));
 sky130_fd_sc_hd__buf_1 _12596_ (.A(net4292),
    .X(_04877_));
 sky130_fd_sc_hd__inv_2 _12597_ (.A(_04877_),
    .Y(_00001_));
 sky130_fd_sc_hd__and3_1 _12598_ (.A(net7531),
    .B(net8904),
    .C(net4389),
    .X(_04878_));
 sky130_fd_sc_hd__clkbuf_1 _12599_ (.A(_04878_),
    .X(_00004_));
 sky130_fd_sc_hd__and2_1 _12600_ (.A(net8864),
    .B(net7463),
    .X(_04879_));
 sky130_fd_sc_hd__clkbuf_1 _12601_ (.A(_04879_),
    .X(_00007_));
 sky130_fd_sc_hd__and3_1 _12602_ (.A(net8864),
    .B(net7530),
    .C(\pid_q.state[0] ),
    .X(_04880_));
 sky130_fd_sc_hd__clkbuf_1 _12603_ (.A(_04880_),
    .X(_00009_));
 sky130_fd_sc_hd__and2_1 _12604_ (.A(net8872),
    .B(net7490),
    .X(_04881_));
 sky130_fd_sc_hd__clkbuf_1 _12605_ (.A(_04881_),
    .X(_04882_));
 sky130_fd_sc_hd__buf_1 _12606_ (.A(net3699),
    .X(_00008_));
 sky130_fd_sc_hd__nand2_1 _12607_ (.A(\matmul0.matmul_stage_inst.state[0] ),
    .B(\matmul0.matmul_stage_inst.start ),
    .Y(_04883_));
 sky130_fd_sc_hd__inv_2 _12608_ (.A(net4279),
    .Y(_04884_));
 sky130_fd_sc_hd__clkbuf_1 _12609_ (.A(net3697),
    .X(_00000_));
 sky130_fd_sc_hd__and2_1 _12610_ (.A(net8909),
    .B(net4341),
    .X(_04885_));
 sky130_fd_sc_hd__clkbuf_2 _12611_ (.A(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__clkbuf_1 _12612_ (.A(net3696),
    .X(_00003_));
 sky130_fd_sc_hd__inv_2 _12613_ (.A(net4315),
    .Y(_04887_));
 sky130_fd_sc_hd__nor2_1 _12614_ (.A(_04865_),
    .B(_04887_),
    .Y(_00002_));
 sky130_fd_sc_hd__and3b_1 _12615_ (.A_N(net6664),
    .B(net6673),
    .C(net6678),
    .X(_04888_));
 sky130_fd_sc_hd__buf_6 _12616_ (.A(_04888_),
    .X(_04889_));
 sky130_fd_sc_hd__clkbuf_1 _12617_ (.A(_04889_),
    .X(_04890_));
 sky130_fd_sc_hd__clkbuf_1 _12618_ (.A(net2992),
    .X(_04891_));
 sky130_fd_sc_hd__buf_6 _12619_ (.A(_04856_),
    .X(_04892_));
 sky130_fd_sc_hd__nor3b_1 _12620_ (.A(net6664),
    .B(net6673),
    .C_N(net6678),
    .Y(_04893_));
 sky130_fd_sc_hd__clkbuf_2 _12621_ (.A(_04893_),
    .X(_04894_));
 sky130_fd_sc_hd__nand3_1 _12622_ (.A(net7314),
    .B(_04892_),
    .C(net3695),
    .Y(_04895_));
 sky130_fd_sc_hd__nor3b_1 _12623_ (.A(net6664),
    .B(net6678),
    .C_N(net6673),
    .Y(_04896_));
 sky130_fd_sc_hd__buf_6 _12624_ (.A(_04896_),
    .X(_04897_));
 sky130_fd_sc_hd__and3_1 _12625_ (.A(net6749),
    .B(net6599),
    .C(net5268),
    .X(_04898_));
 sky130_fd_sc_hd__a22oi_1 _12626_ (.A1(\svm0.vC[5] ),
    .A2(net2990),
    .B1(net3694),
    .B2(net4275),
    .Y(_04899_));
 sky130_fd_sc_hd__and2_1 _12627_ (.A(_04895_),
    .B(net2367),
    .X(_04900_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _12628_ (.A(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__clkbuf_1 _12629_ (.A(net1618),
    .X(_04902_));
 sky130_fd_sc_hd__nand2_1 _12630_ (.A(net7881),
    .B(net1356),
    .Y(_04903_));
 sky130_fd_sc_hd__nand3_1 _12631_ (.A(net7325),
    .B(_04892_),
    .C(net4278),
    .Y(_04904_));
 sky130_fd_sc_hd__clkbuf_1 _12632_ (.A(_04904_),
    .X(_04905_));
 sky130_fd_sc_hd__a32oi_1 _12633_ (.A1(net5276),
    .A2(_04856_),
    .A3(_04897_),
    .B1(_04889_),
    .B2(\svm0.vC[4] ),
    .Y(_04906_));
 sky130_fd_sc_hd__clkbuf_1 _12634_ (.A(net2989),
    .X(_04907_));
 sky130_fd_sc_hd__and3_1 _12635_ (.A(net7852),
    .B(net1985),
    .C(net2363),
    .X(_04908_));
 sky130_fd_sc_hd__clkbuf_1 _12636_ (.A(_04894_),
    .X(_04909_));
 sky130_fd_sc_hd__nand3_1 _12637_ (.A(net7337),
    .B(net3030),
    .C(net2988),
    .Y(_04910_));
 sky130_fd_sc_hd__and3_1 _12638_ (.A(net6750),
    .B(net6600),
    .C(net5284),
    .X(_04911_));
 sky130_fd_sc_hd__a22oi_1 _12639_ (.A1(\svm0.vC[3] ),
    .A2(net2990),
    .B1(net3694),
    .B2(net4269),
    .Y(_04912_));
 sky130_fd_sc_hd__clkbuf_1 _12640_ (.A(net2354),
    .X(_04913_));
 sky130_fd_sc_hd__and3_1 _12641_ (.A(net7825),
    .B(net2357),
    .C(net1979),
    .X(_04914_));
 sky130_fd_sc_hd__xnor2_1 _12642_ (.A(_04908_),
    .B(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__xnor2_2 _12643_ (.A(_04903_),
    .B(_04915_),
    .Y(_04916_));
 sky130_fd_sc_hd__nand3_1 _12644_ (.A(net7341),
    .B(net3030),
    .C(net3695),
    .Y(_04917_));
 sky130_fd_sc_hd__a32oi_1 _12645_ (.A1(net5295),
    .A2(_04892_),
    .A3(net3694),
    .B1(net2990),
    .B2(\svm0.vC[2] ),
    .Y(_04918_));
 sky130_fd_sc_hd__and2_1 _12646_ (.A(net2353),
    .B(net2348),
    .X(_04919_));
 sky130_fd_sc_hd__buf_1 _12647_ (.A(_04919_),
    .X(_04920_));
 sky130_fd_sc_hd__clkbuf_1 _12648_ (.A(net1616),
    .X(_04921_));
 sky130_fd_sc_hd__nand2_1 _12649_ (.A(net7813),
    .B(net1346),
    .Y(_04922_));
 sky130_fd_sc_hd__nand3_1 _12650_ (.A(net7362),
    .B(net3030),
    .C(net3695),
    .Y(_04923_));
 sky130_fd_sc_hd__buf_1 _12651_ (.A(net2344),
    .X(_04924_));
 sky130_fd_sc_hd__a32oi_1 _12652_ (.A1(net5304),
    .A2(_04892_),
    .A3(net3694),
    .B1(net2990),
    .B2(\svm0.vC[1] ),
    .Y(_04925_));
 sky130_fd_sc_hd__buf_1 _12653_ (.A(net2341),
    .X(_04926_));
 sky130_fd_sc_hd__and3_1 _12654_ (.A(net7797),
    .B(_04924_),
    .C(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__and3_1 _12655_ (.A(net6751),
    .B(net6600),
    .C(net5308),
    .X(_04928_));
 sky130_fd_sc_hd__nand2_1 _12656_ (.A(net3693),
    .B(net4266),
    .Y(_04929_));
 sky130_fd_sc_hd__clkbuf_1 _12657_ (.A(net2977),
    .X(_04930_));
 sky130_fd_sc_hd__a32oi_1 _12658_ (.A1(net7364),
    .A2(_04892_),
    .A3(net4278),
    .B1(net2990),
    .B2(\svm0.vC[0] ),
    .Y(_04931_));
 sky130_fd_sc_hd__buf_1 _12659_ (.A(net2335),
    .X(_04932_));
 sky130_fd_sc_hd__and3_1 _12660_ (.A(net7760),
    .B(net2340),
    .C(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__xnor2_1 _12661_ (.A(_04927_),
    .B(_04933_),
    .Y(_04934_));
 sky130_fd_sc_hd__xnor2_2 _12662_ (.A(_04922_),
    .B(_04934_),
    .Y(_04935_));
 sky130_fd_sc_hd__and3_1 _12663_ (.A(net7813),
    .B(_04924_),
    .C(_04926_),
    .X(_04936_));
 sky130_fd_sc_hd__and3_1 _12664_ (.A(net7777),
    .B(net2340),
    .C(_04932_),
    .X(_04937_));
 sky130_fd_sc_hd__o211a_1 _12665_ (.A1(_04936_),
    .A2(_04937_),
    .B1(net7836),
    .C1(net1346),
    .X(_04938_));
 sky130_fd_sc_hd__a21oi_2 _12666_ (.A1(_04936_),
    .A2(_04937_),
    .B1(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__xnor2_1 _12667_ (.A(_04935_),
    .B(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__xnor2_2 _12668_ (.A(_04916_),
    .B(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__and3_1 _12669_ (.A(net7836),
    .B(net1974),
    .C(net1971),
    .X(_04942_));
 sky130_fd_sc_hd__and3_1 _12670_ (.A(net7813),
    .B(net2338),
    .C(net1968),
    .X(_04943_));
 sky130_fd_sc_hd__o211a_1 _12671_ (.A1(_04942_),
    .A2(_04943_),
    .B1(net7853),
    .C1(net1615),
    .X(_04944_));
 sky130_fd_sc_hd__a21o_2 _12672_ (.A1(_04942_),
    .A2(_04943_),
    .B1(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__nand2_1 _12673_ (.A(net7836),
    .B(net1346),
    .Y(_04946_));
 sky130_fd_sc_hd__xor2_1 _12674_ (.A(_04936_),
    .B(_04937_),
    .X(_04947_));
 sky130_fd_sc_hd__xnor2_1 _12675_ (.A(_04946_),
    .B(_04947_),
    .Y(_04948_));
 sky130_fd_sc_hd__and3_1 _12676_ (.A(net7844),
    .B(net2356),
    .C(net1978),
    .X(_04949_));
 sky130_fd_sc_hd__and3_1 _12677_ (.A(net7915),
    .B(net2368),
    .C(net2365),
    .X(_04950_));
 sky130_fd_sc_hd__and3_1 _12678_ (.A(net7881),
    .B(net1981),
    .C(net2359),
    .X(_04951_));
 sky130_fd_sc_hd__xnor2_1 _12679_ (.A(_04950_),
    .B(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__xnor2_2 _12680_ (.A(_04949_),
    .B(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__o21a_1 _12681_ (.A1(_04945_),
    .A2(net1008),
    .B1(_04953_),
    .X(_04954_));
 sky130_fd_sc_hd__a21oi_4 _12682_ (.A1(_04945_),
    .A2(net1008),
    .B1(_04954_),
    .Y(_04955_));
 sky130_fd_sc_hd__nand3_1 _12683_ (.A(net7283),
    .B(_04856_),
    .C(net4278),
    .Y(_04956_));
 sky130_fd_sc_hd__clkbuf_1 _12684_ (.A(net2976),
    .X(_04957_));
 sky130_fd_sc_hd__a32oi_1 _12685_ (.A1(net5255),
    .A2(_04856_),
    .A3(net4277),
    .B1(_04889_),
    .B2(\svm0.vC[7] ),
    .Y(_04958_));
 sky130_fd_sc_hd__buf_1 _12686_ (.A(net2974),
    .X(_04959_));
 sky130_fd_sc_hd__and2_1 _12687_ (.A(net2330),
    .B(net2325),
    .X(_04960_));
 sky130_fd_sc_hd__nand2_1 _12688_ (.A(net7948),
    .B(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__nand3_1 _12689_ (.A(net7303),
    .B(_04856_),
    .C(net4278),
    .Y(_04962_));
 sky130_fd_sc_hd__a32oi_1 _12690_ (.A1(net5263),
    .A2(_04856_),
    .A3(net4277),
    .B1(_04889_),
    .B2(\svm0.vC[6] ),
    .Y(_04963_));
 sky130_fd_sc_hd__and2_1 _12691_ (.A(net2973),
    .B(net2972),
    .X(_04964_));
 sky130_fd_sc_hd__clkbuf_1 _12692_ (.A(_04964_),
    .X(_04965_));
 sky130_fd_sc_hd__nand2_1 _12693_ (.A(net7905),
    .B(net1963),
    .Y(_04966_));
 sky130_fd_sc_hd__xnor2_1 _12694_ (.A(_04961_),
    .B(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__a21o_1 _12695_ (.A1(_04950_),
    .A2(_04951_),
    .B1(_04949_),
    .X(_04968_));
 sky130_fd_sc_hd__o21ai_2 _12696_ (.A1(_04950_),
    .A2(_04951_),
    .B1(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__xnor2_1 _12697_ (.A(net1343),
    .B(_04969_),
    .Y(_04970_));
 sky130_fd_sc_hd__xnor2_1 _12698_ (.A(_04955_),
    .B(_04970_),
    .Y(_04971_));
 sky130_fd_sc_hd__xnor2_1 _12699_ (.A(_04941_),
    .B(_04971_),
    .Y(_04972_));
 sky130_fd_sc_hd__inv_2 _12700_ (.A(net7943),
    .Y(_04973_));
 sky130_fd_sc_hd__clkbuf_1 _12701_ (.A(net2973),
    .X(_04974_));
 sky130_fd_sc_hd__clkbuf_1 _12702_ (.A(net2972),
    .X(_04975_));
 sky130_fd_sc_hd__nand2_1 _12703_ (.A(net2323),
    .B(net2319),
    .Y(_04976_));
 sky130_fd_sc_hd__nor2_1 _12704_ (.A(net4260),
    .B(net1960),
    .Y(_04977_));
 sky130_fd_sc_hd__xnor2_2 _12705_ (.A(_04945_),
    .B(_04953_),
    .Y(_04978_));
 sky130_fd_sc_hd__xnor2_4 _12706_ (.A(net1008),
    .B(_04978_),
    .Y(_04979_));
 sky130_fd_sc_hd__and3_2 _12707_ (.A(net7854),
    .B(net1974),
    .C(net1971),
    .X(_04980_));
 sky130_fd_sc_hd__and3_2 _12708_ (.A(net7826),
    .B(net2338),
    .C(net1968),
    .X(_04981_));
 sky130_fd_sc_hd__and3_1 _12709_ (.A(net7883),
    .B(net2351),
    .C(net2347),
    .X(_04982_));
 sky130_fd_sc_hd__a21o_1 _12710_ (.A1(_04980_),
    .A2(_04981_),
    .B1(_04982_),
    .X(_04983_));
 sky130_fd_sc_hd__o21ai_4 _12711_ (.A1(_04980_),
    .A2(_04981_),
    .B1(_04983_),
    .Y(_04984_));
 sky130_fd_sc_hd__and3_2 _12712_ (.A(net7939),
    .B(net2368),
    .C(net2365),
    .X(_04985_));
 sky130_fd_sc_hd__and3_1 _12713_ (.A(net7882),
    .B(net2356),
    .C(net1978),
    .X(_04986_));
 sky130_fd_sc_hd__and3_1 _12714_ (.A(net7911),
    .B(net1981),
    .C(net2359),
    .X(_04987_));
 sky130_fd_sc_hd__xor2_2 _12715_ (.A(_04986_),
    .B(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__xnor2_4 _12716_ (.A(_04985_),
    .B(_04988_),
    .Y(_04989_));
 sky130_fd_sc_hd__nand2_1 _12717_ (.A(net7853),
    .B(net1615),
    .Y(_04990_));
 sky130_fd_sc_hd__xnor2_1 _12718_ (.A(_04942_),
    .B(_04943_),
    .Y(_04991_));
 sky130_fd_sc_hd__xnor2_1 _12719_ (.A(_04990_),
    .B(_04991_),
    .Y(_04992_));
 sky130_fd_sc_hd__o21a_1 _12720_ (.A1(_04984_),
    .A2(_04989_),
    .B1(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__a21oi_4 _12721_ (.A1(_04984_),
    .A2(_04989_),
    .B1(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__or2_1 _12722_ (.A(_04986_),
    .B(_04987_),
    .X(_04995_));
 sky130_fd_sc_hd__and2_1 _12723_ (.A(_04986_),
    .B(_04987_),
    .X(_04996_));
 sky130_fd_sc_hd__a21o_2 _12724_ (.A1(_04985_),
    .A2(_04995_),
    .B1(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__nand4_1 _12725_ (.A(net1611),
    .B(_04979_),
    .C(_04994_),
    .D(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hd__a211o_1 _12726_ (.A1(net1611),
    .A2(_04979_),
    .B1(_04994_),
    .C1(_04997_),
    .X(_04999_));
 sky130_fd_sc_hd__a211o_1 _12727_ (.A1(_04994_),
    .A2(_04997_),
    .B1(net1611),
    .C1(_04979_),
    .X(_05000_));
 sky130_fd_sc_hd__and3_1 _12728_ (.A(_04998_),
    .B(_04999_),
    .C(_05000_),
    .X(_05001_));
 sky130_fd_sc_hd__xor2_1 _12729_ (.A(_04972_),
    .B(_05001_),
    .X(_05002_));
 sky130_fd_sc_hd__xor2_1 _12730_ (.A(_04984_),
    .B(_04992_),
    .X(_05003_));
 sky130_fd_sc_hd__xnor2_2 _12731_ (.A(_04989_),
    .B(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__and3_1 _12732_ (.A(net7882),
    .B(net1974),
    .C(net1971),
    .X(_05005_));
 sky130_fd_sc_hd__and3_1 _12733_ (.A(net7853),
    .B(net2338),
    .C(net1968),
    .X(_05006_));
 sky130_fd_sc_hd__a22o_1 _12734_ (.A1(net7917),
    .A2(net1350),
    .B1(_05005_),
    .B2(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__o21a_1 _12735_ (.A1(_05005_),
    .A2(_05006_),
    .B1(_05007_),
    .X(_05008_));
 sky130_fd_sc_hd__xnor2_1 _12736_ (.A(_04980_),
    .B(_04981_),
    .Y(_05009_));
 sky130_fd_sc_hd__xnor2_2 _12737_ (.A(_04982_),
    .B(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__and2_1 _12738_ (.A(net2358),
    .B(net1980),
    .X(_05011_));
 sky130_fd_sc_hd__buf_1 _12739_ (.A(_05011_),
    .X(_05012_));
 sky130_fd_sc_hd__nand2_1 _12740_ (.A(net7916),
    .B(net1342),
    .Y(_05013_));
 sky130_fd_sc_hd__and2_1 _12741_ (.A(_04904_),
    .B(net2989),
    .X(_05014_));
 sky130_fd_sc_hd__buf_1 _12742_ (.A(_05014_),
    .X(_05015_));
 sky130_fd_sc_hd__nand2_1 _12743_ (.A(net7940),
    .B(net1608),
    .Y(_05016_));
 sky130_fd_sc_hd__xnor2_1 _12744_ (.A(_05013_),
    .B(_05016_),
    .Y(_05017_));
 sky130_fd_sc_hd__a21boi_1 _12745_ (.A1(_05008_),
    .A2(_05010_),
    .B1_N(_05017_),
    .Y(_05018_));
 sky130_fd_sc_hd__o21ba_1 _12746_ (.A1(_05008_),
    .A2(_05010_),
    .B1_N(_05018_),
    .X(_05019_));
 sky130_fd_sc_hd__nand2_1 _12747_ (.A(_05004_),
    .B(net851),
    .Y(_05020_));
 sky130_fd_sc_hd__inv_2 _12748_ (.A(net7907),
    .Y(_05021_));
 sky130_fd_sc_hd__nor2_1 _12749_ (.A(net4260),
    .B(_05021_),
    .Y(_05022_));
 sky130_fd_sc_hd__and3_1 _12750_ (.A(net1608),
    .B(net1342),
    .C(net3689),
    .X(_05023_));
 sky130_fd_sc_hd__or2_1 _12751_ (.A(_05004_),
    .B(net851),
    .X(_05024_));
 sky130_fd_sc_hd__nand2_1 _12752_ (.A(net1155),
    .B(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__buf_1 _12753_ (.A(net1354),
    .X(_05026_));
 sky130_fd_sc_hd__o21ai_1 _12754_ (.A1(net1154),
    .A2(_04996_),
    .B1(_04995_),
    .Y(_05027_));
 sky130_fd_sc_hd__mux2_1 _12755_ (.A0(_04997_),
    .A1(_05027_),
    .S(net1611),
    .X(_05028_));
 sky130_fd_sc_hd__xnor2_1 _12756_ (.A(_04994_),
    .B(_05028_),
    .Y(_05029_));
 sky130_fd_sc_hd__xor2_2 _12757_ (.A(_04979_),
    .B(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__a21o_1 _12758_ (.A1(_05020_),
    .A2(_05025_),
    .B1(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__or2_1 _12759_ (.A(_05002_),
    .B(_05031_),
    .X(_05032_));
 sky130_fd_sc_hd__nand2_1 _12760_ (.A(net7850),
    .B(net1356),
    .Y(_05033_));
 sky130_fd_sc_hd__and3_2 _12761_ (.A(net7823),
    .B(_04904_),
    .C(net2989),
    .X(_05034_));
 sky130_fd_sc_hd__nand3_1 _12762_ (.A(net7337),
    .B(_04892_),
    .C(net3695),
    .Y(_05035_));
 sky130_fd_sc_hd__and3_2 _12763_ (.A(net7804),
    .B(net2354),
    .C(net2316),
    .X(_05036_));
 sky130_fd_sc_hd__xor2_1 _12764_ (.A(_05034_),
    .B(_05036_),
    .X(_05037_));
 sky130_fd_sc_hd__xnor2_2 _12765_ (.A(_05033_),
    .B(net1604),
    .Y(_05038_));
 sky130_fd_sc_hd__nand2_1 _12766_ (.A(net7784),
    .B(_04920_),
    .Y(_05039_));
 sky130_fd_sc_hd__and3_1 _12767_ (.A(net7758),
    .B(net2345),
    .C(net2342),
    .X(_05040_));
 sky130_fd_sc_hd__and3_1 _12768_ (.A(net7737),
    .B(net2978),
    .C(net2336),
    .X(_05041_));
 sky130_fd_sc_hd__xor2_1 _12769_ (.A(_05040_),
    .B(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__xnor2_2 _12770_ (.A(_05039_),
    .B(_05042_),
    .Y(_05043_));
 sky130_fd_sc_hd__o211a_1 _12771_ (.A1(_04927_),
    .A2(_04933_),
    .B1(net7800),
    .C1(net1615),
    .X(_05044_));
 sky130_fd_sc_hd__a21oi_1 _12772_ (.A1(_04927_),
    .A2(_04933_),
    .B1(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__xor2_1 _12773_ (.A(_05043_),
    .B(net1147),
    .X(_05046_));
 sky130_fd_sc_hd__xnor2_2 _12774_ (.A(_05038_),
    .B(_05046_),
    .Y(_05047_));
 sky130_fd_sc_hd__a22o_1 _12775_ (.A1(net7881),
    .A2(net1356),
    .B1(_04908_),
    .B2(_04914_),
    .X(_05048_));
 sky130_fd_sc_hd__o21ai_1 _12776_ (.A1(_04908_),
    .A2(_04914_),
    .B1(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__and3b_1 _12777_ (.A_N(net6673),
    .B(net6678),
    .C(net7275),
    .X(_05050_));
 sky130_fd_sc_hd__and3b_1 _12778_ (.A_N(net6678),
    .B(net5244),
    .C(net6673),
    .X(_05051_));
 sky130_fd_sc_hd__and3b_1 _12779_ (.A_N(net6665),
    .B(net6599),
    .C(net6748),
    .X(_05052_));
 sky130_fd_sc_hd__o21ai_1 _12780_ (.A1(_05050_),
    .A2(_05051_),
    .B1(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__nand2_1 _12781_ (.A(\svm0.vC[8] ),
    .B(_04889_),
    .Y(_05054_));
 sky130_fd_sc_hd__and2_1 _12782_ (.A(_05053_),
    .B(_05054_),
    .X(_05055_));
 sky130_fd_sc_hd__clkbuf_1 _12783_ (.A(_05055_),
    .X(_05056_));
 sky130_fd_sc_hd__buf_1 _12784_ (.A(net1958),
    .X(_05057_));
 sky130_fd_sc_hd__xnor2_1 _12785_ (.A(net7875),
    .B(net1602),
    .Y(_05058_));
 sky130_fd_sc_hd__a31oi_1 _12786_ (.A1(net7284),
    .A2(_04892_),
    .A3(_04894_),
    .B1(_05021_),
    .Y(_05059_));
 sky130_fd_sc_hd__nand2_1 _12787_ (.A(_04959_),
    .B(_05059_),
    .Y(_05060_));
 sky130_fd_sc_hd__and4_1 _12788_ (.A(net4260),
    .B(net7876),
    .C(_04974_),
    .D(_04975_),
    .X(_05061_));
 sky130_fd_sc_hd__a311oi_1 _12789_ (.A1(net7932),
    .A2(net1959),
    .A3(net1960),
    .B1(_05060_),
    .C1(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__and3_1 _12790_ (.A(net7875),
    .B(_04962_),
    .C(net2971),
    .X(_05063_));
 sky130_fd_sc_hd__buf_1 _12791_ (.A(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__o221a_1 _12792_ (.A1(net1959),
    .A2(_04965_),
    .B1(_05064_),
    .B2(net7935),
    .C1(_05060_),
    .X(_05065_));
 sky130_fd_sc_hd__o2bb2a_1 _12793_ (.A1_N(_04977_),
    .A2_N(_05058_),
    .B1(_05062_),
    .B2(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__xnor2_1 _12794_ (.A(_05049_),
    .B(net1144),
    .Y(_05067_));
 sky130_fd_sc_hd__or2_1 _12795_ (.A(_04935_),
    .B(_04939_),
    .X(_05068_));
 sky130_fd_sc_hd__a21o_1 _12796_ (.A1(_04935_),
    .A2(_04939_),
    .B1(_04916_),
    .X(_05069_));
 sky130_fd_sc_hd__nand2_1 _12797_ (.A(_05068_),
    .B(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__xnor2_1 _12798_ (.A(_05067_),
    .B(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__xnor2_2 _12799_ (.A(_05047_),
    .B(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__nand2_1 _12800_ (.A(net1343),
    .B(_04969_),
    .Y(_05073_));
 sky130_fd_sc_hd__inv_2 _12801_ (.A(_05073_),
    .Y(_05074_));
 sky130_fd_sc_hd__or2_1 _12802_ (.A(net1343),
    .B(_04969_),
    .X(_05075_));
 sky130_fd_sc_hd__a21o_1 _12803_ (.A1(_04955_),
    .A2(_05075_),
    .B1(_05074_),
    .X(_05076_));
 sky130_fd_sc_hd__nor3_1 _12804_ (.A(_04955_),
    .B(_04941_),
    .C(_05075_),
    .Y(_05077_));
 sky130_fd_sc_hd__a221o_1 _12805_ (.A1(_04955_),
    .A2(_05074_),
    .B1(_05076_),
    .B2(_04941_),
    .C1(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__xor2_2 _12806_ (.A(_05072_),
    .B(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__a21o_1 _12807_ (.A1(_04979_),
    .A2(_04997_),
    .B1(_04994_),
    .X(_05080_));
 sky130_fd_sc_hd__o21a_1 _12808_ (.A1(_04979_),
    .A2(_04997_),
    .B1(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__o31a_1 _12809_ (.A1(_04979_),
    .A2(_04994_),
    .A3(_04997_),
    .B1(net1611),
    .X(_05082_));
 sky130_fd_sc_hd__a2bb2o_1 _12810_ (.A1_N(_05081_),
    .A2_N(_05082_),
    .B1(_04998_),
    .B2(_04972_),
    .X(_05083_));
 sky130_fd_sc_hd__and2_1 _12811_ (.A(_05079_),
    .B(_05083_),
    .X(_05084_));
 sky130_fd_sc_hd__a21o_1 _12812_ (.A1(_04955_),
    .A2(net1343),
    .B1(_04941_),
    .X(_05085_));
 sky130_fd_sc_hd__a31o_1 _12813_ (.A1(_04955_),
    .A2(_04941_),
    .A3(net1343),
    .B1(_04969_),
    .X(_05086_));
 sky130_fd_sc_hd__o211ai_1 _12814_ (.A1(_04955_),
    .A2(net1343),
    .B1(_05085_),
    .C1(_05086_),
    .Y(_05087_));
 sky130_fd_sc_hd__a21oi_1 _12815_ (.A1(_05072_),
    .A2(_05087_),
    .B1(_05077_),
    .Y(_05088_));
 sky130_fd_sc_hd__nand2_1 _12816_ (.A(net7804),
    .B(net1610),
    .Y(_05089_));
 sky130_fd_sc_hd__and3_1 _12817_ (.A(net7824),
    .B(net2370),
    .C(net2367),
    .X(_05090_));
 sky130_fd_sc_hd__and3_1 _12818_ (.A(net7779),
    .B(net2354),
    .C(net2316),
    .X(_05091_));
 sky130_fd_sc_hd__xnor2_1 _12819_ (.A(_05090_),
    .B(_05091_),
    .Y(_05092_));
 sky130_fd_sc_hd__xnor2_2 _12820_ (.A(_05089_),
    .B(_05092_),
    .Y(_05093_));
 sky130_fd_sc_hd__nand2_1 _12821_ (.A(net7759),
    .B(_04919_),
    .Y(_05094_));
 sky130_fd_sc_hd__and3_1 _12822_ (.A(net7737),
    .B(net2345),
    .C(net2342),
    .X(_05095_));
 sky130_fd_sc_hd__and3_1 _12823_ (.A(net7727),
    .B(net2978),
    .C(net2336),
    .X(_05096_));
 sky130_fd_sc_hd__xnor2_1 _12824_ (.A(_05095_),
    .B(_05096_),
    .Y(_05097_));
 sky130_fd_sc_hd__xnor2_1 _12825_ (.A(_05094_),
    .B(_05097_),
    .Y(_05098_));
 sky130_fd_sc_hd__a22o_1 _12826_ (.A1(net7784),
    .A2(_04919_),
    .B1(_05040_),
    .B2(_05041_),
    .X(_05099_));
 sky130_fd_sc_hd__o21ai_2 _12827_ (.A1(_05040_),
    .A2(_05041_),
    .B1(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__xnor2_1 _12828_ (.A(net1336),
    .B(_05100_),
    .Y(_05101_));
 sky130_fd_sc_hd__xnor2_1 _12829_ (.A(_05093_),
    .B(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__nand2_1 _12830_ (.A(net7906),
    .B(net1603),
    .Y(_05103_));
 sky130_fd_sc_hd__and3_1 _12831_ (.A(net7875),
    .B(_04956_),
    .C(net2975),
    .X(_05104_));
 sky130_fd_sc_hd__and3_1 _12832_ (.A(net7848),
    .B(_04962_),
    .C(net2971),
    .X(_05105_));
 sky130_fd_sc_hd__xnor2_1 _12833_ (.A(_05104_),
    .B(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__xnor2_1 _12834_ (.A(_05103_),
    .B(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__a22oi_4 _12835_ (.A1(net7849),
    .A2(_04901_),
    .B1(_05034_),
    .B2(_05036_),
    .Y(_05108_));
 sky130_fd_sc_hd__nor2_1 _12836_ (.A(_05034_),
    .B(_05036_),
    .Y(_05109_));
 sky130_fd_sc_hd__and2_1 _12837_ (.A(net2975),
    .B(_05059_),
    .X(_05110_));
 sky130_fd_sc_hd__clkbuf_2 _12838_ (.A(net1956),
    .X(_05111_));
 sky130_fd_sc_hd__a22o_1 _12839_ (.A1(net7931),
    .A2(net1958),
    .B1(net1957),
    .B2(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__or2_1 _12840_ (.A(net1957),
    .B(_05111_),
    .X(_05113_));
 sky130_fd_sc_hd__o211ai_1 _12841_ (.A1(_05108_),
    .A2(_05109_),
    .B1(_05112_),
    .C1(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__a211o_1 _12842_ (.A1(_05112_),
    .A2(_05113_),
    .B1(_05108_),
    .C1(_05109_),
    .X(_05115_));
 sky130_fd_sc_hd__and3_1 _12843_ (.A(_05107_),
    .B(_05114_),
    .C(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__a21oi_1 _12844_ (.A1(_05114_),
    .A2(_05115_),
    .B1(_05107_),
    .Y(_05117_));
 sky130_fd_sc_hd__nor2_1 _12845_ (.A(net1006),
    .B(net1005),
    .Y(_05118_));
 sky130_fd_sc_hd__nand2_1 _12846_ (.A(_05038_),
    .B(_05043_),
    .Y(_05119_));
 sky130_fd_sc_hd__o21bai_1 _12847_ (.A1(_05038_),
    .A2(_05043_),
    .B1_N(net1147),
    .Y(_05120_));
 sky130_fd_sc_hd__nand2_1 _12848_ (.A(_05119_),
    .B(_05120_),
    .Y(_05121_));
 sky130_fd_sc_hd__xnor2_1 _12849_ (.A(_05118_),
    .B(_05121_),
    .Y(_05122_));
 sky130_fd_sc_hd__xnor2_1 _12850_ (.A(_05102_),
    .B(_05122_),
    .Y(_05123_));
 sky130_fd_sc_hd__nand3b_1 _12851_ (.A_N(_05067_),
    .B(_05068_),
    .C(_05069_),
    .Y(_05124_));
 sky130_fd_sc_hd__a21boi_1 _12852_ (.A1(_05068_),
    .A2(_05069_),
    .B1_N(_05067_),
    .Y(_05125_));
 sky130_fd_sc_hd__a21oi_2 _12853_ (.A1(_05047_),
    .A2(_05124_),
    .B1(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__and3_1 _12854_ (.A(net6749),
    .B(net6599),
    .C(net5236),
    .X(_05127_));
 sky130_fd_sc_hd__nand2_1 _12855_ (.A(net3693),
    .B(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__clkbuf_1 _12856_ (.A(net2966),
    .X(_05129_));
 sky130_fd_sc_hd__a32oi_1 _12857_ (.A1(net7272),
    .A2(_04892_),
    .A3(net3695),
    .B1(net2991),
    .B2(net7548),
    .Y(_05130_));
 sky130_fd_sc_hd__clkbuf_1 _12858_ (.A(net2305),
    .X(_05131_));
 sky130_fd_sc_hd__nand2_1 _12859_ (.A(net2310),
    .B(net1955),
    .Y(_05132_));
 sky130_fd_sc_hd__nor2_1 _12860_ (.A(net4261),
    .B(net1596),
    .Y(_05133_));
 sky130_fd_sc_hd__nand2_1 _12861_ (.A(net2334),
    .B(net2329),
    .Y(_05134_));
 sky130_fd_sc_hd__or3b_1 _12862_ (.A(net1960),
    .B(_05134_),
    .C_N(net3688),
    .X(_05135_));
 sky130_fd_sc_hd__xnor2_1 _12863_ (.A(net1957),
    .B(_05111_),
    .Y(_05136_));
 sky130_fd_sc_hd__and3_1 _12864_ (.A(net7931),
    .B(_05057_),
    .C(_05136_),
    .X(_05137_));
 sky130_fd_sc_hd__a21oi_1 _12865_ (.A1(net7931),
    .A2(_05057_),
    .B1(_05136_),
    .Y(_05138_));
 sky130_fd_sc_hd__a2bb2o_1 _12866_ (.A1_N(_05137_),
    .A2_N(_05138_),
    .B1(net1594),
    .B2(net1007),
    .X(_05139_));
 sky130_fd_sc_hd__o21ai_1 _12867_ (.A1(net1007),
    .A2(net1594),
    .B1(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__xnor2_1 _12868_ (.A(net1333),
    .B(_05140_),
    .Y(_05141_));
 sky130_fd_sc_hd__xnor2_1 _12869_ (.A(_05126_),
    .B(net791),
    .Y(_05142_));
 sky130_fd_sc_hd__xnor2_1 _12870_ (.A(net736),
    .B(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__and2_1 _12871_ (.A(_05088_),
    .B(_05143_),
    .X(_05144_));
 sky130_fd_sc_hd__nor2_1 _12872_ (.A(_05088_),
    .B(_05143_),
    .Y(_05145_));
 sky130_fd_sc_hd__or2_1 _12873_ (.A(_05144_),
    .B(_05145_),
    .X(_05146_));
 sky130_fd_sc_hd__o21a_1 _12874_ (.A1(_05032_),
    .A2(_05084_),
    .B1(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__nand2_1 _12875_ (.A(_05083_),
    .B(_05032_),
    .Y(_05148_));
 sky130_fd_sc_hd__and3b_1 _12876_ (.A_N(_05079_),
    .B(_05083_),
    .C(_05032_),
    .X(_05149_));
 sky130_fd_sc_hd__a211oi_1 _12877_ (.A1(_05079_),
    .A2(_05148_),
    .B1(_05149_),
    .C1(_05146_),
    .Y(_05150_));
 sky130_fd_sc_hd__o22a_1 _12878_ (.A1(_05079_),
    .A2(_05083_),
    .B1(_05143_),
    .B2(_05088_),
    .X(_05151_));
 sky130_fd_sc_hd__nor2_1 _12879_ (.A(_05151_),
    .B(_05144_),
    .Y(_05152_));
 sky130_fd_sc_hd__nor2_1 _12880_ (.A(net1336),
    .B(_05100_),
    .Y(_05153_));
 sky130_fd_sc_hd__a21oi_1 _12881_ (.A1(net1336),
    .A2(_05100_),
    .B1(_05093_),
    .Y(_05154_));
 sky130_fd_sc_hd__nand2_1 _12882_ (.A(net7874),
    .B(net1958),
    .Y(_05155_));
 sky130_fd_sc_hd__and3_1 _12883_ (.A(net7848),
    .B(_04956_),
    .C(net2975),
    .X(_05156_));
 sky130_fd_sc_hd__and3_1 _12884_ (.A(net7823),
    .B(_04962_),
    .C(net2971),
    .X(_05157_));
 sky130_fd_sc_hd__xnor2_1 _12885_ (.A(_05156_),
    .B(_05157_),
    .Y(_05158_));
 sky130_fd_sc_hd__xnor2_2 _12886_ (.A(_05155_),
    .B(_05158_),
    .Y(_05159_));
 sky130_fd_sc_hd__a22o_1 _12887_ (.A1(net7906),
    .A2(net1958),
    .B1(_05104_),
    .B2(_05105_),
    .X(_05160_));
 sky130_fd_sc_hd__or2_1 _12888_ (.A(_05104_),
    .B(_05105_),
    .X(_05161_));
 sky130_fd_sc_hd__a31oi_2 _12889_ (.A1(net7804),
    .A2(net1610),
    .A3(_05091_),
    .B1(_05090_),
    .Y(_05162_));
 sky130_fd_sc_hd__a21oi_2 _12890_ (.A1(net7804),
    .A2(net1610),
    .B1(_05091_),
    .Y(_05163_));
 sky130_fd_sc_hd__a211o_1 _12891_ (.A1(_05160_),
    .A2(_05161_),
    .B1(_05162_),
    .C1(_05163_),
    .X(_05164_));
 sky130_fd_sc_hd__o211ai_2 _12892_ (.A1(_05162_),
    .A2(_05163_),
    .B1(_05160_),
    .C1(_05161_),
    .Y(_05165_));
 sky130_fd_sc_hd__and3_1 _12893_ (.A(_05159_),
    .B(_05164_),
    .C(_05165_),
    .X(_05166_));
 sky130_fd_sc_hd__a21oi_2 _12894_ (.A1(_05164_),
    .A2(_05165_),
    .B1(_05159_),
    .Y(_05167_));
 sky130_fd_sc_hd__o22ai_2 _12895_ (.A1(_05153_),
    .A2(_05154_),
    .B1(_05166_),
    .B2(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__or4_2 _12896_ (.A(_05153_),
    .B(_05154_),
    .C(_05166_),
    .D(_05167_),
    .X(_05169_));
 sky130_fd_sc_hd__nand2_1 _12897_ (.A(net7737),
    .B(net1617),
    .Y(_05170_));
 sky130_fd_sc_hd__and3_1 _12898_ (.A(net7727),
    .B(net2344),
    .C(net2341),
    .X(_05171_));
 sky130_fd_sc_hd__and3_1 _12899_ (.A(net7715),
    .B(net2978),
    .C(net2335),
    .X(_05172_));
 sky130_fd_sc_hd__xor2_1 _12900_ (.A(_05171_),
    .B(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__xnor2_1 _12901_ (.A(_05170_),
    .B(_05173_),
    .Y(_05174_));
 sky130_fd_sc_hd__a22o_1 _12902_ (.A1(net7759),
    .A2(net1617),
    .B1(_05095_),
    .B2(_05096_),
    .X(_05175_));
 sky130_fd_sc_hd__o21a_1 _12903_ (.A1(_05095_),
    .A2(_05096_),
    .B1(_05175_),
    .X(_05176_));
 sky130_fd_sc_hd__nand2_1 _12904_ (.A(net7803),
    .B(_04902_),
    .Y(_05177_));
 sky130_fd_sc_hd__and3_1 _12905_ (.A(net7779),
    .B(_04905_),
    .C(_04907_),
    .X(_05178_));
 sky130_fd_sc_hd__and3_1 _12906_ (.A(net7758),
    .B(_04913_),
    .C(net2315),
    .X(_05179_));
 sky130_fd_sc_hd__xor2_1 _12907_ (.A(_05178_),
    .B(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__xnor2_2 _12908_ (.A(_05177_),
    .B(_05180_),
    .Y(_05181_));
 sky130_fd_sc_hd__xor2_1 _12909_ (.A(_05176_),
    .B(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__xnor2_1 _12910_ (.A(net1143),
    .B(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__a21o_1 _12911_ (.A1(_05168_),
    .A2(_05169_),
    .B1(net850),
    .X(_05184_));
 sky130_fd_sc_hd__nand3_1 _12912_ (.A(net850),
    .B(_05168_),
    .C(_05169_),
    .Y(_05185_));
 sky130_fd_sc_hd__and2_1 _12913_ (.A(_05184_),
    .B(_05185_),
    .X(_05186_));
 sky130_fd_sc_hd__and2_1 _12914_ (.A(net2310),
    .B(net1955),
    .X(_05187_));
 sky130_fd_sc_hd__nand2_1 _12915_ (.A(net7909),
    .B(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__nand3_1 _12916_ (.A(net7256),
    .B(_04892_),
    .C(net3695),
    .Y(_05189_));
 sky130_fd_sc_hd__a32oi_1 _12917_ (.A1(net5232),
    .A2(_04856_),
    .A3(_04897_),
    .B1(_04889_),
    .B2(\svm0.vC[10] ),
    .Y(_05190_));
 sky130_fd_sc_hd__and2_1 _12918_ (.A(net2304),
    .B(net2964),
    .X(_05191_));
 sky130_fd_sc_hd__nand2_1 _12919_ (.A(net7933),
    .B(net1949),
    .Y(_05192_));
 sky130_fd_sc_hd__xnor2_1 _12920_ (.A(_05188_),
    .B(_05192_),
    .Y(_05193_));
 sky130_fd_sc_hd__a22oi_1 _12921_ (.A1(net7931),
    .A2(net1958),
    .B1(net1957),
    .B2(_05111_),
    .Y(_05194_));
 sky130_fd_sc_hd__nor2_1 _12922_ (.A(net1957),
    .B(_05111_),
    .Y(_05195_));
 sky130_fd_sc_hd__or4_1 _12923_ (.A(_05194_),
    .B(_05195_),
    .C(_05108_),
    .D(_05109_),
    .X(_05196_));
 sky130_fd_sc_hd__o22a_1 _12924_ (.A1(_05194_),
    .A2(_05195_),
    .B1(_05108_),
    .B2(_05109_),
    .X(_05197_));
 sky130_fd_sc_hd__a21o_1 _12925_ (.A1(_05196_),
    .A2(_05107_),
    .B1(_05197_),
    .X(_05198_));
 sky130_fd_sc_hd__xnor2_2 _12926_ (.A(net1140),
    .B(net1004),
    .Y(_05199_));
 sky130_fd_sc_hd__a211o_1 _12927_ (.A1(_05119_),
    .A2(_05120_),
    .B1(net1006),
    .C1(net1005),
    .X(_05200_));
 sky130_fd_sc_hd__o211a_1 _12928_ (.A1(net1006),
    .A2(net1005),
    .B1(_05119_),
    .C1(_05120_),
    .X(_05201_));
 sky130_fd_sc_hd__a21oi_2 _12929_ (.A1(_05102_),
    .A2(_05200_),
    .B1(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__xnor2_2 _12930_ (.A(_05199_),
    .B(_05202_),
    .Y(_05203_));
 sky130_fd_sc_hd__xnor2_2 _12931_ (.A(_05186_),
    .B(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__nand2_1 _12932_ (.A(net1333),
    .B(_05140_),
    .Y(_05205_));
 sky130_fd_sc_hd__or2_1 _12933_ (.A(_05126_),
    .B(net791),
    .X(_05206_));
 sky130_fd_sc_hd__and2_1 _12934_ (.A(_05126_),
    .B(net791),
    .X(_05207_));
 sky130_fd_sc_hd__a21o_1 _12935_ (.A1(_05206_),
    .A2(net736),
    .B1(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__xnor2_1 _12936_ (.A(net790),
    .B(_05208_),
    .Y(_05209_));
 sky130_fd_sc_hd__xor2_1 _12937_ (.A(_05204_),
    .B(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__xnor2_1 _12938_ (.A(_05152_),
    .B(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__nand2_1 _12939_ (.A(net7917),
    .B(net1350),
    .Y(_05212_));
 sky130_fd_sc_hd__xor2_1 _12940_ (.A(_05005_),
    .B(_05006_),
    .X(_05213_));
 sky130_fd_sc_hd__xnor2_2 _12941_ (.A(_05212_),
    .B(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__and3_1 _12942_ (.A(net7939),
    .B(net2356),
    .C(net1978),
    .X(_05215_));
 sky130_fd_sc_hd__and2_1 _12943_ (.A(net1974),
    .B(net1971),
    .X(_05216_));
 sky130_fd_sc_hd__and2_1 _12944_ (.A(net2338),
    .B(net1968),
    .X(_05217_));
 sky130_fd_sc_hd__and4_1 _12945_ (.A(net7916),
    .B(net7883),
    .C(_05216_),
    .D(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__a41o_1 _12946_ (.A1(net7940),
    .A2(net7889),
    .A3(net1350),
    .A4(_05217_),
    .B1(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__a41o_1 _12947_ (.A1(net7940),
    .A2(net7917),
    .A3(net1350),
    .A4(_05216_),
    .B1(_05219_),
    .X(_05220_));
 sky130_fd_sc_hd__o21ai_1 _12948_ (.A1(_05214_),
    .A2(net1593),
    .B1(net1003),
    .Y(_05221_));
 sky130_fd_sc_hd__nand2_1 _12949_ (.A(_05214_),
    .B(net1593),
    .Y(_05222_));
 sky130_fd_sc_hd__xnor2_1 _12950_ (.A(_05008_),
    .B(_05017_),
    .Y(_05223_));
 sky130_fd_sc_hd__xnor2_1 _12951_ (.A(_05010_),
    .B(_05223_),
    .Y(_05224_));
 sky130_fd_sc_hd__a21oi_1 _12952_ (.A1(_05221_),
    .A2(_05222_),
    .B1(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__xnor2_1 _12953_ (.A(net789),
    .B(_05031_),
    .Y(_05226_));
 sky130_fd_sc_hd__nand2_1 _12954_ (.A(_05002_),
    .B(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__or2_1 _12955_ (.A(_05002_),
    .B(_05226_),
    .X(_05228_));
 sky130_fd_sc_hd__nor2_1 _12956_ (.A(net7889),
    .B(net1350),
    .Y(_05229_));
 sky130_fd_sc_hd__o2111a_1 _12957_ (.A1(_04982_),
    .A2(_05229_),
    .B1(_05216_),
    .C1(_05217_),
    .D1(net3689),
    .X(_05230_));
 sky130_fd_sc_hd__xor2_1 _12958_ (.A(_05214_),
    .B(net1593),
    .X(_05231_));
 sky130_fd_sc_hd__o21ai_1 _12959_ (.A1(net1003),
    .A2(_05231_),
    .B1(_05221_),
    .Y(_05232_));
 sky130_fd_sc_hd__nor2_1 _12960_ (.A(_05224_),
    .B(_05232_),
    .Y(_05233_));
 sky130_fd_sc_hd__a41o_1 _12961_ (.A1(_05224_),
    .A2(net1003),
    .A3(_05214_),
    .A4(net1593),
    .B1(_05233_),
    .X(_05234_));
 sky130_fd_sc_hd__nand2_1 _12962_ (.A(net1002),
    .B(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__xnor2_1 _12963_ (.A(_05004_),
    .B(net851),
    .Y(_05236_));
 sky130_fd_sc_hd__or2_1 _12964_ (.A(_05030_),
    .B(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__mux2_1 _12965_ (.A0(_05024_),
    .A1(_05020_),
    .S(_05030_),
    .X(_05238_));
 sky130_fd_sc_hd__mux2_1 _12966_ (.A0(_05237_),
    .A1(_05238_),
    .S(net1155),
    .X(_05239_));
 sky130_fd_sc_hd__a211o_1 _12967_ (.A1(_05227_),
    .A2(_05228_),
    .B1(_05235_),
    .C1(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__nor2_1 _12968_ (.A(net1140),
    .B(net1004),
    .Y(_05241_));
 sky130_fd_sc_hd__xor2_1 _12969_ (.A(net1140),
    .B(net1004),
    .X(_05242_));
 sky130_fd_sc_hd__a211oi_1 _12970_ (.A1(_05168_),
    .A2(_05169_),
    .B1(net850),
    .C1(_05242_),
    .Y(_05243_));
 sky130_fd_sc_hd__and4_1 _12971_ (.A(net850),
    .B(_05199_),
    .C(_05168_),
    .D(_05169_),
    .X(_05244_));
 sky130_fd_sc_hd__nor3b_1 _12972_ (.A(_05243_),
    .B(_05244_),
    .C_N(_05202_),
    .Y(_05245_));
 sky130_fd_sc_hd__nand2_1 _12973_ (.A(_05241_),
    .B(net735),
    .Y(_05246_));
 sky130_fd_sc_hd__and3_1 _12974_ (.A(_05242_),
    .B(_05184_),
    .C(_05185_),
    .X(_05247_));
 sky130_fd_sc_hd__or3_1 _12975_ (.A(_05241_),
    .B(_05247_),
    .C(net735),
    .X(_05248_));
 sky130_fd_sc_hd__nand2_1 _12976_ (.A(net7785),
    .B(net1355),
    .Y(_05249_));
 sky130_fd_sc_hd__and3_1 _12977_ (.A(net7759),
    .B(net1986),
    .C(net2364),
    .X(_05250_));
 sky130_fd_sc_hd__nand2_1 _12978_ (.A(net7748),
    .B(_05012_),
    .Y(_05251_));
 sky130_fd_sc_hd__xor2_1 _12979_ (.A(_05250_),
    .B(_05251_),
    .X(_05252_));
 sky130_fd_sc_hd__xnor2_2 _12980_ (.A(_05249_),
    .B(_05252_),
    .Y(_05253_));
 sky130_fd_sc_hd__o211a_1 _12981_ (.A1(_05171_),
    .A2(_05172_),
    .B1(net7738),
    .C1(net1617),
    .X(_05254_));
 sky130_fd_sc_hd__a21o_1 _12982_ (.A1(_05171_),
    .A2(_05172_),
    .B1(_05254_),
    .X(_05255_));
 sky130_fd_sc_hd__nand2_1 _12983_ (.A(net7728),
    .B(net1616),
    .Y(_05256_));
 sky130_fd_sc_hd__and3_1 _12984_ (.A(net7688),
    .B(net2977),
    .C(net2335),
    .X(_05257_));
 sky130_fd_sc_hd__and3_1 _12985_ (.A(net7715),
    .B(net2344),
    .C(net2341),
    .X(_05258_));
 sky130_fd_sc_hd__xor2_1 _12986_ (.A(_05257_),
    .B(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__xnor2_2 _12987_ (.A(_05256_),
    .B(_05259_),
    .Y(_05260_));
 sky130_fd_sc_hd__xnor2_1 _12988_ (.A(_05255_),
    .B(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__xnor2_2 _12989_ (.A(_05253_),
    .B(_05261_),
    .Y(_05262_));
 sky130_fd_sc_hd__a21o_1 _12990_ (.A1(_05176_),
    .A2(_05181_),
    .B1(net1143),
    .X(_05263_));
 sky130_fd_sc_hd__o21a_1 _12991_ (.A1(_05176_),
    .A2(_05181_),
    .B1(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__nand2_1 _12992_ (.A(net7847),
    .B(net1602),
    .Y(_05265_));
 sky130_fd_sc_hd__and3_1 _12993_ (.A(net7802),
    .B(net2324),
    .C(net2320),
    .X(_05266_));
 sky130_fd_sc_hd__and3_1 _12994_ (.A(net7822),
    .B(_04957_),
    .C(_04959_),
    .X(_05267_));
 sky130_fd_sc_hd__xor2_1 _12995_ (.A(_05266_),
    .B(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__xnor2_2 _12996_ (.A(_05265_),
    .B(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__a22o_1 _12997_ (.A1(net7803),
    .A2(net1619),
    .B1(_05178_),
    .B2(_05179_),
    .X(_05270_));
 sky130_fd_sc_hd__or2_1 _12998_ (.A(_05178_),
    .B(_05179_),
    .X(_05271_));
 sky130_fd_sc_hd__and2_1 _12999_ (.A(_05156_),
    .B(_05157_),
    .X(_05272_));
 sky130_fd_sc_hd__o211a_1 _13000_ (.A1(_05156_),
    .A2(_05157_),
    .B1(net7874),
    .C1(net1959),
    .X(_05273_));
 sky130_fd_sc_hd__a211oi_1 _13001_ (.A1(_05270_),
    .A2(_05271_),
    .B1(_05272_),
    .C1(_05273_),
    .Y(_05274_));
 sky130_fd_sc_hd__o211a_1 _13002_ (.A1(_05272_),
    .A2(_05273_),
    .B1(_05270_),
    .C1(_05271_),
    .X(_05275_));
 sky130_fd_sc_hd__nor2_1 _13003_ (.A(_05274_),
    .B(_05275_),
    .Y(_05276_));
 sky130_fd_sc_hd__xnor2_2 _13004_ (.A(_05269_),
    .B(_05276_),
    .Y(_05277_));
 sky130_fd_sc_hd__xnor2_1 _13005_ (.A(_05264_),
    .B(_05277_),
    .Y(_05278_));
 sky130_fd_sc_hd__xnor2_1 _13006_ (.A(_05262_),
    .B(_05278_),
    .Y(_05279_));
 sky130_fd_sc_hd__nor2_1 _13007_ (.A(_05153_),
    .B(_05154_),
    .Y(_05280_));
 sky130_fd_sc_hd__or2_1 _13008_ (.A(net1336),
    .B(_05100_),
    .X(_05281_));
 sky130_fd_sc_hd__a21o_1 _13009_ (.A1(net1336),
    .A2(_05100_),
    .B1(_05093_),
    .X(_05282_));
 sky130_fd_sc_hd__o211a_1 _13010_ (.A1(_05166_),
    .A2(_05167_),
    .B1(_05281_),
    .C1(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__o32a_1 _13011_ (.A1(_05280_),
    .A2(_05166_),
    .A3(_05167_),
    .B1(net850),
    .B2(_05283_),
    .X(_05284_));
 sky130_fd_sc_hd__clkbuf_2 _13012_ (.A(net3693),
    .X(_05285_));
 sky130_fd_sc_hd__a32o_1 _13013_ (.A1(net7246),
    .A2(_04892_),
    .A3(_04894_),
    .B1(net2991),
    .B2(net7546),
    .X(_05286_));
 sky130_fd_sc_hd__a31oi_4 _13014_ (.A1(net5215),
    .A2(net3029),
    .A3(_05285_),
    .B1(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__xnor2_1 _13015_ (.A(net7878),
    .B(_05287_),
    .Y(_05288_));
 sky130_fd_sc_hd__and3_1 _13016_ (.A(net7908),
    .B(_05189_),
    .C(net2965),
    .X(_05289_));
 sky130_fd_sc_hd__clkbuf_2 _13017_ (.A(_05289_),
    .X(_05290_));
 sky130_fd_sc_hd__and3_1 _13018_ (.A(net4259),
    .B(net7878),
    .C(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__a211o_1 _13019_ (.A1(net7933),
    .A2(_05288_),
    .B1(_05291_),
    .C1(net1596),
    .X(_05292_));
 sky130_fd_sc_hd__clkbuf_1 _13020_ (.A(net1948),
    .X(_05293_));
 sky130_fd_sc_hd__buf_1 _13021_ (.A(_05187_),
    .X(_05294_));
 sky130_fd_sc_hd__a31o_1 _13022_ (.A1(net7933),
    .A2(_05290_),
    .A3(net1592),
    .B1(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__and3_1 _13023_ (.A(net7878),
    .B(net2966),
    .C(net2305),
    .X(_05296_));
 sky130_fd_sc_hd__o22a_1 _13024_ (.A1(net7933),
    .A2(_05296_),
    .B1(net1592),
    .B2(_05294_),
    .X(_05297_));
 sky130_fd_sc_hd__nor2_1 _13025_ (.A(_05290_),
    .B(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__a21oi_1 _13026_ (.A1(_05292_),
    .A2(_05295_),
    .B1(_05298_),
    .Y(_05299_));
 sky130_fd_sc_hd__nand2_1 _13027_ (.A(_05160_),
    .B(_05161_),
    .Y(_05300_));
 sky130_fd_sc_hd__a211o_1 _13028_ (.A1(_05159_),
    .A2(_05300_),
    .B1(_05162_),
    .C1(_05163_),
    .X(_05301_));
 sky130_fd_sc_hd__o21ai_2 _13029_ (.A1(_05159_),
    .A2(_05300_),
    .B1(_05301_),
    .Y(_05302_));
 sky130_fd_sc_hd__xnor2_2 _13030_ (.A(net920),
    .B(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__xor2_1 _13031_ (.A(_05284_),
    .B(_05303_),
    .X(_05304_));
 sky130_fd_sc_hd__xnor2_1 _13032_ (.A(_05279_),
    .B(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__a21o_1 _13033_ (.A1(_05246_),
    .A2(_05248_),
    .B1(net684),
    .X(_05306_));
 sky130_fd_sc_hd__or2_1 _13034_ (.A(net1140),
    .B(net1004),
    .X(_05307_));
 sky130_fd_sc_hd__o21ai_1 _13035_ (.A1(_05247_),
    .A2(net735),
    .B1(_05307_),
    .Y(_05308_));
 sky130_fd_sc_hd__or2_1 _13036_ (.A(_05307_),
    .B(net735),
    .X(_05309_));
 sky130_fd_sc_hd__a21bo_1 _13037_ (.A1(_05308_),
    .A2(_05309_),
    .B1_N(net684),
    .X(_05310_));
 sky130_fd_sc_hd__or2_1 _13038_ (.A(net791),
    .B(net736),
    .X(_05311_));
 sky130_fd_sc_hd__a21o_1 _13039_ (.A1(net791),
    .A2(net736),
    .B1(_05126_),
    .X(_05312_));
 sky130_fd_sc_hd__nand3b_1 _13040_ (.A_N(net790),
    .B(_05185_),
    .C(_05184_),
    .Y(_05313_));
 sky130_fd_sc_hd__a21o_1 _13041_ (.A1(_05184_),
    .A2(_05185_),
    .B1(net790),
    .X(_05314_));
 sky130_fd_sc_hd__mux2_1 _13042_ (.A0(_05313_),
    .A1(_05314_),
    .S(_05203_),
    .X(_05315_));
 sky130_fd_sc_hd__a32o_1 _13043_ (.A1(_05311_),
    .A2(_05312_),
    .A3(_05315_),
    .B1(net790),
    .B2(_05204_),
    .X(_05316_));
 sky130_fd_sc_hd__a21o_1 _13044_ (.A1(_05306_),
    .A2(_05310_),
    .B1(_05316_),
    .X(_05317_));
 sky130_fd_sc_hd__and2_1 _13045_ (.A(_05306_),
    .B(_05310_),
    .X(_05318_));
 sky130_fd_sc_hd__nand2_1 _13046_ (.A(_05318_),
    .B(_05316_),
    .Y(_05319_));
 sky130_fd_sc_hd__or4bb_1 _13047_ (.A(_05211_),
    .B(net535),
    .C_N(_05317_),
    .D_N(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__nor2_1 _13048_ (.A(net789),
    .B(_05004_),
    .Y(_05321_));
 sky130_fd_sc_hd__nand2_1 _13049_ (.A(net789),
    .B(_05004_),
    .Y(_05322_));
 sky130_fd_sc_hd__inv_2 _13050_ (.A(net851),
    .Y(_05323_));
 sky130_fd_sc_hd__a21o_1 _13051_ (.A1(_05030_),
    .A2(_05322_),
    .B1(_05323_),
    .X(_05324_));
 sky130_fd_sc_hd__o21ai_1 _13052_ (.A1(_05030_),
    .A2(_05321_),
    .B1(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__o21a_1 _13053_ (.A1(_05323_),
    .A2(_05321_),
    .B1(_05322_),
    .X(_05326_));
 sky130_fd_sc_hd__o2bb2a_1 _13054_ (.A1_N(_05325_),
    .A2_N(net1155),
    .B1(_05326_),
    .B2(_05030_),
    .X(_05327_));
 sky130_fd_sc_hd__or3_1 _13055_ (.A(_05079_),
    .B(_05327_),
    .C(_05002_),
    .X(_05328_));
 sky130_fd_sc_hd__nand2_1 _13056_ (.A(net790),
    .B(_05208_),
    .Y(_05329_));
 sky130_fd_sc_hd__mux2_1 _13057_ (.A0(_05329_),
    .A1(_05209_),
    .S(_05204_),
    .X(_05330_));
 sky130_fd_sc_hd__or3_1 _13058_ (.A(_05204_),
    .B(net790),
    .C(_05208_),
    .X(_05331_));
 sky130_fd_sc_hd__mux2_1 _13059_ (.A0(_05330_),
    .A1(_05331_),
    .S(_05318_),
    .X(_05332_));
 sky130_fd_sc_hd__a211o_1 _13060_ (.A1(_05151_),
    .A2(_05328_),
    .B1(_05144_),
    .C1(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__o31a_1 _13061_ (.A1(_05147_),
    .A2(_05150_),
    .A3(_05320_),
    .B1(_05333_),
    .X(_05334_));
 sky130_fd_sc_hd__nand2_1 _13062_ (.A(_05284_),
    .B(_05303_),
    .Y(_05335_));
 sky130_fd_sc_hd__nor2_1 _13063_ (.A(_05284_),
    .B(_05303_),
    .Y(_05336_));
 sky130_fd_sc_hd__a21oi_1 _13064_ (.A1(_05279_),
    .A2(_05335_),
    .B1(_05336_),
    .Y(_05337_));
 sky130_fd_sc_hd__and3_1 _13065_ (.A(net7846),
    .B(net2966),
    .C(net2305),
    .X(_05338_));
 sky130_fd_sc_hd__nand2_1 _13066_ (.A(net7908),
    .B(net1948),
    .Y(_05339_));
 sky130_fd_sc_hd__nand2_1 _13067_ (.A(net7877),
    .B(_05191_),
    .Y(_05340_));
 sky130_fd_sc_hd__xnor2_1 _13068_ (.A(_05339_),
    .B(_05340_),
    .Y(_05341_));
 sky130_fd_sc_hd__xnor2_2 _13069_ (.A(_05338_),
    .B(_05341_),
    .Y(_05342_));
 sky130_fd_sc_hd__and3b_1 _13070_ (.A_N(net6673),
    .B(net6677),
    .C(net7232),
    .X(_05343_));
 sky130_fd_sc_hd__and3b_1 _13071_ (.A_N(net6677),
    .B(net5204),
    .C(net6673),
    .X(_05344_));
 sky130_fd_sc_hd__o21ai_1 _13072_ (.A1(_05343_),
    .A2(_05344_),
    .B1(_05052_),
    .Y(_05345_));
 sky130_fd_sc_hd__buf_1 _13073_ (.A(_05345_),
    .X(_05346_));
 sky130_fd_sc_hd__nand4b_1 _13074_ (.A_N(net6664),
    .B(net6673),
    .C(net6677),
    .D(\svm0.vC[12] ),
    .Y(_05347_));
 sky130_fd_sc_hd__and2_1 _13075_ (.A(_05346_),
    .B(net4255),
    .X(_05348_));
 sky130_fd_sc_hd__nand2_1 _13076_ (.A(_05290_),
    .B(_05296_),
    .Y(_05349_));
 sky130_fd_sc_hd__o21ai_1 _13077_ (.A1(_05290_),
    .A2(_05296_),
    .B1(_05287_),
    .Y(_05350_));
 sky130_fd_sc_hd__nand2_1 _13078_ (.A(_05345_),
    .B(net4255),
    .Y(_05351_));
 sky130_fd_sc_hd__o221a_1 _13079_ (.A1(_05290_),
    .A2(_05296_),
    .B1(_05351_),
    .B2(net4259),
    .C1(_05287_),
    .X(_05352_));
 sky130_fd_sc_hd__a31o_1 _13080_ (.A1(net2303),
    .A2(_05349_),
    .A3(_05350_),
    .B1(_05352_),
    .X(_05353_));
 sky130_fd_sc_hd__nor2_1 _13081_ (.A(net4259),
    .B(_05351_),
    .Y(_05354_));
 sky130_fd_sc_hd__o2bb2a_1 _13082_ (.A1_N(net7933),
    .A2_N(_05353_),
    .B1(_05349_),
    .B2(_05354_),
    .X(_05355_));
 sky130_fd_sc_hd__xnor2_1 _13083_ (.A(_05342_),
    .B(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__and4_1 _13084_ (.A(_05294_),
    .B(net1949),
    .C(_05288_),
    .D(net3688),
    .X(_05357_));
 sky130_fd_sc_hd__a211o_1 _13085_ (.A1(_05270_),
    .A2(_05271_),
    .B1(_05272_),
    .C1(_05273_),
    .X(_05358_));
 sky130_fd_sc_hd__a21oi_1 _13086_ (.A1(_05269_),
    .A2(_05358_),
    .B1(_05275_),
    .Y(_05359_));
 sky130_fd_sc_hd__xnor2_1 _13087_ (.A(_05357_),
    .B(net1001),
    .Y(_05360_));
 sky130_fd_sc_hd__xor2_1 _13088_ (.A(net919),
    .B(_05360_),
    .X(_05361_));
 sky130_fd_sc_hd__or2_1 _13089_ (.A(_05262_),
    .B(_05277_),
    .X(_05362_));
 sky130_fd_sc_hd__a21bo_1 _13090_ (.A1(_05262_),
    .A2(_05277_),
    .B1_N(_05264_),
    .X(_05363_));
 sky130_fd_sc_hd__nand3_1 _13091_ (.A(_05361_),
    .B(_05362_),
    .C(_05363_),
    .Y(_05364_));
 sky130_fd_sc_hd__a21o_1 _13092_ (.A1(_05362_),
    .A2(_05363_),
    .B1(_05361_),
    .X(_05365_));
 sky130_fd_sc_hd__and3_1 _13093_ (.A(net7688),
    .B(net1973),
    .C(net1970),
    .X(_05366_));
 sky130_fd_sc_hd__and3_1 _13094_ (.A(net7672),
    .B(net2339),
    .C(net1967),
    .X(_05367_));
 sky130_fd_sc_hd__and3_1 _13095_ (.A(net7716),
    .B(net2351),
    .C(net2347),
    .X(_05368_));
 sky130_fd_sc_hd__xnor2_1 _13096_ (.A(_05367_),
    .B(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__xnor2_1 _13097_ (.A(_05366_),
    .B(_05369_),
    .Y(_05370_));
 sky130_fd_sc_hd__a22o_1 _13098_ (.A1(net7728),
    .A2(net1616),
    .B1(_05257_),
    .B2(_05258_),
    .X(_05371_));
 sky130_fd_sc_hd__o21a_1 _13099_ (.A1(_05257_),
    .A2(_05258_),
    .B1(_05371_),
    .X(_05372_));
 sky130_fd_sc_hd__nand2_1 _13100_ (.A(net7757),
    .B(net1620),
    .Y(_05373_));
 sky130_fd_sc_hd__and3_1 _13101_ (.A(net7725),
    .B(net2355),
    .C(_05035_),
    .X(_05374_));
 sky130_fd_sc_hd__and3_1 _13102_ (.A(net7735),
    .B(_04904_),
    .C(net2989),
    .X(_05375_));
 sky130_fd_sc_hd__xor2_1 _13103_ (.A(_05374_),
    .B(_05375_),
    .X(_05376_));
 sky130_fd_sc_hd__xnor2_1 _13104_ (.A(_05373_),
    .B(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__xor2_1 _13105_ (.A(_05372_),
    .B(net1138),
    .X(_05378_));
 sky130_fd_sc_hd__xnor2_1 _13106_ (.A(_05370_),
    .B(_05378_),
    .Y(_05379_));
 sky130_fd_sc_hd__nand2_1 _13107_ (.A(_05255_),
    .B(_05260_),
    .Y(_05380_));
 sky130_fd_sc_hd__nor2_1 _13108_ (.A(_05255_),
    .B(_05260_),
    .Y(_05381_));
 sky130_fd_sc_hd__a21o_1 _13109_ (.A1(_05253_),
    .A2(_05380_),
    .B1(_05381_),
    .X(_05382_));
 sky130_fd_sc_hd__and3_1 _13110_ (.A(net7778),
    .B(net2973),
    .C(net2971),
    .X(_05383_));
 sky130_fd_sc_hd__and3_1 _13111_ (.A(net7822),
    .B(_05053_),
    .C(_05054_),
    .X(_05384_));
 sky130_fd_sc_hd__and3_1 _13112_ (.A(net7801),
    .B(net2976),
    .C(net2974),
    .X(_05385_));
 sky130_fd_sc_hd__xor2_1 _13113_ (.A(_05384_),
    .B(_05385_),
    .X(_05386_));
 sky130_fd_sc_hd__xnor2_1 _13114_ (.A(_05383_),
    .B(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__nand2_1 _13115_ (.A(_05266_),
    .B(_05267_),
    .Y(_05388_));
 sky130_fd_sc_hd__o211ai_2 _13116_ (.A1(_05266_),
    .A2(_05267_),
    .B1(net7847),
    .C1(net1601),
    .Y(_05389_));
 sky130_fd_sc_hd__nand2_1 _13117_ (.A(_05388_),
    .B(_05389_),
    .Y(_05390_));
 sky130_fd_sc_hd__a32oi_2 _13118_ (.A1(net7736),
    .A2(_05011_),
    .A3(_05250_),
    .B1(net1619),
    .B2(net7783),
    .Y(_05391_));
 sky130_fd_sc_hd__a21oi_1 _13119_ (.A1(net7736),
    .A2(_05012_),
    .B1(_05250_),
    .Y(_05392_));
 sky130_fd_sc_hd__or2_1 _13120_ (.A(_05391_),
    .B(_05392_),
    .X(_05393_));
 sky130_fd_sc_hd__xor2_1 _13121_ (.A(_05390_),
    .B(_05393_),
    .X(_05394_));
 sky130_fd_sc_hd__xnor2_1 _13122_ (.A(net1585),
    .B(_05394_),
    .Y(_05395_));
 sky130_fd_sc_hd__xnor2_1 _13123_ (.A(_05382_),
    .B(net849),
    .Y(_05396_));
 sky130_fd_sc_hd__xnor2_1 _13124_ (.A(_05379_),
    .B(_05396_),
    .Y(_05397_));
 sky130_fd_sc_hd__a21oi_1 _13125_ (.A1(_05364_),
    .A2(_05365_),
    .B1(net734),
    .Y(_05398_));
 sky130_fd_sc_hd__and3_1 _13126_ (.A(net734),
    .B(_05364_),
    .C(_05365_),
    .X(_05399_));
 sky130_fd_sc_hd__or2_1 _13127_ (.A(_05398_),
    .B(_05399_),
    .X(_05400_));
 sky130_fd_sc_hd__clkbuf_2 _13128_ (.A(_05400_),
    .X(_05401_));
 sky130_fd_sc_hd__nand2_1 _13129_ (.A(net920),
    .B(_05302_),
    .Y(_05402_));
 sky130_fd_sc_hd__or3_1 _13130_ (.A(_05398_),
    .B(_05399_),
    .C(net848),
    .X(_05403_));
 sky130_fd_sc_hd__or2_1 _13131_ (.A(net683),
    .B(net848),
    .X(_05404_));
 sky130_fd_sc_hd__o211ai_2 _13132_ (.A1(net683),
    .A2(_05401_),
    .B1(_05403_),
    .C1(_05404_),
    .Y(_05405_));
 sky130_fd_sc_hd__nand2_1 _13133_ (.A(_05349_),
    .B(_05350_),
    .Y(_05406_));
 sky130_fd_sc_hd__a21o_1 _13134_ (.A1(_05342_),
    .A2(net2303),
    .B1(_05406_),
    .X(_05407_));
 sky130_fd_sc_hd__a31o_1 _13135_ (.A1(_05290_),
    .A2(_05296_),
    .A3(_05342_),
    .B1(net7936),
    .X(_05408_));
 sky130_fd_sc_hd__o211ai_1 _13136_ (.A1(_05342_),
    .A2(net2303),
    .B1(_05407_),
    .C1(_05408_),
    .Y(_05409_));
 sky130_fd_sc_hd__a211o_1 _13137_ (.A1(_05388_),
    .A2(_05389_),
    .B1(_05391_),
    .C1(_05392_),
    .X(_05410_));
 sky130_fd_sc_hd__a32o_1 _13138_ (.A1(_05388_),
    .A2(_05389_),
    .A3(_05393_),
    .B1(_05410_),
    .B2(net1585),
    .X(_05411_));
 sky130_fd_sc_hd__nand2_1 _13139_ (.A(net7873),
    .B(net1947),
    .Y(_05412_));
 sky130_fd_sc_hd__and3_1 _13140_ (.A(net7821),
    .B(net2966),
    .C(net2305),
    .X(_05413_));
 sky130_fd_sc_hd__and3_1 _13141_ (.A(net7845),
    .B(net2304),
    .C(net2964),
    .X(_05414_));
 sky130_fd_sc_hd__xnor2_1 _13142_ (.A(_05413_),
    .B(_05414_),
    .Y(_05415_));
 sky130_fd_sc_hd__xnor2_1 _13143_ (.A(_05412_),
    .B(_05415_),
    .Y(_05416_));
 sky130_fd_sc_hd__a32o_1 _13144_ (.A1(net7877),
    .A2(net1949),
    .A3(_05338_),
    .B1(net1947),
    .B2(net7909),
    .X(_05417_));
 sky130_fd_sc_hd__a21o_1 _13145_ (.A1(net7877),
    .A2(net1949),
    .B1(_05338_),
    .X(_05418_));
 sky130_fd_sc_hd__and3_1 _13146_ (.A(net7215),
    .B(net3029),
    .C(_04894_),
    .X(_05419_));
 sky130_fd_sc_hd__a32o_1 _13147_ (.A1(net5199),
    .A2(net3028),
    .A3(net3693),
    .B1(net2992),
    .B2(\svm0.vC[13] ),
    .X(_05420_));
 sky130_fd_sc_hd__or3_1 _13148_ (.A(net4261),
    .B(net2302),
    .C(net2298),
    .X(_05421_));
 sky130_fd_sc_hd__and3_1 _13149_ (.A(net7909),
    .B(net2956),
    .C(net4254),
    .X(_05422_));
 sky130_fd_sc_hd__xnor2_1 _13150_ (.A(_05421_),
    .B(_05422_),
    .Y(_05423_));
 sky130_fd_sc_hd__nand3_1 _13151_ (.A(_05417_),
    .B(_05418_),
    .C(_05423_),
    .Y(_05424_));
 sky130_fd_sc_hd__a21o_1 _13152_ (.A1(_05417_),
    .A2(_05418_),
    .B1(_05423_),
    .X(_05425_));
 sky130_fd_sc_hd__nand3_1 _13153_ (.A(_05416_),
    .B(_05424_),
    .C(_05425_),
    .Y(_05426_));
 sky130_fd_sc_hd__a21o_1 _13154_ (.A1(_05424_),
    .A2(_05425_),
    .B1(_05416_),
    .X(_05427_));
 sky130_fd_sc_hd__and3_1 _13155_ (.A(net917),
    .B(_05426_),
    .C(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__a21o_1 _13156_ (.A1(_05426_),
    .A2(_05427_),
    .B1(net917),
    .X(_05429_));
 sky130_fd_sc_hd__and2b_1 _13157_ (.A_N(_05428_),
    .B(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__xnor2_1 _13158_ (.A(net918),
    .B(_05430_),
    .Y(_05431_));
 sky130_fd_sc_hd__nor2_1 _13159_ (.A(_05372_),
    .B(net1138),
    .Y(_05432_));
 sky130_fd_sc_hd__a21oi_1 _13160_ (.A1(_05372_),
    .A2(net1138),
    .B1(_05370_),
    .Y(_05433_));
 sky130_fd_sc_hd__a21o_1 _13161_ (.A1(_05383_),
    .A2(_05385_),
    .B1(_05384_),
    .X(_05434_));
 sky130_fd_sc_hd__or2_1 _13162_ (.A(_05383_),
    .B(_05385_),
    .X(_05435_));
 sky130_fd_sc_hd__and2_1 _13163_ (.A(_05374_),
    .B(_05375_),
    .X(_05436_));
 sky130_fd_sc_hd__o211a_1 _13164_ (.A1(_05374_),
    .A2(_05375_),
    .B1(net7757),
    .C1(net1620),
    .X(_05437_));
 sky130_fd_sc_hd__a211o_1 _13165_ (.A1(_05434_),
    .A2(_05435_),
    .B1(_05436_),
    .C1(_05437_),
    .X(_05438_));
 sky130_fd_sc_hd__o211ai_1 _13166_ (.A1(_05436_),
    .A2(_05437_),
    .B1(_05434_),
    .C1(_05435_),
    .Y(_05439_));
 sky130_fd_sc_hd__and3_1 _13167_ (.A(net7756),
    .B(net2324),
    .C(net2320),
    .X(_05440_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13168_ (.A(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__and3_1 _13169_ (.A(net7802),
    .B(net3687),
    .C(net2970),
    .X(_05442_));
 sky130_fd_sc_hd__and3_1 _13170_ (.A(net7778),
    .B(net2334),
    .C(net2974),
    .X(_05443_));
 sky130_fd_sc_hd__xnor2_1 _13171_ (.A(_05442_),
    .B(_05443_),
    .Y(_05444_));
 sky130_fd_sc_hd__xnor2_1 _13172_ (.A(_05441_),
    .B(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__a21oi_1 _13173_ (.A1(net1137),
    .A2(net1136),
    .B1(_05445_),
    .Y(_05446_));
 sky130_fd_sc_hd__and3_1 _13174_ (.A(_05445_),
    .B(net1137),
    .C(net1136),
    .X(_05447_));
 sky130_fd_sc_hd__or4_1 _13175_ (.A(_05432_),
    .B(_05433_),
    .C(net1000),
    .D(net999),
    .X(_05448_));
 sky130_fd_sc_hd__o22ai_2 _13176_ (.A1(_05432_),
    .A2(_05433_),
    .B1(net1000),
    .B2(net999),
    .Y(_05449_));
 sky130_fd_sc_hd__nand2_1 _13177_ (.A(net7740),
    .B(net1353),
    .Y(_05450_));
 sky130_fd_sc_hd__and3_1 _13178_ (.A(net7714),
    .B(net1976),
    .C(net2312),
    .X(_05451_));
 sky130_fd_sc_hd__and3_1 _13179_ (.A(net7732),
    .B(net1983),
    .C(net2361),
    .X(_05452_));
 sky130_fd_sc_hd__xor2_1 _13180_ (.A(_05451_),
    .B(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__xnor2_1 _13181_ (.A(_05450_),
    .B(_05453_),
    .Y(_05454_));
 sky130_fd_sc_hd__a21o_1 _13182_ (.A1(_05366_),
    .A2(_05367_),
    .B1(_05368_),
    .X(_05455_));
 sky130_fd_sc_hd__o21a_1 _13183_ (.A1(_05366_),
    .A2(_05367_),
    .B1(_05455_),
    .X(_05456_));
 sky130_fd_sc_hd__nand2_1 _13184_ (.A(net7672),
    .B(_05216_),
    .Y(_05457_));
 sky130_fd_sc_hd__and3_1 _13185_ (.A(net7650),
    .B(net2339),
    .C(net1967),
    .X(_05458_));
 sky130_fd_sc_hd__and3_1 _13186_ (.A(net7689),
    .B(net2350),
    .C(net2346),
    .X(_05459_));
 sky130_fd_sc_hd__xor2_1 _13187_ (.A(_05458_),
    .B(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__xnor2_2 _13188_ (.A(_05457_),
    .B(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__xnor2_1 _13189_ (.A(_05456_),
    .B(_05461_),
    .Y(_05462_));
 sky130_fd_sc_hd__xnor2_1 _13190_ (.A(_05454_),
    .B(_05462_),
    .Y(_05463_));
 sky130_fd_sc_hd__a21o_1 _13191_ (.A1(_05448_),
    .A2(_05449_),
    .B1(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__nand3_1 _13192_ (.A(_05463_),
    .B(_05448_),
    .C(_05449_),
    .Y(_05465_));
 sky130_fd_sc_hd__nand2_1 _13193_ (.A(_05464_),
    .B(_05465_),
    .Y(_05466_));
 sky130_fd_sc_hd__nor2_1 _13194_ (.A(_05382_),
    .B(net849),
    .Y(_05467_));
 sky130_fd_sc_hd__a21oi_1 _13195_ (.A1(_05382_),
    .A2(net849),
    .B1(_05379_),
    .Y(_05468_));
 sky130_fd_sc_hd__or2_1 _13196_ (.A(_05467_),
    .B(_05468_),
    .X(_05469_));
 sky130_fd_sc_hd__xor2_1 _13197_ (.A(_05466_),
    .B(_05469_),
    .X(_05470_));
 sky130_fd_sc_hd__xnor2_2 _13198_ (.A(net733),
    .B(net682),
    .Y(_05471_));
 sky130_fd_sc_hd__xnor2_1 _13199_ (.A(net919),
    .B(_05360_),
    .Y(_05472_));
 sky130_fd_sc_hd__a21o_1 _13200_ (.A1(_05362_),
    .A2(_05363_),
    .B1(_05472_),
    .X(_05473_));
 sky130_fd_sc_hd__and3_1 _13201_ (.A(_05472_),
    .B(_05362_),
    .C(_05363_),
    .X(_05474_));
 sky130_fd_sc_hd__a21oi_2 _13202_ (.A1(net734),
    .A2(_05473_),
    .B1(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__inv_2 _13203_ (.A(net1001),
    .Y(_05476_));
 sky130_fd_sc_hd__and2_1 _13204_ (.A(net919),
    .B(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__o21a_1 _13205_ (.A1(net919),
    .A2(_05476_),
    .B1(_05357_),
    .X(_05478_));
 sky130_fd_sc_hd__or2_1 _13206_ (.A(_05477_),
    .B(_05478_),
    .X(_05479_));
 sky130_fd_sc_hd__xnor2_1 _13207_ (.A(_05475_),
    .B(_05479_),
    .Y(_05480_));
 sky130_fd_sc_hd__xnor2_1 _13208_ (.A(_05471_),
    .B(_05480_),
    .Y(_05481_));
 sky130_fd_sc_hd__nand2_1 _13209_ (.A(_05405_),
    .B(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__and2b_1 _13210_ (.A_N(_05431_),
    .B(_05479_),
    .X(_05483_));
 sky130_fd_sc_hd__and2_1 _13211_ (.A(_05431_),
    .B(_05479_),
    .X(_05484_));
 sky130_fd_sc_hd__mux2_1 _13212_ (.A0(_05483_),
    .A1(_05484_),
    .S(net682),
    .X(_05485_));
 sky130_fd_sc_hd__o32ai_4 _13213_ (.A1(_05471_),
    .A2(_05477_),
    .A3(_05478_),
    .B1(_05485_),
    .B2(_05475_),
    .Y(_05486_));
 sky130_fd_sc_hd__and3_1 _13214_ (.A(net7728),
    .B(net2368),
    .C(net2365),
    .X(_05487_));
 sky130_fd_sc_hd__nand2_1 _13215_ (.A(net7690),
    .B(net1340),
    .Y(_05488_));
 sky130_fd_sc_hd__nand2_1 _13216_ (.A(net7713),
    .B(net1606),
    .Y(_05489_));
 sky130_fd_sc_hd__xor2_1 _13217_ (.A(_05488_),
    .B(_05489_),
    .X(_05490_));
 sky130_fd_sc_hd__xor2_2 _13218_ (.A(net1946),
    .B(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__a21o_1 _13219_ (.A1(net7672),
    .A2(_05216_),
    .B1(_05458_),
    .X(_05492_));
 sky130_fd_sc_hd__and3_1 _13220_ (.A(net7672),
    .B(_05216_),
    .C(_05458_),
    .X(_05493_));
 sky130_fd_sc_hd__a21o_1 _13221_ (.A1(_05459_),
    .A2(_05492_),
    .B1(_05493_),
    .X(_05494_));
 sky130_fd_sc_hd__and3_1 _13222_ (.A(net7650),
    .B(net1972),
    .C(net1969),
    .X(_05495_));
 sky130_fd_sc_hd__and3_1 _13223_ (.A(net7640),
    .B(net2339),
    .C(net1967),
    .X(_05496_));
 sky130_fd_sc_hd__and3_1 _13224_ (.A(net7674),
    .B(net2350),
    .C(net2346),
    .X(_05497_));
 sky130_fd_sc_hd__xor2_1 _13225_ (.A(_05496_),
    .B(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__xnor2_1 _13226_ (.A(_05495_),
    .B(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__xor2_1 _13227_ (.A(net1135),
    .B(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__xnor2_2 _13228_ (.A(_05491_),
    .B(_05500_),
    .Y(_05501_));
 sky130_fd_sc_hd__a21o_1 _13229_ (.A1(_05456_),
    .A2(_05461_),
    .B1(_05454_),
    .X(_05502_));
 sky130_fd_sc_hd__o21a_1 _13230_ (.A1(_05456_),
    .A2(_05461_),
    .B1(_05502_),
    .X(_05503_));
 sky130_fd_sc_hd__clkbuf_1 _13231_ (.A(_04960_),
    .X(_05504_));
 sky130_fd_sc_hd__nand2_1 _13232_ (.A(net7755),
    .B(_05504_),
    .Y(_05505_));
 sky130_fd_sc_hd__and3_1 _13233_ (.A(net7780),
    .B(net3685),
    .C(net2967),
    .X(_05506_));
 sky130_fd_sc_hd__and3_1 _13234_ (.A(net7745),
    .B(net2321),
    .C(net2317),
    .X(_05507_));
 sky130_fd_sc_hd__xnor2_1 _13235_ (.A(_05506_),
    .B(_05507_),
    .Y(_05508_));
 sky130_fd_sc_hd__xnor2_2 _13236_ (.A(_05505_),
    .B(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hd__a22o_1 _13237_ (.A1(net7740),
    .A2(net1353),
    .B1(_05451_),
    .B2(_05452_),
    .X(_05510_));
 sky130_fd_sc_hd__o21a_1 _13238_ (.A1(_05451_),
    .A2(_05452_),
    .B1(_05510_),
    .X(_05511_));
 sky130_fd_sc_hd__a21o_1 _13239_ (.A1(_05441_),
    .A2(_05443_),
    .B1(_05442_),
    .X(_05512_));
 sky130_fd_sc_hd__o21a_1 _13240_ (.A1(_05441_),
    .A2(_05443_),
    .B1(_05512_),
    .X(_05513_));
 sky130_fd_sc_hd__xor2_1 _13241_ (.A(_05511_),
    .B(net1133),
    .X(_05514_));
 sky130_fd_sc_hd__xnor2_2 _13242_ (.A(_05509_),
    .B(_05514_),
    .Y(_05515_));
 sky130_fd_sc_hd__xor2_1 _13243_ (.A(net847),
    .B(_05515_),
    .X(_05516_));
 sky130_fd_sc_hd__xnor2_1 _13244_ (.A(_05501_),
    .B(_05516_),
    .Y(_05517_));
 sky130_fd_sc_hd__and2_1 _13245_ (.A(net7845),
    .B(net1947),
    .X(_05518_));
 sky130_fd_sc_hd__and3_1 _13246_ (.A(net7808),
    .B(net2309),
    .C(net1954),
    .X(_05519_));
 sky130_fd_sc_hd__clkbuf_2 _13247_ (.A(_05519_),
    .X(_05520_));
 sky130_fd_sc_hd__and3_1 _13248_ (.A(net7821),
    .B(net2304),
    .C(net2964),
    .X(_05521_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _13249_ (.A(_05521_),
    .X(_05522_));
 sky130_fd_sc_hd__xor2_1 _13250_ (.A(_05520_),
    .B(_05522_),
    .X(_05523_));
 sky130_fd_sc_hd__xnor2_1 _13251_ (.A(_05518_),
    .B(_05523_),
    .Y(_05524_));
 sky130_fd_sc_hd__a22o_1 _13252_ (.A1(net7879),
    .A2(net1948),
    .B1(_05413_),
    .B2(_05414_),
    .X(_05525_));
 sky130_fd_sc_hd__o21a_1 _13253_ (.A1(_05413_),
    .A2(_05414_),
    .B1(_05525_),
    .X(_05526_));
 sky130_fd_sc_hd__nor2_1 _13254_ (.A(net2301),
    .B(net2297),
    .Y(_05527_));
 sky130_fd_sc_hd__and2_1 _13255_ (.A(net7923),
    .B(_05527_),
    .X(_05528_));
 sky130_fd_sc_hd__and3b_1 _13256_ (.A_N(net6672),
    .B(net6678),
    .C(net7208),
    .X(_05529_));
 sky130_fd_sc_hd__and3b_1 _13257_ (.A_N(net6677),
    .B(net5193),
    .C(net6672),
    .X(_05530_));
 sky130_fd_sc_hd__o21ai_1 _13258_ (.A1(_05529_),
    .A2(_05530_),
    .B1(_05052_),
    .Y(_05531_));
 sky130_fd_sc_hd__nand2_1 _13259_ (.A(\svm0.vC[14] ),
    .B(net2992),
    .Y(_05532_));
 sky130_fd_sc_hd__and3_1 _13260_ (.A(net7946),
    .B(net3682),
    .C(net2294),
    .X(_05533_));
 sky130_fd_sc_hd__and3_1 _13261_ (.A(net7879),
    .B(net3684),
    .C(net4254),
    .X(_05534_));
 sky130_fd_sc_hd__xnor2_1 _13262_ (.A(_05533_),
    .B(_05534_),
    .Y(_05535_));
 sky130_fd_sc_hd__xnor2_2 _13263_ (.A(_05528_),
    .B(_05535_),
    .Y(_05536_));
 sky130_fd_sc_hd__xor2_1 _13264_ (.A(net1330),
    .B(_05536_),
    .X(_05537_));
 sky130_fd_sc_hd__xor2_1 _13265_ (.A(_05524_),
    .B(_05537_),
    .X(_05538_));
 sky130_fd_sc_hd__and2_1 _13266_ (.A(_05417_),
    .B(_05418_),
    .X(_05539_));
 sky130_fd_sc_hd__xor2_1 _13267_ (.A(_05412_),
    .B(_05415_),
    .X(_05540_));
 sky130_fd_sc_hd__or2_1 _13268_ (.A(_05539_),
    .B(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__a21o_1 _13269_ (.A1(_05539_),
    .A2(_05540_),
    .B1(_05423_),
    .X(_05542_));
 sky130_fd_sc_hd__xor2_1 _13270_ (.A(_05441_),
    .B(_05444_),
    .X(_05543_));
 sky130_fd_sc_hd__a21bo_1 _13271_ (.A1(_05543_),
    .A2(net1136),
    .B1_N(net1137),
    .X(_05544_));
 sky130_fd_sc_hd__a21oi_1 _13272_ (.A1(_05541_),
    .A2(_05542_),
    .B1(_05544_),
    .Y(_05545_));
 sky130_fd_sc_hd__and3_1 _13273_ (.A(_05544_),
    .B(_05541_),
    .C(_05542_),
    .X(_05546_));
 sky130_fd_sc_hd__or3_1 _13274_ (.A(_05538_),
    .B(_05545_),
    .C(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__o21ai_1 _13275_ (.A1(_05545_),
    .A2(_05546_),
    .B1(_05538_),
    .Y(_05548_));
 sky130_fd_sc_hd__a21boi_1 _13276_ (.A1(_05463_),
    .A2(_05449_),
    .B1_N(_05448_),
    .Y(_05549_));
 sky130_fd_sc_hd__and3_1 _13277_ (.A(_05547_),
    .B(_05548_),
    .C(net846),
    .X(_05550_));
 sky130_fd_sc_hd__a21oi_1 _13278_ (.A1(_05547_),
    .A2(_05548_),
    .B1(net846),
    .Y(_05551_));
 sky130_fd_sc_hd__nor2_1 _13279_ (.A(_05550_),
    .B(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__xnor2_2 _13280_ (.A(net732),
    .B(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__a21oi_2 _13281_ (.A1(net918),
    .A2(_05429_),
    .B1(_05428_),
    .Y(_05554_));
 sky130_fd_sc_hd__clkbuf_1 _13282_ (.A(_05527_),
    .X(_05555_));
 sky130_fd_sc_hd__clkbuf_1 _13283_ (.A(net1575),
    .X(_05556_));
 sky130_fd_sc_hd__and3_1 _13284_ (.A(net3688),
    .B(net2303),
    .C(net1321),
    .X(_05557_));
 sky130_fd_sc_hd__xnor2_2 _13285_ (.A(_05554_),
    .B(net1132),
    .Y(_05558_));
 sky130_fd_sc_hd__a211o_1 _13286_ (.A1(_05464_),
    .A2(_05465_),
    .B1(_05468_),
    .C1(_05467_),
    .X(_05559_));
 sky130_fd_sc_hd__o211a_1 _13287_ (.A1(_05467_),
    .A2(_05468_),
    .B1(_05465_),
    .C1(_05464_),
    .X(_05560_));
 sky130_fd_sc_hd__a21o_1 _13288_ (.A1(net733),
    .A2(_05559_),
    .B1(_05560_),
    .X(_05561_));
 sky130_fd_sc_hd__xnor2_1 _13289_ (.A(_05558_),
    .B(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__xnor2_1 _13290_ (.A(_05553_),
    .B(_05562_),
    .Y(_05563_));
 sky130_fd_sc_hd__xor2_1 _13291_ (.A(_05486_),
    .B(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__nand2_1 _13292_ (.A(_05482_),
    .B(_05564_),
    .Y(_05565_));
 sky130_fd_sc_hd__or2_1 _13293_ (.A(_05482_),
    .B(_05564_),
    .X(_05566_));
 sky130_fd_sc_hd__xor2_1 _13294_ (.A(net732),
    .B(_05552_),
    .X(_05567_));
 sky130_fd_sc_hd__and2b_1 _13295_ (.A_N(_05561_),
    .B(_05558_),
    .X(_05568_));
 sky130_fd_sc_hd__or2b_1 _13296_ (.A(_05558_),
    .B_N(_05561_),
    .X(_05569_));
 sky130_fd_sc_hd__o21ai_2 _13297_ (.A1(_05567_),
    .A2(_05568_),
    .B1(_05569_),
    .Y(_05570_));
 sky130_fd_sc_hd__inv_2 _13298_ (.A(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__a21o_1 _13299_ (.A1(_05501_),
    .A2(_05515_),
    .B1(net847),
    .X(_05572_));
 sky130_fd_sc_hd__o21a_1 _13300_ (.A1(_05501_),
    .A2(_05515_),
    .B1(_05572_),
    .X(_05573_));
 sky130_fd_sc_hd__or2b_1 _13301_ (.A(net1135),
    .B_N(_05499_),
    .X(_05574_));
 sky130_fd_sc_hd__and2b_1 _13302_ (.A_N(_05499_),
    .B(net1135),
    .X(_05575_));
 sky130_fd_sc_hd__a21o_1 _13303_ (.A1(_05491_),
    .A2(_05574_),
    .B1(_05575_),
    .X(_05576_));
 sky130_fd_sc_hd__and3_1 _13304_ (.A(net7640),
    .B(net1972),
    .C(net1969),
    .X(_05577_));
 sky130_fd_sc_hd__and3_1 _13305_ (.A(net7619),
    .B(net2339),
    .C(net1967),
    .X(_05578_));
 sky130_fd_sc_hd__and3_1 _13306_ (.A(net7650),
    .B(net2350),
    .C(net2346),
    .X(_05579_));
 sky130_fd_sc_hd__xor2_1 _13307_ (.A(net1572),
    .B(net1945),
    .X(_05580_));
 sky130_fd_sc_hd__xnor2_1 _13308_ (.A(net1574),
    .B(_05580_),
    .Y(_05581_));
 sky130_fd_sc_hd__a21o_1 _13309_ (.A1(_05495_),
    .A2(_05496_),
    .B1(_05497_),
    .X(_05582_));
 sky130_fd_sc_hd__o21ai_1 _13310_ (.A1(_05495_),
    .A2(_05496_),
    .B1(_05582_),
    .Y(_05583_));
 sky130_fd_sc_hd__nand2_1 _13311_ (.A(net7705),
    .B(net1352),
    .Y(_05584_));
 sky130_fd_sc_hd__and3_1 _13312_ (.A(net7671),
    .B(net1975),
    .C(net2311),
    .X(_05585_));
 sky130_fd_sc_hd__and3_1 _13313_ (.A(net7698),
    .B(net1982),
    .C(net2360),
    .X(_05586_));
 sky130_fd_sc_hd__xnor2_1 _13314_ (.A(_05585_),
    .B(_05586_),
    .Y(_05587_));
 sky130_fd_sc_hd__xnor2_2 _13315_ (.A(_05584_),
    .B(_05587_),
    .Y(_05588_));
 sky130_fd_sc_hd__xnor2_1 _13316_ (.A(net1131),
    .B(_05588_),
    .Y(_05589_));
 sky130_fd_sc_hd__xor2_1 _13317_ (.A(_05581_),
    .B(_05589_),
    .X(_05590_));
 sky130_fd_sc_hd__nand2_1 _13318_ (.A(net7769),
    .B(net1598),
    .Y(_05591_));
 sky130_fd_sc_hd__and3_1 _13319_ (.A(net7722),
    .B(net2321),
    .C(net2317),
    .X(_05592_));
 sky130_fd_sc_hd__and3_1 _13320_ (.A(net7747),
    .B(net2330),
    .C(net2325),
    .X(_05593_));
 sky130_fd_sc_hd__xor2_1 _13321_ (.A(_05592_),
    .B(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__xnor2_1 _13322_ (.A(_05591_),
    .B(_05594_),
    .Y(_05595_));
 sky130_fd_sc_hd__a31o_1 _13323_ (.A1(net7774),
    .A2(_04960_),
    .A3(_05507_),
    .B1(_05506_),
    .X(_05596_));
 sky130_fd_sc_hd__a21o_1 _13324_ (.A1(net7774),
    .A2(_04960_),
    .B1(_05507_),
    .X(_05597_));
 sky130_fd_sc_hd__nand2_1 _13325_ (.A(_05596_),
    .B(_05597_),
    .Y(_05598_));
 sky130_fd_sc_hd__a22o_1 _13326_ (.A1(net7710),
    .A2(net1605),
    .B1(net1339),
    .B2(net7687),
    .X(_05599_));
 sky130_fd_sc_hd__a41o_1 _13327_ (.A1(net7713),
    .A2(net7687),
    .A3(net1606),
    .A4(net1339),
    .B1(net1946),
    .X(_05600_));
 sky130_fd_sc_hd__and2_1 _13328_ (.A(_05599_),
    .B(_05600_),
    .X(_05601_));
 sky130_fd_sc_hd__xnor2_1 _13329_ (.A(_05598_),
    .B(_05601_),
    .Y(_05602_));
 sky130_fd_sc_hd__xor2_1 _13330_ (.A(_05595_),
    .B(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__xnor2_1 _13331_ (.A(_05590_),
    .B(net844),
    .Y(_05604_));
 sky130_fd_sc_hd__xnor2_1 _13332_ (.A(net845),
    .B(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hd__nand2_1 _13333_ (.A(net7827),
    .B(net1590),
    .Y(_05606_));
 sky130_fd_sc_hd__and3_1 _13334_ (.A(net7792),
    .B(net2307),
    .C(net1952),
    .X(_05607_));
 sky130_fd_sc_hd__buf_1 _13335_ (.A(net2304),
    .X(_05608_));
 sky130_fd_sc_hd__buf_1 _13336_ (.A(net2964),
    .X(_05609_));
 sky130_fd_sc_hd__and3_1 _13337_ (.A(net7815),
    .B(net1942),
    .C(net2291),
    .X(_05610_));
 sky130_fd_sc_hd__xor2_1 _13338_ (.A(_05607_),
    .B(_05610_),
    .X(_05611_));
 sky130_fd_sc_hd__xnor2_1 _13339_ (.A(_05606_),
    .B(net1320),
    .Y(_05612_));
 sky130_fd_sc_hd__a21oi_1 _13340_ (.A1(_05520_),
    .A2(_05522_),
    .B1(_05518_),
    .Y(_05613_));
 sky130_fd_sc_hd__nor2_1 _13341_ (.A(_05520_),
    .B(_05522_),
    .Y(_05614_));
 sky130_fd_sc_hd__o21a_1 _13342_ (.A1(_05343_),
    .A2(_05344_),
    .B1(_05052_),
    .X(_05615_));
 sky130_fd_sc_hd__nand2_1 _13343_ (.A(net7869),
    .B(net4254),
    .Y(_05616_));
 sky130_fd_sc_hd__buf_1 _13344_ (.A(net2294),
    .X(_05617_));
 sky130_fd_sc_hd__o2111a_1 _13345_ (.A1(net3679),
    .A2(net3675),
    .B1(net3682),
    .C1(net7923),
    .D1(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__buf_1 _13346_ (.A(net3682),
    .X(_05619_));
 sky130_fd_sc_hd__a311oi_2 _13347_ (.A1(net7923),
    .A2(_05619_),
    .A3(net2294),
    .B1(net3675),
    .C1(net3679),
    .Y(_05620_));
 sky130_fd_sc_hd__a211o_1 _13348_ (.A1(net7893),
    .A2(_05527_),
    .B1(_05618_),
    .C1(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__o211ai_2 _13349_ (.A1(_05618_),
    .A2(_05620_),
    .B1(net7893),
    .C1(_05527_),
    .Y(_05622_));
 sky130_fd_sc_hd__o211a_1 _13350_ (.A1(_05613_),
    .A2(_05614_),
    .B1(_05621_),
    .C1(_05622_),
    .X(_05623_));
 sky130_fd_sc_hd__a211o_1 _13351_ (.A1(_05621_),
    .A2(_05622_),
    .B1(_05613_),
    .C1(_05614_),
    .X(_05624_));
 sky130_fd_sc_hd__and2b_1 _13352_ (.A_N(_05623_),
    .B(_05624_),
    .X(_05625_));
 sky130_fd_sc_hd__xnor2_1 _13353_ (.A(_05612_),
    .B(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__nand2_1 _13354_ (.A(_05511_),
    .B(net1133),
    .Y(_05627_));
 sky130_fd_sc_hd__nor2_1 _13355_ (.A(_05511_),
    .B(net1133),
    .Y(_05628_));
 sky130_fd_sc_hd__a21o_1 _13356_ (.A1(_05509_),
    .A2(_05627_),
    .B1(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__a21bo_1 _13357_ (.A1(net1330),
    .A2(_05536_),
    .B1_N(_05524_),
    .X(_05630_));
 sky130_fd_sc_hd__o21a_1 _13358_ (.A1(net1330),
    .A2(_05536_),
    .B1(_05630_),
    .X(_05631_));
 sky130_fd_sc_hd__xor2_1 _13359_ (.A(_05629_),
    .B(net842),
    .X(_05632_));
 sky130_fd_sc_hd__xnor2_2 _13360_ (.A(net843),
    .B(_05632_),
    .Y(_05633_));
 sky130_fd_sc_hd__xor2_1 _13361_ (.A(net731),
    .B(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__xnor2_1 _13362_ (.A(_05573_),
    .B(_05634_),
    .Y(_05635_));
 sky130_fd_sc_hd__o21ba_1 _13363_ (.A1(net732),
    .A2(_05550_),
    .B1_N(_05551_),
    .X(_05636_));
 sky130_fd_sc_hd__a21boi_1 _13364_ (.A1(_05543_),
    .A2(net1136),
    .B1_N(net1137),
    .Y(_05637_));
 sky130_fd_sc_hd__nand3_1 _13365_ (.A(_05637_),
    .B(_05541_),
    .C(_05542_),
    .Y(_05638_));
 sky130_fd_sc_hd__a31o_1 _13366_ (.A1(net7926),
    .A2(net1582),
    .A3(_05534_),
    .B1(_05533_),
    .X(_05639_));
 sky130_fd_sc_hd__o21a_1 _13367_ (.A1(_05528_),
    .A2(_05534_),
    .B1(_05639_),
    .X(_05640_));
 sky130_fd_sc_hd__a22o_1 _13368_ (.A1(net5189),
    .A2(net2963),
    .B1(net2986),
    .B2(net7199),
    .X(_05641_));
 sky130_fd_sc_hd__a22o_1 _13369_ (.A1(\svm0.vC[15] ),
    .A2(net2378),
    .B1(_05641_),
    .B2(net3028),
    .X(_05642_));
 sky130_fd_sc_hd__nand2_1 _13370_ (.A(net7947),
    .B(net1935),
    .Y(_05643_));
 sky130_fd_sc_hd__xor2_1 _13371_ (.A(net1130),
    .B(_05643_),
    .X(_05644_));
 sky130_fd_sc_hd__a21o_1 _13372_ (.A1(_05541_),
    .A2(_05542_),
    .B1(_05637_),
    .X(_05645_));
 sky130_fd_sc_hd__xnor2_1 _13373_ (.A(net1130),
    .B(_05643_),
    .Y(_05646_));
 sky130_fd_sc_hd__nand2_1 _13374_ (.A(_05538_),
    .B(_05638_),
    .Y(_05647_));
 sky130_fd_sc_hd__and3_1 _13375_ (.A(_05645_),
    .B(_05646_),
    .C(_05647_),
    .X(_05648_));
 sky130_fd_sc_hd__nor2_1 _13376_ (.A(_05645_),
    .B(_05646_),
    .Y(_05649_));
 sky130_fd_sc_hd__a311o_1 _13377_ (.A1(_05538_),
    .A2(_05638_),
    .A3(_05644_),
    .B1(_05648_),
    .C1(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__xor2_1 _13378_ (.A(_05636_),
    .B(_05650_),
    .X(_05651_));
 sky130_fd_sc_hd__xnor2_1 _13379_ (.A(net628),
    .B(_05651_),
    .Y(_05652_));
 sky130_fd_sc_hd__nand2_1 _13380_ (.A(_05554_),
    .B(net1132),
    .Y(_05653_));
 sky130_fd_sc_hd__xnor2_1 _13381_ (.A(_05652_),
    .B(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__a221o_1 _13382_ (.A1(_05567_),
    .A2(_05568_),
    .B1(_05571_),
    .B2(_05486_),
    .C1(_05654_),
    .X(_05655_));
 sky130_fd_sc_hd__nand2_1 _13383_ (.A(_05553_),
    .B(_05561_),
    .Y(_05656_));
 sky130_fd_sc_hd__nor2_1 _13384_ (.A(_05486_),
    .B(_05558_),
    .Y(_05657_));
 sky130_fd_sc_hd__xnor2_1 _13385_ (.A(_05553_),
    .B(_05561_),
    .Y(_05658_));
 sky130_fd_sc_hd__o221ai_1 _13386_ (.A1(_05656_),
    .A2(_05657_),
    .B1(_05658_),
    .B2(_05558_),
    .C1(_05654_),
    .Y(_05659_));
 sky130_fd_sc_hd__a22o_1 _13387_ (.A1(_05565_),
    .A2(_05566_),
    .B1(_05655_),
    .B2(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__xnor2_1 _13388_ (.A(_05405_),
    .B(_05481_),
    .Y(_05661_));
 sky130_fd_sc_hd__xor2_2 _13389_ (.A(net683),
    .B(net848),
    .X(_05662_));
 sky130_fd_sc_hd__xor2_1 _13390_ (.A(_05401_),
    .B(_05662_),
    .X(_05663_));
 sky130_fd_sc_hd__nor2_1 _13391_ (.A(_05247_),
    .B(_05245_),
    .Y(_05664_));
 sky130_fd_sc_hd__a21o_1 _13392_ (.A1(net684),
    .A2(_05664_),
    .B1(_05307_),
    .X(_05665_));
 sky130_fd_sc_hd__o21ai_1 _13393_ (.A1(net684),
    .A2(_05664_),
    .B1(_05665_),
    .Y(_05666_));
 sky130_fd_sc_hd__nand3_1 _13394_ (.A(net583),
    .B(_05663_),
    .C(net581),
    .Y(_05667_));
 sky130_fd_sc_hd__xnor2_1 _13395_ (.A(_05401_),
    .B(_05662_),
    .Y(_05668_));
 sky130_fd_sc_hd__or3_1 _13396_ (.A(net583),
    .B(_05668_),
    .C(net581),
    .X(_05669_));
 sky130_fd_sc_hd__or3b_1 _13397_ (.A(net583),
    .B(_05663_),
    .C_N(net581),
    .X(_05670_));
 sky130_fd_sc_hd__mux2_1 _13398_ (.A0(_05669_),
    .A1(_05670_),
    .S(_05661_),
    .X(_05671_));
 sky130_fd_sc_hd__or4b_1 _13399_ (.A(_05663_),
    .B(net581),
    .C(_05661_),
    .D_N(net583),
    .X(_05672_));
 sky130_fd_sc_hd__o211a_1 _13400_ (.A1(_05661_),
    .A2(_05667_),
    .B1(_05671_),
    .C1(_05672_),
    .X(_05673_));
 sky130_fd_sc_hd__nor2_1 _13401_ (.A(_05486_),
    .B(_05563_),
    .Y(_05674_));
 sky130_fd_sc_hd__o2bb2a_1 _13402_ (.A1_N(_05563_),
    .A2_N(_05486_),
    .B1(_05481_),
    .B2(_05405_),
    .X(_05675_));
 sky130_fd_sc_hd__nor2_1 _13403_ (.A(_05674_),
    .B(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__o21bai_1 _13404_ (.A1(_05668_),
    .A2(net581),
    .B1_N(net583),
    .Y(_05677_));
 sky130_fd_sc_hd__a21oi_1 _13405_ (.A1(_05668_),
    .A2(net581),
    .B1(_05674_),
    .Y(_05678_));
 sky130_fd_sc_hd__xnor2_1 _13406_ (.A(_05654_),
    .B(_05570_),
    .Y(_05679_));
 sky130_fd_sc_hd__a31o_1 _13407_ (.A1(_05482_),
    .A2(_05677_),
    .A3(_05678_),
    .B1(_05679_),
    .X(_05680_));
 sky130_fd_sc_hd__o32a_1 _13408_ (.A1(net452),
    .A2(_05660_),
    .A3(_05673_),
    .B1(_05676_),
    .B2(_05680_),
    .X(_05681_));
 sky130_fd_sc_hd__and2b_1 _13409_ (.A_N(_05652_),
    .B(_05656_),
    .X(_05682_));
 sky130_fd_sc_hd__a2bb2o_1 _13410_ (.A1_N(_05653_),
    .A2_N(_05682_),
    .B1(_05570_),
    .B2(_05652_),
    .X(_05683_));
 sky130_fd_sc_hd__a21o_1 _13411_ (.A1(net731),
    .A2(_05633_),
    .B1(_05573_),
    .X(_05684_));
 sky130_fd_sc_hd__o21ai_1 _13412_ (.A1(net731),
    .A2(_05633_),
    .B1(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__and2_1 _13413_ (.A(net2949),
    .B(net1941),
    .X(_05686_));
 sky130_fd_sc_hd__buf_1 _13414_ (.A(_05686_),
    .X(_05687_));
 sky130_fd_sc_hd__nand2_1 _13415_ (.A(net7900),
    .B(net1327),
    .Y(_05688_));
 sky130_fd_sc_hd__or2_1 _13416_ (.A(net3678),
    .B(net3675),
    .X(_05689_));
 sky130_fd_sc_hd__nand2_1 _13417_ (.A(_05688_),
    .B(net2944),
    .Y(_05690_));
 sky130_fd_sc_hd__nor2_1 _13418_ (.A(_05688_),
    .B(net2944),
    .Y(_05691_));
 sky130_fd_sc_hd__a31o_1 _13419_ (.A1(net7921),
    .A2(net1317),
    .A3(_05690_),
    .B1(_05691_),
    .X(_05692_));
 sky130_fd_sc_hd__and3_1 _13420_ (.A(net7921),
    .B(net1929),
    .C(_05692_),
    .X(_05693_));
 sky130_fd_sc_hd__a21o_1 _13421_ (.A1(net7921),
    .A2(net1929),
    .B1(_05692_),
    .X(_05694_));
 sky130_fd_sc_hd__and2b_1 _13422_ (.A_N(_05693_),
    .B(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__o21ba_1 _13423_ (.A1(net843),
    .A2(net842),
    .B1_N(_05629_),
    .X(_05696_));
 sky130_fd_sc_hd__a21o_1 _13424_ (.A1(net843),
    .A2(net842),
    .B1(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__xnor2_2 _13425_ (.A(_05695_),
    .B(net728),
    .Y(_05698_));
 sky130_fd_sc_hd__or2_1 _13426_ (.A(_05590_),
    .B(net844),
    .X(_05699_));
 sky130_fd_sc_hd__nand2_1 _13427_ (.A(net7815),
    .B(net1586),
    .Y(_05700_));
 sky130_fd_sc_hd__and3_1 _13428_ (.A(net7770),
    .B(net2307),
    .C(net1952),
    .X(_05701_));
 sky130_fd_sc_hd__and3_1 _13429_ (.A(net7792),
    .B(net1942),
    .C(net2291),
    .X(_05702_));
 sky130_fd_sc_hd__xnor2_1 _13430_ (.A(_05701_),
    .B(_05702_),
    .Y(_05703_));
 sky130_fd_sc_hd__xnor2_2 _13431_ (.A(_05700_),
    .B(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hd__a22o_1 _13432_ (.A1(net7834),
    .A2(net1587),
    .B1(_05607_),
    .B2(_05610_),
    .X(_05705_));
 sky130_fd_sc_hd__o21ai_1 _13433_ (.A1(_05607_),
    .A2(_05610_),
    .B1(_05705_),
    .Y(_05706_));
 sky130_fd_sc_hd__nand2_1 _13434_ (.A(net7866),
    .B(net1577),
    .Y(_05707_));
 sky130_fd_sc_hd__and3_1 _13435_ (.A(net7901),
    .B(net2946),
    .C(net1938),
    .X(_05708_));
 sky130_fd_sc_hd__clkbuf_1 _13436_ (.A(net4255),
    .X(_05709_));
 sky130_fd_sc_hd__and3_1 _13437_ (.A(net7832),
    .B(net2950),
    .C(net3669),
    .X(_05710_));
 sky130_fd_sc_hd__xnor2_1 _13438_ (.A(_05708_),
    .B(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__xnor2_1 _13439_ (.A(_05707_),
    .B(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__xor2_1 _13440_ (.A(net1129),
    .B(net1128),
    .X(_05713_));
 sky130_fd_sc_hd__xnor2_1 _13441_ (.A(_05704_),
    .B(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__o211a_1 _13442_ (.A1(_05506_),
    .A2(_05507_),
    .B1(net7769),
    .C1(net1584),
    .X(_05715_));
 sky130_fd_sc_hd__and3_1 _13443_ (.A(net7745),
    .B(net1963),
    .C(_05506_),
    .X(_05716_));
 sky130_fd_sc_hd__and4_1 _13444_ (.A(_05596_),
    .B(_05597_),
    .C(_05599_),
    .D(_05600_),
    .X(_05717_));
 sky130_fd_sc_hd__o32a_1 _13445_ (.A1(_05715_),
    .A2(_05716_),
    .A3(_05601_),
    .B1(_05717_),
    .B2(_05595_),
    .X(_05718_));
 sky130_fd_sc_hd__a22o_1 _13446_ (.A1(net7860),
    .A2(net1590),
    .B1(_05520_),
    .B2(_05522_),
    .X(_05719_));
 sky130_fd_sc_hd__or2_1 _13447_ (.A(_05520_),
    .B(_05522_),
    .X(_05720_));
 sky130_fd_sc_hd__a22o_1 _13448_ (.A1(_05719_),
    .A2(_05720_),
    .B1(_05621_),
    .B2(_05622_),
    .X(_05721_));
 sky130_fd_sc_hd__and4_1 _13449_ (.A(_05719_),
    .B(_05720_),
    .C(_05621_),
    .D(_05622_),
    .X(_05722_));
 sky130_fd_sc_hd__a21o_1 _13450_ (.A1(_05612_),
    .A2(_05721_),
    .B1(_05722_),
    .X(_05723_));
 sky130_fd_sc_hd__xnor2_1 _13451_ (.A(net915),
    .B(net913),
    .Y(_05724_));
 sky130_fd_sc_hd__xnor2_1 _13452_ (.A(net916),
    .B(_05724_),
    .Y(_05725_));
 sky130_fd_sc_hd__a21o_1 _13453_ (.A1(_05590_),
    .A2(net844),
    .B1(net845),
    .X(_05726_));
 sky130_fd_sc_hd__and3_1 _13454_ (.A(_05699_),
    .B(_05725_),
    .C(_05726_),
    .X(_05727_));
 sky130_fd_sc_hd__a21oi_1 _13455_ (.A1(_05699_),
    .A2(_05726_),
    .B1(_05725_),
    .Y(_05728_));
 sky130_fd_sc_hd__nor2_1 _13456_ (.A(_05727_),
    .B(_05728_),
    .Y(_05729_));
 sky130_fd_sc_hd__clkbuf_1 _13457_ (.A(net1598),
    .X(_05730_));
 sky130_fd_sc_hd__nand2_1 _13458_ (.A(net7747),
    .B(net1313),
    .Y(_05731_));
 sky130_fd_sc_hd__and3_1 _13459_ (.A(net7710),
    .B(net2321),
    .C(net2317),
    .X(_05732_));
 sky130_fd_sc_hd__and3_1 _13460_ (.A(net7722),
    .B(net2331),
    .C(net2325),
    .X(_05733_));
 sky130_fd_sc_hd__xor2_1 _13461_ (.A(_05732_),
    .B(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__xnor2_1 _13462_ (.A(_05731_),
    .B(_05734_),
    .Y(_05735_));
 sky130_fd_sc_hd__a22o_1 _13463_ (.A1(net7705),
    .A2(net1151),
    .B1(_05585_),
    .B2(_05586_),
    .X(_05736_));
 sky130_fd_sc_hd__o21a_1 _13464_ (.A1(_05585_),
    .A2(_05586_),
    .B1(_05736_),
    .X(_05737_));
 sky130_fd_sc_hd__o211a_1 _13465_ (.A1(_05592_),
    .A2(_05593_),
    .B1(net7769),
    .C1(net1313),
    .X(_05738_));
 sky130_fd_sc_hd__a21o_1 _13466_ (.A1(_05592_),
    .A2(_05593_),
    .B1(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__xor2_1 _13467_ (.A(net912),
    .B(net997),
    .X(_05740_));
 sky130_fd_sc_hd__xnor2_1 _13468_ (.A(net998),
    .B(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__o21a_1 _13469_ (.A1(net1131),
    .A2(_05588_),
    .B1(_05581_),
    .X(_05742_));
 sky130_fd_sc_hd__a21oi_2 _13470_ (.A1(net1131),
    .A2(_05588_),
    .B1(_05742_),
    .Y(_05743_));
 sky130_fd_sc_hd__nand2_1 _13471_ (.A(net7685),
    .B(net1151),
    .Y(_05744_));
 sky130_fd_sc_hd__and3_1 _13472_ (.A(net7655),
    .B(net1975),
    .C(net2311),
    .X(_05745_));
 sky130_fd_sc_hd__and3_1 _13473_ (.A(net7671),
    .B(net1982),
    .C(net2360),
    .X(_05746_));
 sky130_fd_sc_hd__xnor2_1 _13474_ (.A(_05745_),
    .B(_05746_),
    .Y(_05747_));
 sky130_fd_sc_hd__xnor2_2 _13475_ (.A(_05744_),
    .B(_05747_),
    .Y(_05748_));
 sky130_fd_sc_hd__a21o_1 _13476_ (.A1(net1574),
    .A2(net1572),
    .B1(net1945),
    .X(_05749_));
 sky130_fd_sc_hd__or2_1 _13477_ (.A(net1574),
    .B(net1572),
    .X(_05750_));
 sky130_fd_sc_hd__and3_1 _13478_ (.A(net7619),
    .B(net1972),
    .C(net1969),
    .X(_05751_));
 sky130_fd_sc_hd__and3_1 _13479_ (.A(net7640),
    .B(net2350),
    .C(net2346),
    .X(_05752_));
 sky130_fd_sc_hd__xor2_1 _13480_ (.A(_05751_),
    .B(_05752_),
    .X(_05753_));
 sky130_fd_sc_hd__a21o_1 _13481_ (.A1(_05749_),
    .A2(_05750_),
    .B1(net1310),
    .X(_05754_));
 sky130_fd_sc_hd__nand3_1 _13482_ (.A(_05749_),
    .B(_05750_),
    .C(net1310),
    .Y(_05755_));
 sky130_fd_sc_hd__nand2_1 _13483_ (.A(_05754_),
    .B(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__xor2_2 _13484_ (.A(_05748_),
    .B(_05756_),
    .X(_05757_));
 sky130_fd_sc_hd__xnor2_1 _13485_ (.A(_05743_),
    .B(_05757_),
    .Y(_05758_));
 sky130_fd_sc_hd__xnor2_1 _13486_ (.A(_05741_),
    .B(_05758_),
    .Y(_05759_));
 sky130_fd_sc_hd__xor2_1 _13487_ (.A(_05729_),
    .B(_05759_),
    .X(_05760_));
 sky130_fd_sc_hd__xnor2_1 _13488_ (.A(_05698_),
    .B(net622),
    .Y(_05761_));
 sky130_fd_sc_hd__xnor2_1 _13489_ (.A(net625),
    .B(_05761_),
    .Y(_05762_));
 sky130_fd_sc_hd__or2b_1 _13490_ (.A(net1130),
    .B_N(_05643_),
    .X(_05763_));
 sky130_fd_sc_hd__clkbuf_1 _13491_ (.A(net1933),
    .X(_05764_));
 sky130_fd_sc_hd__and3_1 _13492_ (.A(net7947),
    .B(net1130),
    .C(net1564),
    .X(_05765_));
 sky130_fd_sc_hd__a31o_1 _13493_ (.A1(_05645_),
    .A2(_05647_),
    .A3(_05763_),
    .B1(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__and2_1 _13494_ (.A(_05636_),
    .B(_05650_),
    .X(_05767_));
 sky130_fd_sc_hd__or2_1 _13495_ (.A(_05636_),
    .B(_05650_),
    .X(_05768_));
 sky130_fd_sc_hd__o21a_1 _13496_ (.A1(net628),
    .A2(_05767_),
    .B1(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__and2b_1 _13497_ (.A_N(net785),
    .B(net578),
    .X(_05770_));
 sky130_fd_sc_hd__and2b_1 _13498_ (.A_N(net578),
    .B(net785),
    .X(_05771_));
 sky130_fd_sc_hd__nor2_1 _13499_ (.A(_05770_),
    .B(_05771_),
    .Y(_05772_));
 sky130_fd_sc_hd__xnor2_2 _13500_ (.A(net534),
    .B(_05772_),
    .Y(_05773_));
 sky130_fd_sc_hd__xnor2_1 _13501_ (.A(net504),
    .B(_05773_),
    .Y(_05774_));
 sky130_fd_sc_hd__xor2_1 _13502_ (.A(net367),
    .B(_05774_),
    .X(_05775_));
 sky130_fd_sc_hd__nor2_1 _13503_ (.A(\svm0.state[1] ),
    .B(\svm0.state[0] ),
    .Y(_05776_));
 sky130_fd_sc_hd__or2_1 _13504_ (.A(net2961),
    .B(net2984),
    .X(_05777_));
 sky130_fd_sc_hd__clkbuf_1 _13505_ (.A(_05777_),
    .X(_00411_));
 sky130_fd_sc_hd__or2_1 _13506_ (.A(_05776_),
    .B(_00411_),
    .X(_05778_));
 sky130_fd_sc_hd__clkbuf_2 _13507_ (.A(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__clkbuf_1 _13508_ (.A(net1308),
    .X(_05780_));
 sky130_fd_sc_hd__a22o_1 _13509_ (.A1(net2374),
    .A2(net324),
    .B1(net1127),
    .B2(net9152),
    .X(_00017_));
 sky130_fd_sc_hd__o21bai_1 _13510_ (.A1(net534),
    .A2(_05770_),
    .B1_N(_05771_),
    .Y(_05781_));
 sky130_fd_sc_hd__a21o_1 _13511_ (.A1(_05698_),
    .A2(net622),
    .B1(net625),
    .X(_05782_));
 sky130_fd_sc_hd__o21a_1 _13512_ (.A1(_05698_),
    .A2(net622),
    .B1(_05782_),
    .X(_05783_));
 sky130_fd_sc_hd__a21o_1 _13513_ (.A1(_05694_),
    .A2(net728),
    .B1(_05693_),
    .X(_05784_));
 sky130_fd_sc_hd__nand2_1 _13514_ (.A(net7786),
    .B(net1586),
    .Y(_05785_));
 sky130_fd_sc_hd__and3_1 _13515_ (.A(net7746),
    .B(net2307),
    .C(net1952),
    .X(_05786_));
 sky130_fd_sc_hd__and3_1 _13516_ (.A(net7770),
    .B(net1942),
    .C(net2291),
    .X(_05787_));
 sky130_fd_sc_hd__xor2_1 _13517_ (.A(_05786_),
    .B(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__xnor2_2 _13518_ (.A(_05785_),
    .B(_05788_),
    .Y(_05789_));
 sky130_fd_sc_hd__o211a_1 _13519_ (.A1(_05701_),
    .A2(_05702_),
    .B1(net7814),
    .C1(net1586),
    .X(_05790_));
 sky130_fd_sc_hd__a21o_1 _13520_ (.A1(_05701_),
    .A2(_05702_),
    .B1(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__nand2_1 _13521_ (.A(net7838),
    .B(net1577),
    .Y(_05792_));
 sky130_fd_sc_hd__and3_1 _13522_ (.A(net7866),
    .B(net2946),
    .C(net1938),
    .X(_05793_));
 sky130_fd_sc_hd__and3_1 _13523_ (.A(net7805),
    .B(net2950),
    .C(net3669),
    .X(_05794_));
 sky130_fd_sc_hd__xor2_1 _13524_ (.A(_05793_),
    .B(_05794_),
    .X(_05795_));
 sky130_fd_sc_hd__xnor2_1 _13525_ (.A(_05792_),
    .B(_05795_),
    .Y(_05796_));
 sky130_fd_sc_hd__xnor2_1 _13526_ (.A(_05791_),
    .B(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__xnor2_2 _13527_ (.A(_05789_),
    .B(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__nor2_1 _13528_ (.A(_05704_),
    .B(net1128),
    .Y(_05799_));
 sky130_fd_sc_hd__a21oi_1 _13529_ (.A1(_05704_),
    .A2(net1128),
    .B1(net1129),
    .Y(_05800_));
 sky130_fd_sc_hd__or2_1 _13530_ (.A(net912),
    .B(net997),
    .X(_05801_));
 sky130_fd_sc_hd__a21o_1 _13531_ (.A1(net912),
    .A2(net997),
    .B1(net998),
    .X(_05802_));
 sky130_fd_sc_hd__o211ai_2 _13532_ (.A1(_05799_),
    .A2(_05800_),
    .B1(_05801_),
    .C1(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__a211o_1 _13533_ (.A1(_05801_),
    .A2(_05802_),
    .B1(_05799_),
    .C1(_05800_),
    .X(_05804_));
 sky130_fd_sc_hd__nand2_1 _13534_ (.A(_05803_),
    .B(_05804_),
    .Y(_05805_));
 sky130_fd_sc_hd__xnor2_2 _13535_ (.A(_05798_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__o21ba_1 _13536_ (.A1(_05743_),
    .A2(_05757_),
    .B1_N(_05741_),
    .X(_05807_));
 sky130_fd_sc_hd__a21o_1 _13537_ (.A1(_05743_),
    .A2(_05757_),
    .B1(_05807_),
    .X(_05808_));
 sky130_fd_sc_hd__nand2_1 _13538_ (.A(net7722),
    .B(net1313),
    .Y(_05809_));
 sky130_fd_sc_hd__and3_1 _13539_ (.A(net7686),
    .B(net2321),
    .C(net2317),
    .X(_05810_));
 sky130_fd_sc_hd__and3_1 _13540_ (.A(net7710),
    .B(net2331),
    .C(net2326),
    .X(_05811_));
 sky130_fd_sc_hd__xor2_1 _13541_ (.A(_05810_),
    .B(_05811_),
    .X(_05812_));
 sky130_fd_sc_hd__xnor2_2 _13542_ (.A(_05809_),
    .B(_05812_),
    .Y(_05813_));
 sky130_fd_sc_hd__a22oi_2 _13543_ (.A1(net7747),
    .A2(net1598),
    .B1(_05732_),
    .B2(_05733_),
    .Y(_05814_));
 sky130_fd_sc_hd__nor2_1 _13544_ (.A(_05732_),
    .B(_05733_),
    .Y(_05815_));
 sky130_fd_sc_hd__a22oi_2 _13545_ (.A1(net7698),
    .A2(net1352),
    .B1(_05745_),
    .B2(_05746_),
    .Y(_05816_));
 sky130_fd_sc_hd__nor2_1 _13546_ (.A(_05745_),
    .B(_05746_),
    .Y(_05817_));
 sky130_fd_sc_hd__nor4_1 _13547_ (.A(_05814_),
    .B(_05815_),
    .C(_05816_),
    .D(_05817_),
    .Y(_05818_));
 sky130_fd_sc_hd__o22a_1 _13548_ (.A1(_05814_),
    .A2(_05815_),
    .B1(_05816_),
    .B2(_05817_),
    .X(_05819_));
 sky130_fd_sc_hd__nor2_1 _13549_ (.A(_05818_),
    .B(_05819_),
    .Y(_05820_));
 sky130_fd_sc_hd__xor2_2 _13550_ (.A(_05813_),
    .B(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__a21bo_1 _13551_ (.A1(_05748_),
    .A2(_05755_),
    .B1_N(_05754_),
    .X(_05822_));
 sky130_fd_sc_hd__and3b_1 _13552_ (.A_N(net1573),
    .B(net1347),
    .C(net7617),
    .X(_05823_));
 sky130_fd_sc_hd__nand2_1 _13553_ (.A(net7671),
    .B(net1150),
    .Y(_05824_));
 sky130_fd_sc_hd__and3_1 _13554_ (.A(net7655),
    .B(net1982),
    .C(net2360),
    .X(_05825_));
 sky130_fd_sc_hd__and3_1 _13555_ (.A(net7638),
    .B(net1975),
    .C(net2311),
    .X(_05826_));
 sky130_fd_sc_hd__xor2_1 _13556_ (.A(_05825_),
    .B(_05826_),
    .X(_05827_));
 sky130_fd_sc_hd__xnor2_1 _13557_ (.A(_05824_),
    .B(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__xnor2_1 _13558_ (.A(_05823_),
    .B(_05828_),
    .Y(_05829_));
 sky130_fd_sc_hd__nor2_1 _13559_ (.A(_05822_),
    .B(_05829_),
    .Y(_05830_));
 sky130_fd_sc_hd__nand2_1 _13560_ (.A(_05822_),
    .B(_05829_),
    .Y(_05831_));
 sky130_fd_sc_hd__or2b_1 _13561_ (.A(_05830_),
    .B_N(_05831_),
    .X(_05832_));
 sky130_fd_sc_hd__xnor2_2 _13562_ (.A(_05821_),
    .B(_05832_),
    .Y(_05833_));
 sky130_fd_sc_hd__xnor2_1 _13563_ (.A(net681),
    .B(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__xnor2_1 _13564_ (.A(_05806_),
    .B(_05834_),
    .Y(_05835_));
 sky130_fd_sc_hd__o21ba_1 _13565_ (.A1(_05728_),
    .A2(_05759_),
    .B1_N(_05727_),
    .X(_05836_));
 sky130_fd_sc_hd__a21o_1 _13566_ (.A1(net7865),
    .A2(net1577),
    .B1(_05710_),
    .X(_05837_));
 sky130_fd_sc_hd__and3_1 _13567_ (.A(net7865),
    .B(net1577),
    .C(_05710_),
    .X(_05838_));
 sky130_fd_sc_hd__a21o_1 _13568_ (.A1(_05708_),
    .A2(_05837_),
    .B1(_05838_),
    .X(_05839_));
 sky130_fd_sc_hd__and3_1 _13569_ (.A(net7895),
    .B(net1928),
    .C(_05839_),
    .X(_05840_));
 sky130_fd_sc_hd__a21o_1 _13570_ (.A1(net7895),
    .A2(net1928),
    .B1(_05839_),
    .X(_05841_));
 sky130_fd_sc_hd__or2b_1 _13571_ (.A(_05840_),
    .B_N(_05841_),
    .X(_05842_));
 sky130_fd_sc_hd__a21o_1 _13572_ (.A1(net916),
    .A2(net913),
    .B1(net915),
    .X(_05843_));
 sky130_fd_sc_hd__o21a_1 _13573_ (.A1(net916),
    .A2(net913),
    .B1(_05843_),
    .X(_05844_));
 sky130_fd_sc_hd__xnor2_2 _13574_ (.A(_05842_),
    .B(net783),
    .Y(_05845_));
 sky130_fd_sc_hd__xor2_1 _13575_ (.A(net679),
    .B(_05845_),
    .X(_05846_));
 sky130_fd_sc_hd__xnor2_1 _13576_ (.A(net577),
    .B(_05846_),
    .Y(_05847_));
 sky130_fd_sc_hd__xnor2_1 _13577_ (.A(_05784_),
    .B(net533),
    .Y(_05848_));
 sky130_fd_sc_hd__xnor2_1 _13578_ (.A(_05783_),
    .B(_05848_),
    .Y(_05849_));
 sky130_fd_sc_hd__or2b_1 _13579_ (.A(_05781_),
    .B_N(_05849_),
    .X(_05850_));
 sky130_fd_sc_hd__or2b_1 _13580_ (.A(_05849_),
    .B_N(_05781_),
    .X(_05851_));
 sky130_fd_sc_hd__nand2_1 _13581_ (.A(_05850_),
    .B(_05851_),
    .Y(_05852_));
 sky130_fd_sc_hd__nor2_1 _13582_ (.A(net504),
    .B(_05773_),
    .Y(_05853_));
 sky130_fd_sc_hd__nand2_1 _13583_ (.A(net504),
    .B(_05773_),
    .Y(_05854_));
 sky130_fd_sc_hd__o21ai_1 _13584_ (.A1(net367),
    .A2(_05853_),
    .B1(_05854_),
    .Y(_05855_));
 sky130_fd_sc_hd__xnor2_1 _13585_ (.A(_05852_),
    .B(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__clkbuf_1 _13586_ (.A(net2371),
    .X(_05857_));
 sky130_fd_sc_hd__a22o_1 _13587_ (.A1(\svm0.tC[1] ),
    .A2(net1127),
    .B1(net287),
    .B2(net1927),
    .X(_00018_));
 sky130_fd_sc_hd__inv_2 _13588_ (.A(net504),
    .Y(_05858_));
 sky130_fd_sc_hd__and2b_1 _13589_ (.A_N(_05771_),
    .B(_05849_),
    .X(_05859_));
 sky130_fd_sc_hd__or3b_1 _13590_ (.A(_05849_),
    .B(_05770_),
    .C_N(net504),
    .X(_05860_));
 sky130_fd_sc_hd__o31a_1 _13591_ (.A1(_05858_),
    .A2(net534),
    .A3(_05859_),
    .B1(_05860_),
    .X(_05861_));
 sky130_fd_sc_hd__o311a_1 _13592_ (.A1(net367),
    .A2(_05774_),
    .A3(_05852_),
    .B1(_05861_),
    .C1(_05851_),
    .X(_05862_));
 sky130_fd_sc_hd__o21ai_1 _13593_ (.A1(_05840_),
    .A2(net783),
    .B1(_05841_),
    .Y(_05863_));
 sky130_fd_sc_hd__o21ba_1 _13594_ (.A1(net577),
    .A2(_05845_),
    .B1_N(net679),
    .X(_05864_));
 sky130_fd_sc_hd__a21oi_1 _13595_ (.A1(net577),
    .A2(_05845_),
    .B1(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__and2_1 _13596_ (.A(_05863_),
    .B(_05865_),
    .X(_05866_));
 sky130_fd_sc_hd__or2_1 _13597_ (.A(_05863_),
    .B(_05865_),
    .X(_05867_));
 sky130_fd_sc_hd__inv_2 _13598_ (.A(_05867_),
    .Y(_05868_));
 sky130_fd_sc_hd__nor2_1 _13599_ (.A(_05866_),
    .B(_05868_),
    .Y(_05869_));
 sky130_fd_sc_hd__nand2_1 _13600_ (.A(_05784_),
    .B(net533),
    .Y(_05870_));
 sky130_fd_sc_hd__nor2_1 _13601_ (.A(_05784_),
    .B(net533),
    .Y(_05871_));
 sky130_fd_sc_hd__a21o_2 _13602_ (.A1(_05783_),
    .A2(_05870_),
    .B1(_05871_),
    .X(_05872_));
 sky130_fd_sc_hd__buf_1 _13603_ (.A(net1589),
    .X(_05873_));
 sky130_fd_sc_hd__nand2_1 _13604_ (.A(net7770),
    .B(net1306),
    .Y(_05874_));
 sky130_fd_sc_hd__and3_1 _13605_ (.A(net7723),
    .B(net2307),
    .C(net1952),
    .X(_05875_));
 sky130_fd_sc_hd__and3_1 _13606_ (.A(net7746),
    .B(net1942),
    .C(net2291),
    .X(_05876_));
 sky130_fd_sc_hd__xnor2_1 _13607_ (.A(_05875_),
    .B(_05876_),
    .Y(_05877_));
 sky130_fd_sc_hd__xnor2_1 _13608_ (.A(_05874_),
    .B(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__a22oi_2 _13609_ (.A1(net7792),
    .A2(net1306),
    .B1(_05786_),
    .B2(_05787_),
    .Y(_05879_));
 sky130_fd_sc_hd__nor2_1 _13610_ (.A(_05786_),
    .B(_05787_),
    .Y(_05880_));
 sky130_fd_sc_hd__nor2_1 _13611_ (.A(_05879_),
    .B(_05880_),
    .Y(_05881_));
 sky130_fd_sc_hd__and2_1 _13612_ (.A(net7811),
    .B(net1578),
    .X(_05882_));
 sky130_fd_sc_hd__and3_1 _13613_ (.A(net7832),
    .B(net2946),
    .C(net1938),
    .X(_05883_));
 sky130_fd_sc_hd__and3_1 _13614_ (.A(net7790),
    .B(net2950),
    .C(net3669),
    .X(_05884_));
 sky130_fd_sc_hd__xor2_1 _13615_ (.A(_05883_),
    .B(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__xnor2_1 _13616_ (.A(_05882_),
    .B(_05885_),
    .Y(_05886_));
 sky130_fd_sc_hd__xnor2_1 _13617_ (.A(_05881_),
    .B(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__xnor2_1 _13618_ (.A(_05878_),
    .B(_05887_),
    .Y(_05888_));
 sky130_fd_sc_hd__or2_1 _13619_ (.A(_05791_),
    .B(_05796_),
    .X(_05889_));
 sky130_fd_sc_hd__o21ba_1 _13620_ (.A1(_05813_),
    .A2(_05818_),
    .B1_N(_05819_),
    .X(_05890_));
 sky130_fd_sc_hd__a21o_1 _13621_ (.A1(_05791_),
    .A2(_05796_),
    .B1(_05789_),
    .X(_05891_));
 sky130_fd_sc_hd__and3_1 _13622_ (.A(_05889_),
    .B(net911),
    .C(_05891_),
    .X(_05892_));
 sky130_fd_sc_hd__a21o_1 _13623_ (.A1(_05889_),
    .A2(_05891_),
    .B1(net911),
    .X(_05893_));
 sky130_fd_sc_hd__and2b_1 _13624_ (.A_N(_05892_),
    .B(_05893_),
    .X(_05894_));
 sky130_fd_sc_hd__xnor2_1 _13625_ (.A(_05888_),
    .B(_05894_),
    .Y(_05895_));
 sky130_fd_sc_hd__and3_1 _13626_ (.A(net7675),
    .B(net2322),
    .C(net2318),
    .X(_05896_));
 sky130_fd_sc_hd__and3_1 _13627_ (.A(net7709),
    .B(net3685),
    .C(net2967),
    .X(_05897_));
 sky130_fd_sc_hd__and3_1 _13628_ (.A(net7686),
    .B(net2331),
    .C(net2326),
    .X(_05898_));
 sky130_fd_sc_hd__xnor2_1 _13629_ (.A(_05897_),
    .B(_05898_),
    .Y(_05899_));
 sky130_fd_sc_hd__xnor2_2 _13630_ (.A(_05896_),
    .B(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__o211a_1 _13631_ (.A1(_05810_),
    .A2(_05811_),
    .B1(net7722),
    .C1(net1598),
    .X(_05901_));
 sky130_fd_sc_hd__a21o_1 _13632_ (.A1(_05810_),
    .A2(_05811_),
    .B1(_05901_),
    .X(_05902_));
 sky130_fd_sc_hd__o211a_1 _13633_ (.A1(_05825_),
    .A2(_05826_),
    .B1(net7671),
    .C1(net1150),
    .X(_05903_));
 sky130_fd_sc_hd__a21o_1 _13634_ (.A1(_05825_),
    .A2(_05826_),
    .B1(_05903_),
    .X(_05904_));
 sky130_fd_sc_hd__xnor2_1 _13635_ (.A(_05902_),
    .B(_05904_),
    .Y(_05905_));
 sky130_fd_sc_hd__xnor2_1 _13636_ (.A(_05900_),
    .B(_05905_),
    .Y(_05906_));
 sky130_fd_sc_hd__nand2_1 _13637_ (.A(net7657),
    .B(net1150),
    .Y(_05907_));
 sky130_fd_sc_hd__nand2_1 _13638_ (.A(net7616),
    .B(net1337),
    .Y(_05908_));
 sky130_fd_sc_hd__and3_1 _13639_ (.A(net7638),
    .B(net1982),
    .C(net2360),
    .X(_05909_));
 sky130_fd_sc_hd__xnor2_1 _13640_ (.A(_05908_),
    .B(_05909_),
    .Y(_05910_));
 sky130_fd_sc_hd__xnor2_1 _13641_ (.A(_05907_),
    .B(_05910_),
    .Y(_05911_));
 sky130_fd_sc_hd__o211a_1 _13642_ (.A1(net1573),
    .A2(_05828_),
    .B1(net7617),
    .C1(net1347),
    .X(_05912_));
 sky130_fd_sc_hd__xnor2_1 _13643_ (.A(_05911_),
    .B(_05912_),
    .Y(_05913_));
 sky130_fd_sc_hd__xnor2_1 _13644_ (.A(_05906_),
    .B(_05913_),
    .Y(_05914_));
 sky130_fd_sc_hd__a21o_1 _13645_ (.A1(_05821_),
    .A2(_05831_),
    .B1(_05830_),
    .X(_05915_));
 sky130_fd_sc_hd__nor2_1 _13646_ (.A(_05914_),
    .B(_05915_),
    .Y(_05916_));
 sky130_fd_sc_hd__nand2_1 _13647_ (.A(_05914_),
    .B(_05915_),
    .Y(_05917_));
 sky130_fd_sc_hd__and2b_1 _13648_ (.A_N(_05916_),
    .B(_05917_),
    .X(_05918_));
 sky130_fd_sc_hd__xnor2_1 _13649_ (.A(_05895_),
    .B(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__nand2_1 _13650_ (.A(_05798_),
    .B(_05804_),
    .Y(_05920_));
 sky130_fd_sc_hd__nand2_2 _13651_ (.A(_05803_),
    .B(_05920_),
    .Y(_05921_));
 sky130_fd_sc_hd__a21o_1 _13652_ (.A1(net7832),
    .A2(net1328),
    .B1(_05794_),
    .X(_05922_));
 sky130_fd_sc_hd__and3_1 _13653_ (.A(net7832),
    .B(net1328),
    .C(_05794_),
    .X(_05923_));
 sky130_fd_sc_hd__a21o_1 _13654_ (.A1(_05793_),
    .A2(_05922_),
    .B1(_05923_),
    .X(_05924_));
 sky130_fd_sc_hd__nand2_1 _13655_ (.A(net7866),
    .B(net1928),
    .Y(_05925_));
 sky130_fd_sc_hd__xnor2_1 _13656_ (.A(_05924_),
    .B(_05925_),
    .Y(_05926_));
 sky130_fd_sc_hd__xnor2_2 _13657_ (.A(_05921_),
    .B(_05926_),
    .Y(_05927_));
 sky130_fd_sc_hd__a21o_1 _13658_ (.A1(_05806_),
    .A2(_05833_),
    .B1(net681),
    .X(_05928_));
 sky130_fd_sc_hd__o21ai_2 _13659_ (.A1(_05806_),
    .A2(_05833_),
    .B1(_05928_),
    .Y(_05929_));
 sky130_fd_sc_hd__nand2_1 _13660_ (.A(_05927_),
    .B(_05929_),
    .Y(_05930_));
 sky130_fd_sc_hd__or2_1 _13661_ (.A(_05927_),
    .B(_05929_),
    .X(_05931_));
 sky130_fd_sc_hd__and2_1 _13662_ (.A(_05930_),
    .B(_05931_),
    .X(_05932_));
 sky130_fd_sc_hd__xnor2_1 _13663_ (.A(_05919_),
    .B(_05932_),
    .Y(_05933_));
 sky130_fd_sc_hd__xor2_1 _13664_ (.A(_05872_),
    .B(net451),
    .X(_05934_));
 sky130_fd_sc_hd__xor2_1 _13665_ (.A(_05869_),
    .B(_05934_),
    .X(_05935_));
 sky130_fd_sc_hd__xnor2_1 _13666_ (.A(net322),
    .B(_05935_),
    .Y(_05936_));
 sky130_fd_sc_hd__a22o_1 _13667_ (.A1(net9149),
    .A2(net1127),
    .B1(net284),
    .B2(net1927),
    .X(_00019_));
 sky130_fd_sc_hd__o21a_1 _13668_ (.A1(_05895_),
    .A2(_05916_),
    .B1(_05917_),
    .X(_05937_));
 sky130_fd_sc_hd__nand2_1 _13669_ (.A(net7746),
    .B(net1306),
    .Y(_05938_));
 sky130_fd_sc_hd__and3_2 _13670_ (.A(net7700),
    .B(net2308),
    .C(net1953),
    .X(_05939_));
 sky130_fd_sc_hd__and3_2 _13671_ (.A(net7717),
    .B(net1943),
    .C(net2292),
    .X(_05940_));
 sky130_fd_sc_hd__xor2_2 _13672_ (.A(_05939_),
    .B(_05940_),
    .X(_05941_));
 sky130_fd_sc_hd__xnor2_2 _13673_ (.A(_05938_),
    .B(_05941_),
    .Y(_05942_));
 sky130_fd_sc_hd__a22o_1 _13674_ (.A1(net7770),
    .A2(net1306),
    .B1(_05875_),
    .B2(_05876_),
    .X(_05943_));
 sky130_fd_sc_hd__or2_1 _13675_ (.A(_05875_),
    .B(_05876_),
    .X(_05944_));
 sky130_fd_sc_hd__nand2_1 _13676_ (.A(_05943_),
    .B(_05944_),
    .Y(_05945_));
 sky130_fd_sc_hd__nor3b_1 _13677_ (.A(net2300),
    .B(net2296),
    .C_N(net7789),
    .Y(_05946_));
 sky130_fd_sc_hd__nand2_1 _13678_ (.A(net7768),
    .B(net3670),
    .Y(_05947_));
 sky130_fd_sc_hd__o2111a_1 _13679_ (.A1(net3677),
    .A2(_05947_),
    .B1(net2947),
    .C1(net7810),
    .D1(net1939),
    .X(_05948_));
 sky130_fd_sc_hd__a311oi_1 _13680_ (.A1(net7810),
    .A2(net2947),
    .A3(net1939),
    .B1(_05947_),
    .C1(net3677),
    .Y(_05949_));
 sky130_fd_sc_hd__or3_1 _13681_ (.A(net1923),
    .B(_05948_),
    .C(_05949_),
    .X(_05950_));
 sky130_fd_sc_hd__o21ai_1 _13682_ (.A1(_05948_),
    .A2(_05949_),
    .B1(net1923),
    .Y(_05951_));
 sky130_fd_sc_hd__and2_1 _13683_ (.A(_05950_),
    .B(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__xnor2_1 _13684_ (.A(_05945_),
    .B(_05952_),
    .Y(_05953_));
 sky130_fd_sc_hd__xnor2_2 _13685_ (.A(_05942_),
    .B(_05953_),
    .Y(_05954_));
 sky130_fd_sc_hd__or3_1 _13686_ (.A(_05879_),
    .B(_05880_),
    .C(_05886_),
    .X(_05955_));
 sky130_fd_sc_hd__and2b_1 _13687_ (.A_N(_05881_),
    .B(_05886_),
    .X(_05956_));
 sky130_fd_sc_hd__a21o_1 _13688_ (.A1(_05878_),
    .A2(_05955_),
    .B1(_05956_),
    .X(_05957_));
 sky130_fd_sc_hd__o21a_1 _13689_ (.A1(_05900_),
    .A2(_05902_),
    .B1(_05904_),
    .X(_05958_));
 sky130_fd_sc_hd__a21o_1 _13690_ (.A1(_05900_),
    .A2(_05902_),
    .B1(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__xor2_1 _13691_ (.A(_05957_),
    .B(net782),
    .X(_05960_));
 sky130_fd_sc_hd__xnor2_1 _13692_ (.A(_05954_),
    .B(_05960_),
    .Y(_05961_));
 sky130_fd_sc_hd__nand2_1 _13693_ (.A(net7621),
    .B(net1605),
    .Y(_05962_));
 sky130_fd_sc_hd__nand2_1 _13694_ (.A(net7637),
    .B(net1149),
    .Y(_05963_));
 sky130_fd_sc_hd__xnor2_1 _13695_ (.A(_05962_),
    .B(_05963_),
    .Y(_05964_));
 sky130_fd_sc_hd__a21oi_1 _13696_ (.A1(_05896_),
    .A2(_05898_),
    .B1(_05897_),
    .Y(_05965_));
 sky130_fd_sc_hd__nor2_1 _13697_ (.A(_05896_),
    .B(_05898_),
    .Y(_05966_));
 sky130_fd_sc_hd__nor2_1 _13698_ (.A(_05965_),
    .B(_05966_),
    .Y(_05967_));
 sky130_fd_sc_hd__a32oi_4 _13699_ (.A1(net7615),
    .A2(net1338),
    .A3(net1563),
    .B1(net1148),
    .B2(net7654),
    .Y(_05968_));
 sky130_fd_sc_hd__a21oi_1 _13700_ (.A1(net7615),
    .A2(net1338),
    .B1(net1563),
    .Y(_05969_));
 sky130_fd_sc_hd__nor2_1 _13701_ (.A(_05968_),
    .B(_05969_),
    .Y(_05970_));
 sky130_fd_sc_hd__xnor2_1 _13702_ (.A(_05967_),
    .B(_05970_),
    .Y(_05971_));
 sky130_fd_sc_hd__inv_2 _13703_ (.A(net7647),
    .Y(_05972_));
 sky130_fd_sc_hd__nor2_1 _13704_ (.A(net4248),
    .B(net1961),
    .Y(_05973_));
 sky130_fd_sc_hd__and3_1 _13705_ (.A(net7697),
    .B(net3685),
    .C(net2967),
    .X(_05974_));
 sky130_fd_sc_hd__and3_1 _13706_ (.A(net7660),
    .B(net2332),
    .C(net2326),
    .X(_05975_));
 sky130_fd_sc_hd__xor2_1 _13707_ (.A(_05974_),
    .B(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__xnor2_1 _13708_ (.A(net1562),
    .B(_05976_),
    .Y(_05977_));
 sky130_fd_sc_hd__xnor2_1 _13709_ (.A(_05971_),
    .B(_05977_),
    .Y(_05978_));
 sky130_fd_sc_hd__xnor2_2 _13710_ (.A(net909),
    .B(net781),
    .Y(_05979_));
 sky130_fd_sc_hd__and2_1 _13711_ (.A(_05911_),
    .B(_05912_),
    .X(_05980_));
 sky130_fd_sc_hd__or2_1 _13712_ (.A(_05911_),
    .B(_05912_),
    .X(_05981_));
 sky130_fd_sc_hd__o21ai_1 _13713_ (.A1(_05906_),
    .A2(_05980_),
    .B1(_05981_),
    .Y(_05982_));
 sky130_fd_sc_hd__xnor2_1 _13714_ (.A(_05979_),
    .B(net727),
    .Y(_05983_));
 sky130_fd_sc_hd__xnor2_1 _13715_ (.A(_05961_),
    .B(_05983_),
    .Y(_05984_));
 sky130_fd_sc_hd__o21a_1 _13716_ (.A1(_05888_),
    .A2(_05892_),
    .B1(_05893_),
    .X(_05985_));
 sky130_fd_sc_hd__a22o_1 _13717_ (.A1(net7831),
    .A2(net1317),
    .B1(_05882_),
    .B2(_05884_),
    .X(_05986_));
 sky130_fd_sc_hd__o21a_1 _13718_ (.A1(_05882_),
    .A2(_05884_),
    .B1(_05986_),
    .X(_05987_));
 sky130_fd_sc_hd__nand2_1 _13719_ (.A(net7831),
    .B(net1929),
    .Y(_05988_));
 sky130_fd_sc_hd__xnor2_1 _13720_ (.A(_05987_),
    .B(_05988_),
    .Y(_05989_));
 sky130_fd_sc_hd__xnor2_2 _13721_ (.A(net780),
    .B(_05989_),
    .Y(_05990_));
 sky130_fd_sc_hd__xnor2_1 _13722_ (.A(_05984_),
    .B(_05990_),
    .Y(_05991_));
 sky130_fd_sc_hd__xnor2_1 _13723_ (.A(net621),
    .B(_05991_),
    .Y(_05992_));
 sky130_fd_sc_hd__or2_1 _13724_ (.A(_05921_),
    .B(_05924_),
    .X(_05993_));
 sky130_fd_sc_hd__nand2_1 _13725_ (.A(_05925_),
    .B(_05929_),
    .Y(_05994_));
 sky130_fd_sc_hd__o21ba_1 _13726_ (.A1(_05921_),
    .A2(_05924_),
    .B1_N(_05925_),
    .X(_05995_));
 sky130_fd_sc_hd__a21oi_1 _13727_ (.A1(_05921_),
    .A2(_05924_),
    .B1(_05995_),
    .Y(_05996_));
 sky130_fd_sc_hd__and2b_1 _13728_ (.A_N(_05919_),
    .B(_05996_),
    .X(_05997_));
 sky130_fd_sc_hd__a2bb2o_1 _13729_ (.A1_N(_05993_),
    .A2_N(_05994_),
    .B1(_05997_),
    .B2(_05931_),
    .X(_05998_));
 sky130_fd_sc_hd__o21ba_1 _13730_ (.A1(_05927_),
    .A2(_05929_),
    .B1_N(_05919_),
    .X(_05999_));
 sky130_fd_sc_hd__a211o_1 _13731_ (.A1(_05927_),
    .A2(_05929_),
    .B1(_05996_),
    .C1(_05999_),
    .X(_06000_));
 sky130_fd_sc_hd__or2b_1 _13732_ (.A(net503),
    .B_N(_06000_),
    .X(_06001_));
 sky130_fd_sc_hd__xnor2_1 _13733_ (.A(_05992_),
    .B(_06001_),
    .Y(_06002_));
 sky130_fd_sc_hd__a21o_1 _13734_ (.A1(_05867_),
    .A2(net451),
    .B1(_05866_),
    .X(_06003_));
 sky130_fd_sc_hd__or2_1 _13735_ (.A(_05867_),
    .B(net451),
    .X(_06004_));
 sky130_fd_sc_hd__o21a_1 _13736_ (.A1(_05872_),
    .A2(_06003_),
    .B1(_06004_),
    .X(_06005_));
 sky130_fd_sc_hd__nand2_1 _13737_ (.A(_05866_),
    .B(net451),
    .Y(_06006_));
 sky130_fd_sc_hd__a21bo_1 _13738_ (.A1(_05872_),
    .A2(_06003_),
    .B1_N(_06006_),
    .X(_06007_));
 sky130_fd_sc_hd__nand2_1 _13739_ (.A(net322),
    .B(_06007_),
    .Y(_06008_));
 sky130_fd_sc_hd__mux2_1 _13740_ (.A0(_06004_),
    .A1(_06006_),
    .S(_05872_),
    .X(_06009_));
 sky130_fd_sc_hd__o211a_1 _13741_ (.A1(net322),
    .A2(_06005_),
    .B1(_06008_),
    .C1(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__xnor2_1 _13742_ (.A(net404),
    .B(_06010_),
    .Y(_06011_));
 sky130_fd_sc_hd__a22o_1 _13743_ (.A1(net9147),
    .A2(net1126),
    .B1(net223),
    .B2(net1926),
    .X(_00020_));
 sky130_fd_sc_hd__and2_1 _13744_ (.A(_05872_),
    .B(net451),
    .X(_06012_));
 sky130_fd_sc_hd__nor2_1 _13745_ (.A(_05872_),
    .B(net451),
    .Y(_06013_));
 sky130_fd_sc_hd__mux2_1 _13746_ (.A0(_06012_),
    .A1(_06013_),
    .S(net404),
    .X(_06014_));
 sky130_fd_sc_hd__mux2_1 _13747_ (.A0(_05866_),
    .A1(_05868_),
    .S(net404),
    .X(_06015_));
 sky130_fd_sc_hd__a22oi_1 _13748_ (.A1(_05869_),
    .A2(_06014_),
    .B1(_06015_),
    .B2(_05934_),
    .Y(_06016_));
 sky130_fd_sc_hd__or2_1 _13749_ (.A(net404),
    .B(_06003_),
    .X(_06017_));
 sky130_fd_sc_hd__a21bo_1 _13750_ (.A1(_05867_),
    .A2(net404),
    .B1_N(_06013_),
    .X(_06018_));
 sky130_fd_sc_hd__o311a_1 _13751_ (.A1(_05866_),
    .A2(_05872_),
    .A3(net404),
    .B1(_06017_),
    .C1(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__o21ai_1 _13752_ (.A1(_05862_),
    .A2(net321),
    .B1(net320),
    .Y(_06020_));
 sky130_fd_sc_hd__o21ai_1 _13753_ (.A1(_05992_),
    .A2(net503),
    .B1(_06000_),
    .Y(_06021_));
 sky130_fd_sc_hd__or2_1 _13754_ (.A(_05979_),
    .B(net727),
    .X(_06022_));
 sky130_fd_sc_hd__and2_1 _13755_ (.A(_05979_),
    .B(net727),
    .X(_06023_));
 sky130_fd_sc_hd__a21oi_1 _13756_ (.A1(_05961_),
    .A2(_06022_),
    .B1(_06023_),
    .Y(_06024_));
 sky130_fd_sc_hd__nand2_1 _13757_ (.A(_05939_),
    .B(_05940_),
    .Y(_06025_));
 sky130_fd_sc_hd__o211ai_2 _13758_ (.A1(_05939_),
    .A2(_05940_),
    .B1(net7741),
    .C1(net1588),
    .Y(_06026_));
 sky130_fd_sc_hd__or3b_1 _13759_ (.A(net2300),
    .B(net2296),
    .C_N(net7768),
    .X(_06027_));
 sky130_fd_sc_hd__nand2_1 _13760_ (.A(net7741),
    .B(net3670),
    .Y(_06028_));
 sky130_fd_sc_hd__o2111ai_1 _13761_ (.A1(net3676),
    .A2(_06028_),
    .B1(net2948),
    .C1(net7789),
    .D1(net1940),
    .Y(_06029_));
 sky130_fd_sc_hd__a311o_1 _13762_ (.A1(net7789),
    .A2(net2948),
    .A3(net1940),
    .B1(_06028_),
    .C1(net3676),
    .X(_06030_));
 sky130_fd_sc_hd__and3_1 _13763_ (.A(_06027_),
    .B(_06029_),
    .C(_06030_),
    .X(_06031_));
 sky130_fd_sc_hd__a21oi_1 _13764_ (.A1(_06029_),
    .A2(_06030_),
    .B1(_06027_),
    .Y(_06032_));
 sky130_fd_sc_hd__a211o_1 _13765_ (.A1(_06025_),
    .A2(_06026_),
    .B1(_06031_),
    .C1(_06032_),
    .X(_06033_));
 sky130_fd_sc_hd__o211ai_2 _13766_ (.A1(_06031_),
    .A2(_06032_),
    .B1(_06025_),
    .C1(_06026_),
    .Y(_06034_));
 sky130_fd_sc_hd__nand2_1 _13767_ (.A(net7721),
    .B(net1307),
    .Y(_06035_));
 sky130_fd_sc_hd__and3_1 _13768_ (.A(net7696),
    .B(net2308),
    .C(net1953),
    .X(_06036_));
 sky130_fd_sc_hd__and3_1 _13769_ (.A(net7700),
    .B(net1943),
    .C(net2292),
    .X(_06037_));
 sky130_fd_sc_hd__xnor2_1 _13770_ (.A(_06036_),
    .B(_06037_),
    .Y(_06038_));
 sky130_fd_sc_hd__xnor2_1 _13771_ (.A(_06035_),
    .B(_06038_),
    .Y(_06039_));
 sky130_fd_sc_hd__a21oi_1 _13772_ (.A1(_06033_),
    .A2(_06034_),
    .B1(_06039_),
    .Y(_06040_));
 sky130_fd_sc_hd__and3_1 _13773_ (.A(_06039_),
    .B(_06033_),
    .C(_06034_),
    .X(_06041_));
 sky130_fd_sc_hd__or2_1 _13774_ (.A(_06040_),
    .B(_06041_),
    .X(_06042_));
 sky130_fd_sc_hd__or4_1 _13775_ (.A(_05965_),
    .B(_05966_),
    .C(_05968_),
    .D(_05969_),
    .X(_06043_));
 sky130_fd_sc_hd__o22a_1 _13776_ (.A1(_05965_),
    .A2(_05966_),
    .B1(_05968_),
    .B2(_05969_),
    .X(_06044_));
 sky130_fd_sc_hd__a21o_1 _13777_ (.A1(_05977_),
    .A2(_06043_),
    .B1(_06044_),
    .X(_06045_));
 sky130_fd_sc_hd__a22o_1 _13778_ (.A1(_05943_),
    .A2(_05944_),
    .B1(_05950_),
    .B2(_05951_),
    .X(_06046_));
 sky130_fd_sc_hd__and4_1 _13779_ (.A(_05943_),
    .B(_05944_),
    .C(_05950_),
    .D(_05951_),
    .X(_06047_));
 sky130_fd_sc_hd__a21oi_2 _13780_ (.A1(_05942_),
    .A2(_06046_),
    .B1(_06047_),
    .Y(_06048_));
 sky130_fd_sc_hd__xnor2_1 _13781_ (.A(net841),
    .B(_06048_),
    .Y(_06049_));
 sky130_fd_sc_hd__xnor2_2 _13782_ (.A(_06042_),
    .B(_06049_),
    .Y(_06050_));
 sky130_fd_sc_hd__or2_1 _13783_ (.A(net909),
    .B(net781),
    .X(_06051_));
 sky130_fd_sc_hd__nand2_1 _13784_ (.A(net7665),
    .B(net1312),
    .Y(_06052_));
 sky130_fd_sc_hd__and3_1 _13785_ (.A(net7636),
    .B(net2322),
    .C(net2318),
    .X(_06053_));
 sky130_fd_sc_hd__and3_1 _13786_ (.A(net7641),
    .B(net2332),
    .C(net2327),
    .X(_06054_));
 sky130_fd_sc_hd__xnor2_1 _13787_ (.A(_06053_),
    .B(_06054_),
    .Y(_06055_));
 sky130_fd_sc_hd__xnor2_1 _13788_ (.A(_06052_),
    .B(_06055_),
    .Y(_06056_));
 sky130_fd_sc_hd__a31o_1 _13789_ (.A1(net7653),
    .A2(net1962),
    .A3(_05975_),
    .B1(_05974_),
    .X(_06057_));
 sky130_fd_sc_hd__a21o_1 _13790_ (.A1(net7653),
    .A2(net1962),
    .B1(_05975_),
    .X(_06058_));
 sky130_fd_sc_hd__nand2_1 _13791_ (.A(_06057_),
    .B(_06058_),
    .Y(_06059_));
 sky130_fd_sc_hd__xnor2_1 _13792_ (.A(_06056_),
    .B(_06059_),
    .Y(_06060_));
 sky130_fd_sc_hd__nand3b_1 _13793_ (.A_N(net1563),
    .B(net1148),
    .C(net7615),
    .Y(_06061_));
 sky130_fd_sc_hd__xor2_1 _13794_ (.A(_06060_),
    .B(_06061_),
    .X(_06062_));
 sky130_fd_sc_hd__xnor2_1 _13795_ (.A(_06051_),
    .B(net840),
    .Y(_06063_));
 sky130_fd_sc_hd__xnor2_2 _13796_ (.A(_06050_),
    .B(_06063_),
    .Y(_06064_));
 sky130_fd_sc_hd__nor2_1 _13797_ (.A(_05954_),
    .B(_05957_),
    .Y(_06065_));
 sky130_fd_sc_hd__nand2_1 _13798_ (.A(_05954_),
    .B(_05957_),
    .Y(_06066_));
 sky130_fd_sc_hd__o21ai_2 _13799_ (.A1(net782),
    .A2(_06065_),
    .B1(_06066_),
    .Y(_06067_));
 sky130_fd_sc_hd__nor2_1 _13800_ (.A(net3677),
    .B(_05947_),
    .Y(_06068_));
 sky130_fd_sc_hd__a22o_1 _13801_ (.A1(net7810),
    .A2(net1319),
    .B1(net1923),
    .B2(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__o21a_1 _13802_ (.A1(net1923),
    .A2(_06068_),
    .B1(_06069_),
    .X(_06070_));
 sky130_fd_sc_hd__nand2_1 _13803_ (.A(net7807),
    .B(net1568),
    .Y(_06071_));
 sky130_fd_sc_hd__xor2_1 _13804_ (.A(net996),
    .B(_06071_),
    .X(_06072_));
 sky130_fd_sc_hd__xnor2_2 _13805_ (.A(_06067_),
    .B(_06072_),
    .Y(_06073_));
 sky130_fd_sc_hd__xor2_1 _13806_ (.A(_06064_),
    .B(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__xnor2_1 _13807_ (.A(_06024_),
    .B(_06074_),
    .Y(_06075_));
 sky130_fd_sc_hd__o21a_1 _13808_ (.A1(net621),
    .A2(_05990_),
    .B1(_05984_),
    .X(_06076_));
 sky130_fd_sc_hd__a21o_1 _13809_ (.A1(net621),
    .A2(_05990_),
    .B1(_06076_),
    .X(_06077_));
 sky130_fd_sc_hd__a21bo_1 _13810_ (.A1(net780),
    .A2(_05987_),
    .B1_N(_05988_),
    .X(_06078_));
 sky130_fd_sc_hd__o21ai_1 _13811_ (.A1(net780),
    .A2(_05987_),
    .B1(_06078_),
    .Y(_06079_));
 sky130_fd_sc_hd__or2_1 _13812_ (.A(net531),
    .B(net678),
    .X(_06080_));
 sky130_fd_sc_hd__and2_1 _13813_ (.A(net531),
    .B(net678),
    .X(_06081_));
 sky130_fd_sc_hd__inv_2 _13814_ (.A(_06081_),
    .Y(_06082_));
 sky130_fd_sc_hd__nand2_1 _13815_ (.A(_06080_),
    .B(_06082_),
    .Y(_06083_));
 sky130_fd_sc_hd__xor2_1 _13816_ (.A(net532),
    .B(_06083_),
    .X(_06084_));
 sky130_fd_sc_hd__xnor2_1 _13817_ (.A(net449),
    .B(_06084_),
    .Y(_06085_));
 sky130_fd_sc_hd__xnor2_1 _13818_ (.A(net283),
    .B(_06085_),
    .Y(_06086_));
 sky130_fd_sc_hd__a22o_1 _13819_ (.A1(net9137),
    .A2(net1126),
    .B1(net256),
    .B2(net1926),
    .X(_00021_));
 sky130_fd_sc_hd__a21bo_1 _13820_ (.A1(_06064_),
    .A2(_06073_),
    .B1_N(_06024_),
    .X(_06087_));
 sky130_fd_sc_hd__o21ai_1 _13821_ (.A1(_06064_),
    .A2(_06073_),
    .B1(_06087_),
    .Y(_06088_));
 sky130_fd_sc_hd__nor2_1 _13822_ (.A(_06050_),
    .B(net840),
    .Y(_06089_));
 sky130_fd_sc_hd__nand2_1 _13823_ (.A(_06050_),
    .B(net840),
    .Y(_06090_));
 sky130_fd_sc_hd__o21a_1 _13824_ (.A1(_06051_),
    .A2(_06089_),
    .B1(_06090_),
    .X(_06091_));
 sky130_fd_sc_hd__nand2_1 _13825_ (.A(net7708),
    .B(net1307),
    .Y(_06092_));
 sky130_fd_sc_hd__and3_1 _13826_ (.A(net7669),
    .B(net2308),
    .C(net1953),
    .X(_06093_));
 sky130_fd_sc_hd__and3_1 _13827_ (.A(net7679),
    .B(net1943),
    .C(net2292),
    .X(_06094_));
 sky130_fd_sc_hd__xor2_1 _13828_ (.A(_06093_),
    .B(_06094_),
    .X(_06095_));
 sky130_fd_sc_hd__xnor2_2 _13829_ (.A(_06092_),
    .B(_06095_),
    .Y(_06096_));
 sky130_fd_sc_hd__o211a_1 _13830_ (.A1(_06036_),
    .A2(_06037_),
    .B1(net7721),
    .C1(net1307),
    .X(_06097_));
 sky130_fd_sc_hd__a21o_1 _13831_ (.A1(_06036_),
    .A2(_06037_),
    .B1(_06097_),
    .X(_06098_));
 sky130_fd_sc_hd__and2_1 _13832_ (.A(net7744),
    .B(net1580),
    .X(_06099_));
 sky130_fd_sc_hd__and3_1 _13833_ (.A(net7766),
    .B(net2948),
    .C(net1940),
    .X(_06100_));
 sky130_fd_sc_hd__and3_1 _13834_ (.A(net7720),
    .B(net2952),
    .C(net3671),
    .X(_06101_));
 sky130_fd_sc_hd__xnor2_1 _13835_ (.A(_06100_),
    .B(_06101_),
    .Y(_06102_));
 sky130_fd_sc_hd__xnor2_1 _13836_ (.A(_06099_),
    .B(_06102_),
    .Y(_06103_));
 sky130_fd_sc_hd__xnor2_1 _13837_ (.A(_06098_),
    .B(_06103_),
    .Y(_06104_));
 sky130_fd_sc_hd__xnor2_2 _13838_ (.A(_06096_),
    .B(_06104_),
    .Y(_06105_));
 sky130_fd_sc_hd__and3_1 _13839_ (.A(net7615),
    .B(net1148),
    .C(net1563),
    .X(_06106_));
 sky130_fd_sc_hd__nand3_1 _13840_ (.A(_06057_),
    .B(_06058_),
    .C(_06106_),
    .Y(_06107_));
 sky130_fd_sc_hd__a21oi_1 _13841_ (.A1(_06057_),
    .A2(_06058_),
    .B1(_06106_),
    .Y(_06108_));
 sky130_fd_sc_hd__a21o_1 _13842_ (.A1(_06056_),
    .A2(_06107_),
    .B1(_06108_),
    .X(_06109_));
 sky130_fd_sc_hd__a21bo_1 _13843_ (.A1(_06039_),
    .A2(_06033_),
    .B1_N(_06034_),
    .X(_06110_));
 sky130_fd_sc_hd__xnor2_1 _13844_ (.A(net839),
    .B(_06110_),
    .Y(_06111_));
 sky130_fd_sc_hd__xnor2_2 _13845_ (.A(_06105_),
    .B(_06111_),
    .Y(_06112_));
 sky130_fd_sc_hd__inv_2 _13846_ (.A(_06106_),
    .Y(_06113_));
 sky130_fd_sc_hd__mux2_1 _13847_ (.A0(_06061_),
    .A1(_06113_),
    .S(_06060_),
    .X(_06114_));
 sky130_fd_sc_hd__nand2_1 _13848_ (.A(net7641),
    .B(net1311),
    .Y(_06115_));
 sky130_fd_sc_hd__nand2_1 _13849_ (.A(net7610),
    .B(net1962),
    .Y(_06116_));
 sky130_fd_sc_hd__inv_2 _13850_ (.A(net7633),
    .Y(_06117_));
 sky130_fd_sc_hd__nor2_1 _13851_ (.A(_06117_),
    .B(net1950),
    .Y(_06118_));
 sky130_fd_sc_hd__xnor2_1 _13852_ (.A(_06116_),
    .B(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__xnor2_1 _13853_ (.A(_06115_),
    .B(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__o211a_1 _13854_ (.A1(_06053_),
    .A2(_06054_),
    .B1(net7669),
    .C1(net1312),
    .X(_06121_));
 sky130_fd_sc_hd__a21o_1 _13855_ (.A1(_06053_),
    .A2(_06054_),
    .B1(_06121_),
    .X(_06122_));
 sky130_fd_sc_hd__xnor2_1 _13856_ (.A(_06120_),
    .B(_06122_),
    .Y(_06123_));
 sky130_fd_sc_hd__xnor2_1 _13857_ (.A(net837),
    .B(net907),
    .Y(_06124_));
 sky130_fd_sc_hd__xnor2_2 _13858_ (.A(_06112_),
    .B(_06124_),
    .Y(_06125_));
 sky130_fd_sc_hd__nand2_1 _13859_ (.A(net841),
    .B(_06048_),
    .Y(_06126_));
 sky130_fd_sc_hd__nor2_1 _13860_ (.A(net841),
    .B(_06048_),
    .Y(_06127_));
 sky130_fd_sc_hd__a21o_1 _13861_ (.A1(_06042_),
    .A2(_06126_),
    .B1(_06127_),
    .X(_06128_));
 sky130_fd_sc_hd__and2_1 _13862_ (.A(net7767),
    .B(net1579),
    .X(_06129_));
 sky130_fd_sc_hd__nor2_1 _13863_ (.A(net3676),
    .B(_06028_),
    .Y(_06130_));
 sky130_fd_sc_hd__a22o_1 _13864_ (.A1(net7788),
    .A2(net1318),
    .B1(_06129_),
    .B2(_06130_),
    .X(_06131_));
 sky130_fd_sc_hd__o21a_1 _13865_ (.A1(_06129_),
    .A2(_06130_),
    .B1(_06131_),
    .X(_06132_));
 sky130_fd_sc_hd__nand2_1 _13866_ (.A(net7788),
    .B(net1930),
    .Y(_06133_));
 sky130_fd_sc_hd__xor2_1 _13867_ (.A(_06132_),
    .B(_06133_),
    .X(_06134_));
 sky130_fd_sc_hd__xnor2_1 _13868_ (.A(_06128_),
    .B(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__xor2_1 _13869_ (.A(_06125_),
    .B(_06135_),
    .X(_06136_));
 sky130_fd_sc_hd__xnor2_2 _13870_ (.A(_06091_),
    .B(_06136_),
    .Y(_06137_));
 sky130_fd_sc_hd__and2b_1 _13871_ (.A_N(net996),
    .B(_06071_),
    .X(_06138_));
 sky130_fd_sc_hd__nor2_1 _13872_ (.A(_06067_),
    .B(_06138_),
    .Y(_06139_));
 sky130_fd_sc_hd__a31o_1 _13873_ (.A1(net7807),
    .A2(net1568),
    .A3(net996),
    .B1(_06139_),
    .X(_06140_));
 sky130_fd_sc_hd__xor2_1 _13874_ (.A(_06137_),
    .B(_06140_),
    .X(_06141_));
 sky130_fd_sc_hd__xnor2_2 _13875_ (.A(net530),
    .B(_06141_),
    .Y(_06142_));
 sky130_fd_sc_hd__and2_1 _13876_ (.A(net532),
    .B(_06080_),
    .X(_06143_));
 sky130_fd_sc_hd__nor2_1 _13877_ (.A(_06081_),
    .B(_06143_),
    .Y(_06144_));
 sky130_fd_sc_hd__nand2_1 _13878_ (.A(net532),
    .B(_06081_),
    .Y(_06145_));
 sky130_fd_sc_hd__o21a_1 _13879_ (.A1(net449),
    .A2(_06144_),
    .B1(_06145_),
    .X(_06146_));
 sky130_fd_sc_hd__or2_1 _13880_ (.A(net532),
    .B(_06080_),
    .X(_06147_));
 sky130_fd_sc_hd__a21bo_1 _13881_ (.A1(net449),
    .A2(_06144_),
    .B1_N(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__nand2_1 _13882_ (.A(net283),
    .B(_06148_),
    .Y(_06149_));
 sky130_fd_sc_hd__mux2_1 _13883_ (.A0(_06145_),
    .A1(_06147_),
    .S(net449),
    .X(_06150_));
 sky130_fd_sc_hd__o211a_1 _13884_ (.A1(net283),
    .A2(_06146_),
    .B1(_06149_),
    .C1(_06150_),
    .X(_06151_));
 sky130_fd_sc_hd__xnor2_1 _13885_ (.A(_06142_),
    .B(_06151_),
    .Y(_06152_));
 sky130_fd_sc_hd__a22o_1 _13886_ (.A1(net9180),
    .A2(net1126),
    .B1(net191),
    .B2(net1926),
    .X(_00022_));
 sky130_fd_sc_hd__or2_1 _13887_ (.A(_06081_),
    .B(_06143_),
    .X(_06153_));
 sky130_fd_sc_hd__o21a_1 _13888_ (.A1(_06081_),
    .A2(_06142_),
    .B1(net532),
    .X(_06154_));
 sky130_fd_sc_hd__a21oi_1 _13889_ (.A1(_06080_),
    .A2(_06142_),
    .B1(_06154_),
    .Y(_06155_));
 sky130_fd_sc_hd__a2bb2o_1 _13890_ (.A1_N(_06142_),
    .A2_N(_06153_),
    .B1(_06155_),
    .B2(net449),
    .X(_06156_));
 sky130_fd_sc_hd__o2bb2a_1 _13891_ (.A1_N(_06142_),
    .A2_N(_06153_),
    .B1(_06155_),
    .B2(net449),
    .X(_06157_));
 sky130_fd_sc_hd__o21ai_1 _13892_ (.A1(net283),
    .A2(_06156_),
    .B1(_06157_),
    .Y(_06158_));
 sky130_fd_sc_hd__nand2_1 _13893_ (.A(_06137_),
    .B(_06140_),
    .Y(_06159_));
 sky130_fd_sc_hd__nand2_1 _13894_ (.A(_06125_),
    .B(_06135_),
    .Y(_06160_));
 sky130_fd_sc_hd__nor2_1 _13895_ (.A(_06125_),
    .B(_06135_),
    .Y(_06161_));
 sky130_fd_sc_hd__a21oi_1 _13896_ (.A1(_06091_),
    .A2(_06160_),
    .B1(_06161_),
    .Y(_06162_));
 sky130_fd_sc_hd__or2b_1 _13897_ (.A(_06132_),
    .B_N(_06133_),
    .X(_06163_));
 sky130_fd_sc_hd__and3_1 _13898_ (.A(net7788),
    .B(net1568),
    .C(_06132_),
    .X(_06164_));
 sky130_fd_sc_hd__a21oi_2 _13899_ (.A1(_06128_),
    .A2(_06163_),
    .B1(_06164_),
    .Y(_06165_));
 sky130_fd_sc_hd__a21bo_1 _13900_ (.A1(net839),
    .A2(_06110_),
    .B1_N(_06105_),
    .X(_06166_));
 sky130_fd_sc_hd__o21a_1 _13901_ (.A1(net839),
    .A2(_06110_),
    .B1(_06166_),
    .X(_06167_));
 sky130_fd_sc_hd__a31o_1 _13902_ (.A1(net7744),
    .A2(net1326),
    .A3(_06101_),
    .B1(_06100_),
    .X(_06168_));
 sky130_fd_sc_hd__o21a_1 _13903_ (.A1(_06099_),
    .A2(_06101_),
    .B1(_06168_),
    .X(_06169_));
 sky130_fd_sc_hd__nand2_1 _13904_ (.A(net7766),
    .B(net1931),
    .Y(_06170_));
 sky130_fd_sc_hd__xor2_1 _13905_ (.A(_06169_),
    .B(_06170_),
    .X(_06171_));
 sky130_fd_sc_hd__xnor2_2 _13906_ (.A(_06167_),
    .B(_06171_),
    .Y(_06172_));
 sky130_fd_sc_hd__nand2_1 _13907_ (.A(net3686),
    .B(net2968),
    .Y(_06173_));
 sky130_fd_sc_hd__nand2_1 _13908_ (.A(net7633),
    .B(net7605),
    .Y(_06174_));
 sky130_fd_sc_hd__or3_1 _13909_ (.A(_06173_),
    .B(net1950),
    .C(_06174_),
    .X(_06175_));
 sky130_fd_sc_hd__o22a_1 _13910_ (.A1(net7632),
    .A2(net1583),
    .B1(_06175_),
    .B2(net1965),
    .X(_06176_));
 sky130_fd_sc_hd__and2_1 _13911_ (.A(net7632),
    .B(net7611),
    .X(_06177_));
 sky130_fd_sc_hd__and3_1 _13912_ (.A(_06117_),
    .B(net1311),
    .C(net1583),
    .X(_06178_));
 sky130_fd_sc_hd__a21oi_1 _13913_ (.A1(net1950),
    .A2(_06177_),
    .B1(_06178_),
    .Y(_06179_));
 sky130_fd_sc_hd__o22a_1 _13914_ (.A1(_06117_),
    .A2(net1311),
    .B1(_06179_),
    .B2(net4248),
    .X(_06180_));
 sky130_fd_sc_hd__o21a_1 _13915_ (.A1(net1965),
    .A2(net1583),
    .B1(net7611),
    .X(_06181_));
 sky130_fd_sc_hd__o21bai_1 _13916_ (.A1(_06173_),
    .A2(_06054_),
    .B1_N(net7610),
    .Y(_06182_));
 sky130_fd_sc_hd__o221a_1 _13917_ (.A1(net1311),
    .A2(net1583),
    .B1(_06181_),
    .B2(net7633),
    .C1(_06182_),
    .X(_06183_));
 sky130_fd_sc_hd__o221a_1 _13918_ (.A1(net7641),
    .A2(_06176_),
    .B1(_06180_),
    .B2(net1961),
    .C1(_06183_),
    .X(_06184_));
 sky130_fd_sc_hd__nand2_1 _13919_ (.A(net7681),
    .B(_05873_),
    .Y(_06185_));
 sky130_fd_sc_hd__nand2_1 _13920_ (.A(net7645),
    .B(net1331),
    .Y(_06186_));
 sky130_fd_sc_hd__and3_1 _13921_ (.A(net7668),
    .B(net1944),
    .C(net2293),
    .X(_06187_));
 sky130_fd_sc_hd__xnor2_1 _13922_ (.A(_06186_),
    .B(_06187_),
    .Y(_06188_));
 sky130_fd_sc_hd__xnor2_2 _13923_ (.A(_06185_),
    .B(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__o211a_1 _13924_ (.A1(_06093_),
    .A2(_06094_),
    .B1(net7704),
    .C1(net1307),
    .X(_06190_));
 sky130_fd_sc_hd__a21oi_2 _13925_ (.A1(_06093_),
    .A2(_06094_),
    .B1(_06190_),
    .Y(_06191_));
 sky130_fd_sc_hd__and2_1 _13926_ (.A(net7721),
    .B(net1581),
    .X(_06192_));
 sky130_fd_sc_hd__nand2_1 _13927_ (.A(net7743),
    .B(net1571),
    .Y(_06193_));
 sky130_fd_sc_hd__and3_1 _13928_ (.A(net7704),
    .B(net2953),
    .C(net3672),
    .X(_06194_));
 sky130_fd_sc_hd__xnor2_1 _13929_ (.A(_06193_),
    .B(_06194_),
    .Y(_06195_));
 sky130_fd_sc_hd__xnor2_2 _13930_ (.A(_06192_),
    .B(_06195_),
    .Y(_06196_));
 sky130_fd_sc_hd__xnor2_1 _13931_ (.A(_06191_),
    .B(_06196_),
    .Y(_06197_));
 sky130_fd_sc_hd__xnor2_2 _13932_ (.A(_06189_),
    .B(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__nand2_1 _13933_ (.A(_06120_),
    .B(_06122_),
    .Y(_06199_));
 sky130_fd_sc_hd__a21o_1 _13934_ (.A1(_06098_),
    .A2(_06103_),
    .B1(_06096_),
    .X(_06200_));
 sky130_fd_sc_hd__o21a_1 _13935_ (.A1(_06098_),
    .A2(_06103_),
    .B1(_06200_),
    .X(_06201_));
 sky130_fd_sc_hd__xor2_1 _13936_ (.A(net906),
    .B(_06201_),
    .X(_06202_));
 sky130_fd_sc_hd__xnor2_1 _13937_ (.A(_06198_),
    .B(_06202_),
    .Y(_06203_));
 sky130_fd_sc_hd__xnor2_1 _13938_ (.A(net836),
    .B(_06203_),
    .Y(_06204_));
 sky130_fd_sc_hd__xnor2_1 _13939_ (.A(_06172_),
    .B(net677),
    .Y(_06205_));
 sky130_fd_sc_hd__nor2_1 _13940_ (.A(net837),
    .B(net907),
    .Y(_06206_));
 sky130_fd_sc_hd__nand2_1 _13941_ (.A(net837),
    .B(net907),
    .Y(_06207_));
 sky130_fd_sc_hd__o21ai_2 _13942_ (.A1(_06112_),
    .A2(_06206_),
    .B1(_06207_),
    .Y(_06208_));
 sky130_fd_sc_hd__xnor2_2 _13943_ (.A(_06205_),
    .B(_06208_),
    .Y(_06209_));
 sky130_fd_sc_hd__xor2_1 _13944_ (.A(_06165_),
    .B(_06209_),
    .X(_06210_));
 sky130_fd_sc_hd__xnor2_1 _13945_ (.A(_06162_),
    .B(_06210_),
    .Y(_06211_));
 sky130_fd_sc_hd__o21ai_1 _13946_ (.A1(_06137_),
    .A2(_06140_),
    .B1(net530),
    .Y(_06212_));
 sky130_fd_sc_hd__and3_1 _13947_ (.A(_06159_),
    .B(_06211_),
    .C(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__a21o_1 _13948_ (.A1(_06159_),
    .A2(_06212_),
    .B1(_06211_),
    .X(_06214_));
 sky130_fd_sc_hd__and2b_1 _13949_ (.A_N(_06213_),
    .B(_06214_),
    .X(_06215_));
 sky130_fd_sc_hd__xnor2_1 _13950_ (.A(_06158_),
    .B(_06215_),
    .Y(_06216_));
 sky130_fd_sc_hd__a22o_1 _13951_ (.A1(net9118),
    .A2(net1126),
    .B1(net220),
    .B2(net1926),
    .X(_00023_));
 sky130_fd_sc_hd__o21a_1 _13952_ (.A1(_06158_),
    .A2(_06213_),
    .B1(_06214_),
    .X(_06217_));
 sky130_fd_sc_hd__buf_1 _13953_ (.A(_05873_),
    .X(_06218_));
 sky130_fd_sc_hd__nand2_1 _13954_ (.A(net7664),
    .B(net1125),
    .Y(_06219_));
 sky130_fd_sc_hd__nor2_1 _13955_ (.A(_06117_),
    .B(net1597),
    .Y(_06220_));
 sky130_fd_sc_hd__buf_2 _13956_ (.A(_05191_),
    .X(_06221_));
 sky130_fd_sc_hd__nand2_1 _13957_ (.A(net7642),
    .B(_06221_),
    .Y(_06222_));
 sky130_fd_sc_hd__xnor2_1 _13958_ (.A(_06220_),
    .B(_06222_),
    .Y(_06223_));
 sky130_fd_sc_hd__xnor2_2 _13959_ (.A(_06219_),
    .B(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__a21o_1 _13960_ (.A1(net7648),
    .A2(net1331),
    .B1(_06187_),
    .X(_06225_));
 sky130_fd_sc_hd__a32o_1 _13961_ (.A1(net7648),
    .A2(net1331),
    .A3(_06187_),
    .B1(_06218_),
    .B2(net7681),
    .X(_06226_));
 sky130_fd_sc_hd__nand2_1 _13962_ (.A(_06225_),
    .B(_06226_),
    .Y(_06227_));
 sky130_fd_sc_hd__nand2_1 _13963_ (.A(net7703),
    .B(net1324),
    .Y(_06228_));
 sky130_fd_sc_hd__nand2_1 _13964_ (.A(net7718),
    .B(net1571),
    .Y(_06229_));
 sky130_fd_sc_hd__and3_1 _13965_ (.A(net7683),
    .B(net2954),
    .C(net3673),
    .X(_06230_));
 sky130_fd_sc_hd__xor2_1 _13966_ (.A(_06229_),
    .B(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__xnor2_2 _13967_ (.A(_06228_),
    .B(_06231_),
    .Y(_06232_));
 sky130_fd_sc_hd__xnor2_1 _13968_ (.A(_06227_),
    .B(_06232_),
    .Y(_06233_));
 sky130_fd_sc_hd__xnor2_2 _13969_ (.A(_06224_),
    .B(_06233_),
    .Y(_06234_));
 sky130_fd_sc_hd__and2_1 _13970_ (.A(_06117_),
    .B(net7604),
    .X(_06235_));
 sky130_fd_sc_hd__nor2_1 _13971_ (.A(net1961),
    .B(net1583),
    .Y(_06236_));
 sky130_fd_sc_hd__mux2_1 _13972_ (.A0(net1583),
    .A1(_06236_),
    .S(net7601),
    .X(_06237_));
 sky130_fd_sc_hd__a32o_1 _13973_ (.A1(net1965),
    .A2(net1583),
    .A3(_06235_),
    .B1(_06237_),
    .B2(net7633),
    .X(_06238_));
 sky130_fd_sc_hd__and3_1 _13974_ (.A(net7642),
    .B(net1311),
    .C(_06238_),
    .X(_06239_));
 sky130_fd_sc_hd__a41o_1 _13975_ (.A1(_06173_),
    .A2(net1965),
    .A3(net1583),
    .A4(_06177_),
    .B1(_06239_),
    .X(_06240_));
 sky130_fd_sc_hd__a21bo_1 _13976_ (.A1(_06191_),
    .A2(_06196_),
    .B1_N(_06189_),
    .X(_06241_));
 sky130_fd_sc_hd__o21ai_2 _13977_ (.A1(_06191_),
    .A2(_06196_),
    .B1(_06241_),
    .Y(_06242_));
 sky130_fd_sc_hd__xor2_1 _13978_ (.A(net835),
    .B(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__xnor2_1 _13979_ (.A(_06234_),
    .B(_06243_),
    .Y(_06244_));
 sky130_fd_sc_hd__or3b_1 _13980_ (.A(_06118_),
    .B(_06173_),
    .C_N(net7610),
    .X(_06245_));
 sky130_fd_sc_hd__or2_1 _13981_ (.A(_06244_),
    .B(net1305),
    .X(_06246_));
 sky130_fd_sc_hd__nand2_1 _13982_ (.A(_06244_),
    .B(net1305),
    .Y(_06247_));
 sky130_fd_sc_hd__and2_1 _13983_ (.A(_06246_),
    .B(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__and2_1 _13984_ (.A(net836),
    .B(_06203_),
    .X(_06249_));
 sky130_fd_sc_hd__a21bo_1 _13985_ (.A1(_06201_),
    .A2(_06198_),
    .B1_N(net906),
    .X(_06250_));
 sky130_fd_sc_hd__o21ai_1 _13986_ (.A1(_06201_),
    .A2(_06198_),
    .B1(_06250_),
    .Y(_06251_));
 sky130_fd_sc_hd__a21bo_1 _13987_ (.A1(_06192_),
    .A2(_06194_),
    .B1_N(_06193_),
    .X(_06252_));
 sky130_fd_sc_hd__o21a_1 _13988_ (.A1(_06192_),
    .A2(_06194_),
    .B1(_06252_),
    .X(_06253_));
 sky130_fd_sc_hd__nand2_1 _13989_ (.A(net7743),
    .B(net1570),
    .Y(_06254_));
 sky130_fd_sc_hd__xnor2_1 _13990_ (.A(_06253_),
    .B(_06254_),
    .Y(_06255_));
 sky130_fd_sc_hd__xnor2_1 _13991_ (.A(_06251_),
    .B(_06255_),
    .Y(_06256_));
 sky130_fd_sc_hd__xor2_1 _13992_ (.A(_06249_),
    .B(_06256_),
    .X(_06257_));
 sky130_fd_sc_hd__xnor2_1 _13993_ (.A(_06248_),
    .B(_06257_),
    .Y(_06258_));
 sky130_fd_sc_hd__a21o_1 _13994_ (.A1(_06172_),
    .A2(net677),
    .B1(_06208_),
    .X(_06259_));
 sky130_fd_sc_hd__o21ai_2 _13995_ (.A1(_06172_),
    .A2(net677),
    .B1(_06259_),
    .Y(_06260_));
 sky130_fd_sc_hd__and2b_1 _13996_ (.A_N(_06169_),
    .B(_06170_),
    .X(_06261_));
 sky130_fd_sc_hd__and3_1 _13997_ (.A(net7766),
    .B(net1569),
    .C(_06169_),
    .X(_06262_));
 sky130_fd_sc_hd__o21ba_1 _13998_ (.A1(_06167_),
    .A2(_06261_),
    .B1_N(_06262_),
    .X(_06263_));
 sky130_fd_sc_hd__xnor2_1 _13999_ (.A(_06260_),
    .B(_06263_),
    .Y(_06264_));
 sky130_fd_sc_hd__xnor2_2 _14000_ (.A(net529),
    .B(_06264_),
    .Y(_06265_));
 sky130_fd_sc_hd__nor2_1 _14001_ (.A(_06165_),
    .B(_06209_),
    .Y(_06266_));
 sky130_fd_sc_hd__nand2_1 _14002_ (.A(_06165_),
    .B(_06209_),
    .Y(_06267_));
 sky130_fd_sc_hd__o21a_1 _14003_ (.A1(_06162_),
    .A2(_06266_),
    .B1(_06267_),
    .X(_06268_));
 sky130_fd_sc_hd__xor2_1 _14004_ (.A(_06265_),
    .B(_06268_),
    .X(_06269_));
 sky130_fd_sc_hd__xnor2_1 _14005_ (.A(_06217_),
    .B(_06269_),
    .Y(_06270_));
 sky130_fd_sc_hd__a22o_1 _14006_ (.A1(\svm0.tC[7] ),
    .A2(net1126),
    .B1(net189),
    .B2(net1926),
    .X(_00024_));
 sky130_fd_sc_hd__nand2_1 _14007_ (.A(_06265_),
    .B(_06268_),
    .Y(_06271_));
 sky130_fd_sc_hd__nor2_1 _14008_ (.A(_06265_),
    .B(_06268_),
    .Y(_06272_));
 sky130_fd_sc_hd__a21oi_1 _14009_ (.A1(_06214_),
    .A2(_06271_),
    .B1(_06272_),
    .Y(_06273_));
 sky130_fd_sc_hd__nor2_1 _14010_ (.A(_06156_),
    .B(_06273_),
    .Y(_06274_));
 sky130_fd_sc_hd__o211ai_1 _14011_ (.A1(_05862_),
    .A2(net321),
    .B1(net320),
    .C1(_06274_),
    .Y(_06275_));
 sky130_fd_sc_hd__a31o_1 _14012_ (.A1(_06157_),
    .A2(_06215_),
    .A3(_06269_),
    .B1(_06273_),
    .X(_06276_));
 sky130_fd_sc_hd__nand2_1 _14013_ (.A(net282),
    .B(net319),
    .Y(_06277_));
 sky130_fd_sc_hd__inv_2 _14014_ (.A(_06260_),
    .Y(_06278_));
 sky130_fd_sc_hd__a21o_1 _14015_ (.A1(_06278_),
    .A2(_06263_),
    .B1(net529),
    .X(_06279_));
 sky130_fd_sc_hd__o21ai_1 _14016_ (.A1(_06278_),
    .A2(_06263_),
    .B1(_06279_),
    .Y(_06280_));
 sky130_fd_sc_hd__a31o_1 _14017_ (.A1(_06246_),
    .A2(_06247_),
    .A3(_06256_),
    .B1(_06249_),
    .X(_06281_));
 sky130_fd_sc_hd__o21a_1 _14018_ (.A1(_06248_),
    .A2(_06256_),
    .B1(_06281_),
    .X(_06282_));
 sky130_fd_sc_hd__o21a_1 _14019_ (.A1(_06234_),
    .A2(_06242_),
    .B1(net835),
    .X(_06283_));
 sky130_fd_sc_hd__a21o_1 _14020_ (.A1(_06234_),
    .A2(_06242_),
    .B1(_06283_),
    .X(_06284_));
 sky130_fd_sc_hd__a32o_1 _14021_ (.A1(net7702),
    .A2(net1324),
    .A3(_06230_),
    .B1(net1316),
    .B2(net7718),
    .X(_06285_));
 sky130_fd_sc_hd__a21o_1 _14022_ (.A1(net7702),
    .A2(net1324),
    .B1(_06230_),
    .X(_06286_));
 sky130_fd_sc_hd__and2_1 _14023_ (.A(_06285_),
    .B(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__nand2_1 _14024_ (.A(net7718),
    .B(net1567),
    .Y(_06288_));
 sky130_fd_sc_hd__xor2_1 _14025_ (.A(_06287_),
    .B(_06288_),
    .X(_06289_));
 sky130_fd_sc_hd__xnor2_2 _14026_ (.A(_06284_),
    .B(_06289_),
    .Y(_06290_));
 sky130_fd_sc_hd__nand2_1 _14027_ (.A(net7646),
    .B(net1124),
    .Y(_06291_));
 sky130_fd_sc_hd__and3_1 _14028_ (.A(net7625),
    .B(_05608_),
    .C(_05609_),
    .X(_06292_));
 sky130_fd_sc_hd__xor2_2 _14029_ (.A(_06291_),
    .B(net1560),
    .X(_06293_));
 sky130_fd_sc_hd__nand2_1 _14030_ (.A(net7604),
    .B(net1332),
    .Y(_06294_));
 sky130_fd_sc_hd__xnor2_2 _14031_ (.A(_06293_),
    .B(_06294_),
    .Y(_06295_));
 sky130_fd_sc_hd__and3_1 _14032_ (.A(net7642),
    .B(_05608_),
    .C(_05609_),
    .X(_06296_));
 sky130_fd_sc_hd__a21bo_1 _14033_ (.A1(_06220_),
    .A2(_06296_),
    .B1_N(_06219_),
    .X(_06297_));
 sky130_fd_sc_hd__o21a_1 _14034_ (.A1(_06220_),
    .A2(_06296_),
    .B1(_06297_),
    .X(_06298_));
 sky130_fd_sc_hd__nand2_1 _14035_ (.A(net7680),
    .B(net1323),
    .Y(_06299_));
 sky130_fd_sc_hd__nand2_1 _14036_ (.A(net7706),
    .B(net1315),
    .Y(_06300_));
 sky130_fd_sc_hd__and3_1 _14037_ (.A(net7663),
    .B(net2955),
    .C(net3674),
    .X(_06301_));
 sky130_fd_sc_hd__xnor2_1 _14038_ (.A(_06300_),
    .B(_06301_),
    .Y(_06302_));
 sky130_fd_sc_hd__xnor2_2 _14039_ (.A(_06299_),
    .B(_06302_),
    .Y(_06303_));
 sky130_fd_sc_hd__xor2_1 _14040_ (.A(_06298_),
    .B(_06303_),
    .X(_06304_));
 sky130_fd_sc_hd__xnor2_2 _14041_ (.A(_06295_),
    .B(_06304_),
    .Y(_06305_));
 sky130_fd_sc_hd__o21ba_1 _14042_ (.A1(_06227_),
    .A2(_06232_),
    .B1_N(_06224_),
    .X(_06306_));
 sky130_fd_sc_hd__a21oi_2 _14043_ (.A1(_06227_),
    .A2(_06232_),
    .B1(_06306_),
    .Y(_06307_));
 sky130_fd_sc_hd__xor2_1 _14044_ (.A(net1561),
    .B(_06307_),
    .X(_06308_));
 sky130_fd_sc_hd__xnor2_2 _14045_ (.A(_06305_),
    .B(_06308_),
    .Y(_06309_));
 sky130_fd_sc_hd__xnor2_1 _14046_ (.A(_06246_),
    .B(_06309_),
    .Y(_06310_));
 sky130_fd_sc_hd__xnor2_1 _14047_ (.A(_06290_),
    .B(_06310_),
    .Y(_06311_));
 sky130_fd_sc_hd__and2b_1 _14048_ (.A_N(_06253_),
    .B(_06254_),
    .X(_06312_));
 sky130_fd_sc_hd__and3_1 _14049_ (.A(net7742),
    .B(net1570),
    .C(_06253_),
    .X(_06313_));
 sky130_fd_sc_hd__o21ba_1 _14050_ (.A1(_06251_),
    .A2(_06312_),
    .B1_N(_06313_),
    .X(_06314_));
 sky130_fd_sc_hd__nand2_1 _14051_ (.A(_06311_),
    .B(_06314_),
    .Y(_06315_));
 sky130_fd_sc_hd__inv_2 _14052_ (.A(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__nor2_1 _14053_ (.A(_06311_),
    .B(_06314_),
    .Y(_06317_));
 sky130_fd_sc_hd__nor2_1 _14054_ (.A(_06316_),
    .B(_06317_),
    .Y(_06318_));
 sky130_fd_sc_hd__xnor2_1 _14055_ (.A(_06282_),
    .B(_06318_),
    .Y(_06319_));
 sky130_fd_sc_hd__xnor2_1 _14056_ (.A(_06280_),
    .B(net366),
    .Y(_06320_));
 sky130_fd_sc_hd__xnor2_1 _14057_ (.A(_06277_),
    .B(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__a22o_1 _14058_ (.A1(net9161),
    .A2(net1127),
    .B1(net219),
    .B2(net1927),
    .X(_00025_));
 sky130_fd_sc_hd__a21bo_1 _14059_ (.A1(_06290_),
    .A2(_06309_),
    .B1_N(_06246_),
    .X(_06322_));
 sky130_fd_sc_hd__o21ai_4 _14060_ (.A1(_06290_),
    .A2(_06309_),
    .B1(_06322_),
    .Y(_06323_));
 sky130_fd_sc_hd__a21bo_1 _14061_ (.A1(_06307_),
    .A2(_06305_),
    .B1_N(net1561),
    .X(_06324_));
 sky130_fd_sc_hd__o21a_1 _14062_ (.A1(_06307_),
    .A2(_06305_),
    .B1(_06324_),
    .X(_06325_));
 sky130_fd_sc_hd__clkbuf_1 _14063_ (.A(net1322),
    .X(_06326_));
 sky130_fd_sc_hd__a32o_1 _14064_ (.A1(net7680),
    .A2(net1122),
    .A3(_06301_),
    .B1(net1315),
    .B2(net7706),
    .X(_06327_));
 sky130_fd_sc_hd__a21o_1 _14065_ (.A1(net7680),
    .A2(net1122),
    .B1(_06301_),
    .X(_06328_));
 sky130_fd_sc_hd__and2_1 _14066_ (.A(_06327_),
    .B(_06328_),
    .X(_06329_));
 sky130_fd_sc_hd__nand2_1 _14067_ (.A(net7701),
    .B(net1567),
    .Y(_06330_));
 sky130_fd_sc_hd__xnor2_1 _14068_ (.A(_06329_),
    .B(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__xnor2_2 _14069_ (.A(_06325_),
    .B(_06331_),
    .Y(_06332_));
 sky130_fd_sc_hd__nand2_1 _14070_ (.A(_06221_),
    .B(net1125),
    .Y(_06333_));
 sky130_fd_sc_hd__o22a_1 _14071_ (.A1(_06221_),
    .A2(_06174_),
    .B1(_06333_),
    .B2(net7625),
    .X(_06334_));
 sky130_fd_sc_hd__o22a_1 _14072_ (.A1(_06117_),
    .A2(net1125),
    .B1(_06334_),
    .B2(net4249),
    .X(_06335_));
 sky130_fd_sc_hd__o32a_1 _14073_ (.A1(net1332),
    .A2(_06174_),
    .A3(_06333_),
    .B1(_06221_),
    .B2(net7625),
    .X(_06336_));
 sky130_fd_sc_hd__o21a_1 _14074_ (.A1(net1332),
    .A2(_06221_),
    .B1(net7604),
    .X(_06337_));
 sky130_fd_sc_hd__a21o_1 _14075_ (.A1(net1125),
    .A2(_06222_),
    .B1(net7604),
    .X(_06338_));
 sky130_fd_sc_hd__o221a_1 _14076_ (.A1(net7646),
    .A2(_06336_),
    .B1(_06337_),
    .B2(net7633),
    .C1(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__o221a_1 _14077_ (.A1(_06221_),
    .A2(net1125),
    .B1(_06335_),
    .B2(net1597),
    .C1(_06339_),
    .X(_06340_));
 sky130_fd_sc_hd__and2_1 _14078_ (.A(net7666),
    .B(net1123),
    .X(_06341_));
 sky130_fd_sc_hd__nand2_1 _14079_ (.A(net7692),
    .B(net1314),
    .Y(_06342_));
 sky130_fd_sc_hd__nor2_1 _14080_ (.A(net4250),
    .B(_05351_),
    .Y(_06343_));
 sky130_fd_sc_hd__xnor2_1 _14081_ (.A(_06342_),
    .B(_06343_),
    .Y(_06344_));
 sky130_fd_sc_hd__xnor2_1 _14082_ (.A(_06341_),
    .B(_06344_),
    .Y(_06345_));
 sky130_fd_sc_hd__xnor2_1 _14083_ (.A(_06340_),
    .B(_06345_),
    .Y(_06346_));
 sky130_fd_sc_hd__a21bo_1 _14084_ (.A1(_06298_),
    .A2(_06303_),
    .B1_N(_06295_),
    .X(_06347_));
 sky130_fd_sc_hd__o21a_1 _14085_ (.A1(_06298_),
    .A2(_06303_),
    .B1(_06347_),
    .X(_06348_));
 sky130_fd_sc_hd__nand2_2 _14086_ (.A(_06346_),
    .B(_06348_),
    .Y(_06349_));
 sky130_fd_sc_hd__or2_1 _14087_ (.A(_06346_),
    .B(_06348_),
    .X(_06350_));
 sky130_fd_sc_hd__nand2_1 _14088_ (.A(_06349_),
    .B(_06350_),
    .Y(_06351_));
 sky130_fd_sc_hd__xnor2_2 _14089_ (.A(_06332_),
    .B(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__a21bo_1 _14090_ (.A1(_06284_),
    .A2(_06287_),
    .B1_N(_06288_),
    .X(_06353_));
 sky130_fd_sc_hd__o21ai_1 _14091_ (.A1(_06284_),
    .A2(_06287_),
    .B1(_06353_),
    .Y(_06354_));
 sky130_fd_sc_hd__xor2_1 _14092_ (.A(_06352_),
    .B(_06354_),
    .X(_06355_));
 sky130_fd_sc_hd__xnor2_1 _14093_ (.A(_06323_),
    .B(_06355_),
    .Y(_06356_));
 sky130_fd_sc_hd__a21o_1 _14094_ (.A1(_06282_),
    .A2(_06315_),
    .B1(_06317_),
    .X(_06357_));
 sky130_fd_sc_hd__xor2_1 _14095_ (.A(_06356_),
    .B(_06357_),
    .X(_06358_));
 sky130_fd_sc_hd__inv_2 _14096_ (.A(net366),
    .Y(_06359_));
 sky130_fd_sc_hd__a31o_1 _14097_ (.A1(net282),
    .A2(net319),
    .A3(_06359_),
    .B1(_06280_),
    .X(_06360_));
 sky130_fd_sc_hd__a21o_1 _14098_ (.A1(net282),
    .A2(net319),
    .B1(_06359_),
    .X(_06361_));
 sky130_fd_sc_hd__nand2_1 _14099_ (.A(net255),
    .B(net254),
    .Y(_06362_));
 sky130_fd_sc_hd__xnor2_1 _14100_ (.A(_06358_),
    .B(_06362_),
    .Y(_06363_));
 sky130_fd_sc_hd__a22o_1 _14101_ (.A1(net9112),
    .A2(_05780_),
    .B1(net188),
    .B2(net2374),
    .X(_00026_));
 sky130_fd_sc_hd__a22o_1 _14102_ (.A1(_06356_),
    .A2(_06357_),
    .B1(net255),
    .B2(net254),
    .X(_06364_));
 sky130_fd_sc_hd__or2_1 _14103_ (.A(_06356_),
    .B(_06357_),
    .X(_06365_));
 sky130_fd_sc_hd__nand2_1 _14104_ (.A(net217),
    .B(net403),
    .Y(_06366_));
 sky130_fd_sc_hd__o21a_1 _14105_ (.A1(_06323_),
    .A2(_06352_),
    .B1(_06354_),
    .X(_06367_));
 sky130_fd_sc_hd__a21oi_4 _14106_ (.A1(_06323_),
    .A2(_06352_),
    .B1(_06367_),
    .Y(_06368_));
 sky130_fd_sc_hd__nor2_2 _14107_ (.A(_06332_),
    .B(_06351_),
    .Y(_06369_));
 sky130_fd_sc_hd__a21bo_1 _14108_ (.A1(_06325_),
    .A2(_06329_),
    .B1_N(_06330_),
    .X(_06370_));
 sky130_fd_sc_hd__o21ai_1 _14109_ (.A1(_06325_),
    .A2(_06329_),
    .B1(_06370_),
    .Y(_06371_));
 sky130_fd_sc_hd__a21bo_1 _14110_ (.A1(_06341_),
    .A2(_06343_),
    .B1_N(_06342_),
    .X(_06372_));
 sky130_fd_sc_hd__o21ai_1 _14111_ (.A1(_06341_),
    .A2(_06343_),
    .B1(_06372_),
    .Y(_06373_));
 sky130_fd_sc_hd__buf_1 _14112_ (.A(net1566),
    .X(_06374_));
 sky130_fd_sc_hd__nand2_1 _14113_ (.A(net7680),
    .B(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__xnor2_1 _14114_ (.A(net834),
    .B(_06375_),
    .Y(_06376_));
 sky130_fd_sc_hd__xnor2_1 _14115_ (.A(_06349_),
    .B(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__nand2_1 _14116_ (.A(net7647),
    .B(net1123),
    .Y(_06378_));
 sky130_fd_sc_hd__nand2_1 _14117_ (.A(net7666),
    .B(net1314),
    .Y(_06379_));
 sky130_fd_sc_hd__nand2_1 _14118_ (.A(net7627),
    .B(_05348_),
    .Y(_06380_));
 sky130_fd_sc_hd__xnor2_1 _14119_ (.A(_06379_),
    .B(_06380_),
    .Y(_06381_));
 sky130_fd_sc_hd__xor2_1 _14120_ (.A(_06378_),
    .B(_06381_),
    .X(_06382_));
 sky130_fd_sc_hd__and3b_1 _14121_ (.A_N(net1560),
    .B(net1124),
    .C(net7603),
    .X(_06383_));
 sky130_fd_sc_hd__xnor2_1 _14122_ (.A(_06382_),
    .B(_06383_),
    .Y(_06384_));
 sky130_fd_sc_hd__inv_2 _14123_ (.A(_06340_),
    .Y(_06385_));
 sky130_fd_sc_hd__nor2_1 _14124_ (.A(net1597),
    .B(_06221_),
    .Y(_06386_));
 sky130_fd_sc_hd__mux2_1 _14125_ (.A0(_06221_),
    .A1(_06386_),
    .S(net7613),
    .X(_06387_));
 sky130_fd_sc_hd__and3_1 _14126_ (.A(net1332),
    .B(_06221_),
    .C(_06235_),
    .X(_06388_));
 sky130_fd_sc_hd__a21oi_1 _14127_ (.A1(net7625),
    .A2(_06387_),
    .B1(_06388_),
    .Y(_06389_));
 sky130_fd_sc_hd__or4b_1 _14128_ (.A(net1597),
    .B(net1125),
    .C(_06174_),
    .D_N(_06221_),
    .X(_06390_));
 sky130_fd_sc_hd__o221a_1 _14129_ (.A1(_06385_),
    .A2(_06345_),
    .B1(_06389_),
    .B2(_06291_),
    .C1(_06390_),
    .X(_06391_));
 sky130_fd_sc_hd__xor2_1 _14130_ (.A(_06384_),
    .B(_06391_),
    .X(_06392_));
 sky130_fd_sc_hd__xor2_1 _14131_ (.A(_06377_),
    .B(_06392_),
    .X(_06393_));
 sky130_fd_sc_hd__or2_2 _14132_ (.A(_06371_),
    .B(_06393_),
    .X(_06394_));
 sky130_fd_sc_hd__nand2_2 _14133_ (.A(_06371_),
    .B(_06393_),
    .Y(_06395_));
 sky130_fd_sc_hd__nand2_1 _14134_ (.A(_06394_),
    .B(_06395_),
    .Y(_06396_));
 sky130_fd_sc_hd__xor2_1 _14135_ (.A(_06369_),
    .B(_06396_),
    .X(_06397_));
 sky130_fd_sc_hd__xnor2_1 _14136_ (.A(_06368_),
    .B(_06397_),
    .Y(_06398_));
 sky130_fd_sc_hd__xnor2_1 _14137_ (.A(_06366_),
    .B(_06398_),
    .Y(_06399_));
 sky130_fd_sc_hd__a22o_1 _14138_ (.A1(net9198),
    .A2(net1308),
    .B1(net174),
    .B2(net2375),
    .X(_00027_));
 sky130_fd_sc_hd__a21o_1 _14139_ (.A1(_06349_),
    .A2(net834),
    .B1(_06375_),
    .X(_06400_));
 sky130_fd_sc_hd__o21a_1 _14140_ (.A1(_06349_),
    .A2(net834),
    .B1(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__and2b_1 _14141_ (.A_N(_06377_),
    .B(_06392_),
    .X(_06402_));
 sky130_fd_sc_hd__nor2_2 _14142_ (.A(_06384_),
    .B(_06391_),
    .Y(_06403_));
 sky130_fd_sc_hd__nand2_1 _14143_ (.A(net7626),
    .B(net1121),
    .Y(_06404_));
 sky130_fd_sc_hd__clkbuf_1 _14144_ (.A(net1314),
    .X(_06405_));
 sky130_fd_sc_hd__nand2_1 _14145_ (.A(net7647),
    .B(net1120),
    .Y(_06406_));
 sky130_fd_sc_hd__and3_1 _14146_ (.A(net7612),
    .B(_05346_),
    .C(_05709_),
    .X(_06407_));
 sky130_fd_sc_hd__xor2_1 _14147_ (.A(_06406_),
    .B(_06407_),
    .X(_06408_));
 sky130_fd_sc_hd__xnor2_2 _14148_ (.A(_06404_),
    .B(_06408_),
    .Y(_06409_));
 sky130_fd_sc_hd__o211ai_1 _14149_ (.A1(net1560),
    .A2(_06382_),
    .B1(net7603),
    .C1(net1124),
    .Y(_06410_));
 sky130_fd_sc_hd__xor2_2 _14150_ (.A(_06409_),
    .B(net833),
    .X(_06411_));
 sky130_fd_sc_hd__nand2_1 _14151_ (.A(_06378_),
    .B(_06380_),
    .Y(_06412_));
 sky130_fd_sc_hd__nor2_1 _14152_ (.A(_06378_),
    .B(_06380_),
    .Y(_06413_));
 sky130_fd_sc_hd__a31o_1 _14153_ (.A1(net7666),
    .A2(_06405_),
    .A3(_06412_),
    .B1(_06413_),
    .X(_06414_));
 sky130_fd_sc_hd__and3_1 _14154_ (.A(net7662),
    .B(_06374_),
    .C(_06414_),
    .X(_06415_));
 sky130_fd_sc_hd__a21oi_1 _14155_ (.A1(net7662),
    .A2(_06374_),
    .B1(_06414_),
    .Y(_06416_));
 sky130_fd_sc_hd__or2_1 _14156_ (.A(_06415_),
    .B(_06416_),
    .X(_06417_));
 sky130_fd_sc_hd__xnor2_1 _14157_ (.A(_06411_),
    .B(_06417_),
    .Y(_06418_));
 sky130_fd_sc_hd__xnor2_2 _14158_ (.A(_06403_),
    .B(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__xnor2_1 _14159_ (.A(_06402_),
    .B(_06419_),
    .Y(_06420_));
 sky130_fd_sc_hd__xnor2_2 _14160_ (.A(_06401_),
    .B(_06420_),
    .Y(_06421_));
 sky130_fd_sc_hd__and2_1 _14161_ (.A(net403),
    .B(_06368_),
    .X(_06422_));
 sky130_fd_sc_hd__nand2_1 _14162_ (.A(net217),
    .B(_06422_),
    .Y(_06423_));
 sky130_fd_sc_hd__a21o_1 _14163_ (.A1(net217),
    .A2(net403),
    .B1(_06368_),
    .X(_06424_));
 sky130_fd_sc_hd__a21boi_1 _14164_ (.A1(_06368_),
    .A2(_06395_),
    .B1_N(_06394_),
    .Y(_06425_));
 sky130_fd_sc_hd__o2bb2a_1 _14165_ (.A1_N(_06366_),
    .A2_N(_06425_),
    .B1(_06395_),
    .B2(_06368_),
    .X(_06426_));
 sky130_fd_sc_hd__inv_2 _14166_ (.A(_06368_),
    .Y(_06427_));
 sky130_fd_sc_hd__o22a_1 _14167_ (.A1(_06427_),
    .A2(_06394_),
    .B1(_06425_),
    .B2(_06366_),
    .X(_06428_));
 sky130_fd_sc_hd__mux2_1 _14168_ (.A0(_06426_),
    .A1(_06428_),
    .S(_06369_),
    .X(_06429_));
 sky130_fd_sc_hd__o221a_1 _14169_ (.A1(_06394_),
    .A2(_06423_),
    .B1(_06424_),
    .B2(_06395_),
    .C1(_06429_),
    .X(_06430_));
 sky130_fd_sc_hd__xor2_1 _14170_ (.A(_06421_),
    .B(_06430_),
    .X(_06431_));
 sky130_fd_sc_hd__a22o_1 _14171_ (.A1(net9222),
    .A2(net1308),
    .B1(net157),
    .B2(net2375),
    .X(_00028_));
 sky130_fd_sc_hd__a211o_1 _14172_ (.A1(net217),
    .A2(net403),
    .B1(_06368_),
    .C1(_06369_),
    .X(_06432_));
 sky130_fd_sc_hd__a31o_1 _14173_ (.A1(net217),
    .A2(_06369_),
    .A3(_06422_),
    .B1(_06421_),
    .X(_06433_));
 sky130_fd_sc_hd__a21bo_1 _14174_ (.A1(_06432_),
    .A2(_06433_),
    .B1_N(_06394_),
    .X(_06434_));
 sky130_fd_sc_hd__a21o_1 _14175_ (.A1(net217),
    .A2(_06422_),
    .B1(_06369_),
    .X(_06435_));
 sky130_fd_sc_hd__a22o_1 _14176_ (.A1(_06395_),
    .A2(_06421_),
    .B1(_06424_),
    .B2(_06435_),
    .X(_06436_));
 sky130_fd_sc_hd__or2_1 _14177_ (.A(_06395_),
    .B(_06421_),
    .X(_06437_));
 sky130_fd_sc_hd__and3_1 _14178_ (.A(_06434_),
    .B(_06436_),
    .C(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__nor2_2 _14179_ (.A(_06409_),
    .B(net833),
    .Y(_06439_));
 sky130_fd_sc_hd__a32o_1 _14180_ (.A1(net7627),
    .A2(net1123),
    .A3(_06407_),
    .B1(net1120),
    .B2(net7647),
    .X(_06440_));
 sky130_fd_sc_hd__a21o_1 _14181_ (.A1(net7627),
    .A2(net1123),
    .B1(_06407_),
    .X(_06441_));
 sky130_fd_sc_hd__and2_1 _14182_ (.A(_06440_),
    .B(_06441_),
    .X(_06442_));
 sky130_fd_sc_hd__nand2_1 _14183_ (.A(net7626),
    .B(net1120),
    .Y(_06443_));
 sky130_fd_sc_hd__nand2_1 _14184_ (.A(net7602),
    .B(net1121),
    .Y(_06444_));
 sky130_fd_sc_hd__xnor2_2 _14185_ (.A(_06443_),
    .B(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__inv_2 _14186_ (.A(net1304),
    .Y(_06446_));
 sky130_fd_sc_hd__nor2_1 _14187_ (.A(_05972_),
    .B(_06446_),
    .Y(_06447_));
 sky130_fd_sc_hd__xor2_1 _14188_ (.A(_06445_),
    .B(_06447_),
    .X(_06448_));
 sky130_fd_sc_hd__xnor2_1 _14189_ (.A(_06442_),
    .B(_06448_),
    .Y(_06449_));
 sky130_fd_sc_hd__xnor2_2 _14190_ (.A(_06439_),
    .B(_06449_),
    .Y(_06450_));
 sky130_fd_sc_hd__inv_2 _14191_ (.A(_06411_),
    .Y(_06451_));
 sky130_fd_sc_hd__o21ba_1 _14192_ (.A1(_06451_),
    .A2(_06416_),
    .B1_N(_06415_),
    .X(_06452_));
 sky130_fd_sc_hd__inv_2 _14193_ (.A(_06403_),
    .Y(_06453_));
 sky130_fd_sc_hd__and3_1 _14194_ (.A(_06403_),
    .B(_06411_),
    .C(_06415_),
    .X(_06454_));
 sky130_fd_sc_hd__a221o_1 _14195_ (.A1(_06451_),
    .A2(_06416_),
    .B1(_06452_),
    .B2(_06453_),
    .C1(_06454_),
    .X(_06455_));
 sky130_fd_sc_hd__xnor2_1 _14196_ (.A(_06450_),
    .B(_06455_),
    .Y(_06456_));
 sky130_fd_sc_hd__a21bo_1 _14197_ (.A1(_06401_),
    .A2(_06419_),
    .B1_N(_06402_),
    .X(_06457_));
 sky130_fd_sc_hd__o21a_1 _14198_ (.A1(_06401_),
    .A2(_06419_),
    .B1(_06457_),
    .X(_06458_));
 sky130_fd_sc_hd__nor2_1 _14199_ (.A(_06456_),
    .B(_06458_),
    .Y(_06459_));
 sky130_fd_sc_hd__nand2_1 _14200_ (.A(_06456_),
    .B(_06458_),
    .Y(_06460_));
 sky130_fd_sc_hd__or2b_1 _14201_ (.A(_06459_),
    .B_N(_06460_),
    .X(_06461_));
 sky130_fd_sc_hd__xnor2_1 _14202_ (.A(_06438_),
    .B(_06461_),
    .Y(_06462_));
 sky130_fd_sc_hd__a22o_1 _14203_ (.A1(net9126),
    .A2(_05779_),
    .B1(net160),
    .B2(net2373),
    .X(_00029_));
 sky130_fd_sc_hd__o21ai_1 _14204_ (.A1(_06438_),
    .A2(_06459_),
    .B1(_06460_),
    .Y(_06463_));
 sky130_fd_sc_hd__or2b_1 _14205_ (.A(_06415_),
    .B_N(_06450_),
    .X(_06464_));
 sky130_fd_sc_hd__a2bb2o_1 _14206_ (.A1_N(_06416_),
    .A2_N(_06450_),
    .B1(_06464_),
    .B2(_06411_),
    .X(_06465_));
 sky130_fd_sc_hd__a2bb2o_1 _14207_ (.A1_N(_06450_),
    .A2_N(_06452_),
    .B1(_06465_),
    .B2(_06403_),
    .X(_06466_));
 sky130_fd_sc_hd__nor2_1 _14208_ (.A(_06439_),
    .B(_06442_),
    .Y(_06467_));
 sky130_fd_sc_hd__nand2_1 _14209_ (.A(_06439_),
    .B(_06442_),
    .Y(_06468_));
 sky130_fd_sc_hd__a21oi_1 _14210_ (.A1(_06445_),
    .A2(_06468_),
    .B1(_06467_),
    .Y(_06469_));
 sky130_fd_sc_hd__o2bb2a_2 _14211_ (.A1_N(_06445_),
    .A2_N(_06467_),
    .B1(_06469_),
    .B2(_06447_),
    .X(_06470_));
 sky130_fd_sc_hd__nand2_1 _14212_ (.A(net7602),
    .B(net1119),
    .Y(_06471_));
 sky130_fd_sc_hd__o21a_1 _14213_ (.A1(net1121),
    .A2(net1304),
    .B1(net7629),
    .X(_06472_));
 sky130_fd_sc_hd__o211a_1 _14214_ (.A1(net1121),
    .A2(_06471_),
    .B1(net1304),
    .C1(net7629),
    .X(_06473_));
 sky130_fd_sc_hd__o21ba_1 _14215_ (.A1(_06471_),
    .A2(_06472_),
    .B1_N(_06473_),
    .X(_06474_));
 sky130_fd_sc_hd__xnor2_1 _14216_ (.A(_06470_),
    .B(_06474_),
    .Y(_06475_));
 sky130_fd_sc_hd__and2_1 _14217_ (.A(_06466_),
    .B(_06475_),
    .X(_06476_));
 sky130_fd_sc_hd__or2_1 _14218_ (.A(_06466_),
    .B(_06475_),
    .X(_06477_));
 sky130_fd_sc_hd__and2b_1 _14219_ (.A_N(_06476_),
    .B(_06477_),
    .X(_06478_));
 sky130_fd_sc_hd__xnor2_1 _14220_ (.A(_06463_),
    .B(_06478_),
    .Y(_06479_));
 sky130_fd_sc_hd__a22o_1 _14221_ (.A1(net9157),
    .A2(_05779_),
    .B1(net156),
    .B2(net2373),
    .X(_00030_));
 sky130_fd_sc_hd__a41o_1 _14222_ (.A1(_06434_),
    .A2(_06436_),
    .A3(_06437_),
    .A4(_06460_),
    .B1(_06459_),
    .X(_06480_));
 sky130_fd_sc_hd__a21oi_1 _14223_ (.A1(_06477_),
    .A2(_06480_),
    .B1(_06476_),
    .Y(_06481_));
 sky130_fd_sc_hd__and3_1 _14224_ (.A(net7629),
    .B(net1304),
    .C(_06470_),
    .X(_06482_));
 sky130_fd_sc_hd__a21o_1 _14225_ (.A1(net1119),
    .A2(_06470_),
    .B1(net7626),
    .X(_06483_));
 sky130_fd_sc_hd__o21ai_1 _14226_ (.A1(net1119),
    .A2(_06470_),
    .B1(_06483_),
    .Y(_06484_));
 sky130_fd_sc_hd__o21ba_1 _14227_ (.A1(_06446_),
    .A2(_06470_),
    .B1_N(_06404_),
    .X(_06485_));
 sky130_fd_sc_hd__a21o_1 _14228_ (.A1(_06446_),
    .A2(_06470_),
    .B1(_06485_),
    .X(_06486_));
 sky130_fd_sc_hd__a22o_1 _14229_ (.A1(net1304),
    .A2(_06484_),
    .B1(_06486_),
    .B2(net1119),
    .X(_06487_));
 sky130_fd_sc_hd__mux2_1 _14230_ (.A0(_06482_),
    .A1(_06487_),
    .S(net7602),
    .X(_06488_));
 sky130_fd_sc_hd__xnor2_1 _14231_ (.A(_06481_),
    .B(_06488_),
    .Y(_06489_));
 sky130_fd_sc_hd__a22o_1 _14232_ (.A1(net9091),
    .A2(_05779_),
    .B1(net154),
    .B2(net2373),
    .X(_00031_));
 sky130_fd_sc_hd__a21bo_1 _14233_ (.A1(_06466_),
    .A2(_06475_),
    .B1_N(_06463_),
    .X(_06490_));
 sky130_fd_sc_hd__a21o_1 _14234_ (.A1(net7629),
    .A2(net1304),
    .B1(net1119),
    .X(_06491_));
 sky130_fd_sc_hd__a22o_1 _14235_ (.A1(net1119),
    .A2(_06472_),
    .B1(_06491_),
    .B2(_06470_),
    .X(_06492_));
 sky130_fd_sc_hd__and2_1 _14236_ (.A(net1304),
    .B(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__nor2_1 _14237_ (.A(_06446_),
    .B(_06481_),
    .Y(_06494_));
 sky130_fd_sc_hd__a311o_1 _14238_ (.A1(_06477_),
    .A2(_06490_),
    .A3(_06492_),
    .B1(_06493_),
    .C1(_06494_),
    .X(_06495_));
 sky130_fd_sc_hd__a32o_1 _14239_ (.A1(net7606),
    .A2(net2373),
    .A3(net153),
    .B1(_05779_),
    .B2(net9194),
    .X(_00032_));
 sky130_fd_sc_hd__o21a_1 _14240_ (.A1(net6456),
    .A2(net6649),
    .B1(net6446),
    .X(_06496_));
 sky130_fd_sc_hd__or3b_1 _14241_ (.A(net6456),
    .B(net6446),
    .C_N(net8319),
    .X(_06497_));
 sky130_fd_sc_hd__a21o_1 _14242_ (.A1(net152),
    .A2(_06497_),
    .B1(net6451),
    .X(_06498_));
 sky130_fd_sc_hd__o21a_1 _14243_ (.A1(net152),
    .A2(_06496_),
    .B1(_06498_),
    .X(_00033_));
 sky130_fd_sc_hd__inv_2 _14244_ (.A(net8062),
    .Y(_06499_));
 sky130_fd_sc_hd__nand2_1 _14245_ (.A(_06499_),
    .B(net7535),
    .Y(_06500_));
 sky130_fd_sc_hd__buf_1 _14246_ (.A(_06500_),
    .X(_06501_));
 sky130_fd_sc_hd__buf_1 _14247_ (.A(_06501_),
    .X(_06502_));
 sky130_fd_sc_hd__or2_1 _14248_ (.A(net6508),
    .B(net6496),
    .X(_06503_));
 sky130_fd_sc_hd__or2_1 _14249_ (.A(net6477),
    .B(net6467),
    .X(_06504_));
 sky130_fd_sc_hd__nor2_1 _14250_ (.A(net4238),
    .B(_06504_),
    .Y(_06505_));
 sky130_fd_sc_hd__nand2_1 _14251_ (.A(net6458),
    .B(_06505_),
    .Y(_06506_));
 sky130_fd_sc_hd__nand2_1 _14252_ (.A(net8047),
    .B(net2932),
    .Y(_06507_));
 sky130_fd_sc_hd__buf_1 _14253_ (.A(net2284),
    .X(_06508_));
 sky130_fd_sc_hd__buf_1 _14254_ (.A(net1916),
    .X(_06509_));
 sky130_fd_sc_hd__nand2_1 _14255_ (.A(net2285),
    .B(net1554),
    .Y(_00034_));
 sky130_fd_sc_hd__nor2_1 _14256_ (.A(net6451),
    .B(_06497_),
    .Y(_06510_));
 sky130_fd_sc_hd__buf_1 _14257_ (.A(net3658),
    .X(_06511_));
 sky130_fd_sc_hd__inv_2 _14258_ (.A(net6451),
    .Y(_06512_));
 sky130_fd_sc_hd__nand2_1 _14259_ (.A(net6455),
    .B(net6445),
    .Y(_06513_));
 sky130_fd_sc_hd__o21ba_1 _14260_ (.A1(net4236),
    .A2(_06513_),
    .B1_N(net3666),
    .X(_06514_));
 sky130_fd_sc_hd__buf_1 _14261_ (.A(net2923),
    .X(_06515_));
 sky130_fd_sc_hd__a22o_1 _14262_ (.A1(net49),
    .A2(net2931),
    .B1(net2278),
    .B2(net9010),
    .X(_00035_));
 sky130_fd_sc_hd__a22o_1 _14263_ (.A1(net56),
    .A2(net2931),
    .B1(net2278),
    .B2(net8986),
    .X(_00036_));
 sky130_fd_sc_hd__a22o_1 _14264_ (.A1(net57),
    .A2(net2931),
    .B1(net2278),
    .B2(net9023),
    .X(_00037_));
 sky130_fd_sc_hd__a22o_1 _14265_ (.A1(net58),
    .A2(_06511_),
    .B1(_06515_),
    .B2(net8985),
    .X(_00038_));
 sky130_fd_sc_hd__a22o_1 _14266_ (.A1(net59),
    .A2(net2931),
    .B1(net2278),
    .B2(net9004),
    .X(_00039_));
 sky130_fd_sc_hd__a22o_1 _14267_ (.A1(net60),
    .A2(_06511_),
    .B1(_06515_),
    .B2(net9014),
    .X(_00040_));
 sky130_fd_sc_hd__a22o_1 _14268_ (.A1(net61),
    .A2(net2931),
    .B1(net2278),
    .B2(net9053),
    .X(_00041_));
 sky130_fd_sc_hd__a22o_1 _14269_ (.A1(net62),
    .A2(net2931),
    .B1(net2278),
    .B2(net9060),
    .X(_00042_));
 sky130_fd_sc_hd__a22o_1 _14270_ (.A1(net63),
    .A2(net2931),
    .B1(net2278),
    .B2(net9103),
    .X(_00043_));
 sky130_fd_sc_hd__a22o_1 _14271_ (.A1(net64),
    .A2(_06511_),
    .B1(_06515_),
    .B2(net8999),
    .X(_00044_));
 sky130_fd_sc_hd__clkbuf_1 _14272_ (.A(net3657),
    .X(_06516_));
 sky130_fd_sc_hd__clkbuf_2 _14273_ (.A(net2922),
    .X(_06517_));
 sky130_fd_sc_hd__a22o_1 _14274_ (.A1(net50),
    .A2(net2914),
    .B1(_06517_),
    .B2(net9078),
    .X(_00045_));
 sky130_fd_sc_hd__a22o_1 _14275_ (.A1(net51),
    .A2(net2902),
    .B1(net2265),
    .B2(net9011),
    .X(_00046_));
 sky130_fd_sc_hd__a22o_1 _14276_ (.A1(net52),
    .A2(net2903),
    .B1(net2266),
    .B2(net7973),
    .X(_00047_));
 sky130_fd_sc_hd__a22o_1 _14277_ (.A1(net53),
    .A2(net2914),
    .B1(_06517_),
    .B2(net9042),
    .X(_00048_));
 sky130_fd_sc_hd__a22o_1 _14278_ (.A1(net54),
    .A2(net2914),
    .B1(_06517_),
    .B2(net8990),
    .X(_00049_));
 sky130_fd_sc_hd__a22o_1 _14279_ (.A1(net55),
    .A2(net2914),
    .B1(_06517_),
    .B2(net7954),
    .X(_00050_));
 sky130_fd_sc_hd__a22o_1 _14280_ (.A1(net65),
    .A2(net2902),
    .B1(net2265),
    .B2(net7934),
    .X(_00051_));
 sky130_fd_sc_hd__a22o_1 _14281_ (.A1(net72),
    .A2(net2902),
    .B1(net2265),
    .B2(net7914),
    .X(_00052_));
 sky130_fd_sc_hd__a22o_1 _14282_ (.A1(net73),
    .A2(net2902),
    .B1(net2265),
    .B2(net7880),
    .X(_00053_));
 sky130_fd_sc_hd__a22o_1 _14283_ (.A1(net8118),
    .A2(net2902),
    .B1(net2265),
    .B2(net7855),
    .X(_00054_));
 sky130_fd_sc_hd__clkbuf_2 _14284_ (.A(net3649),
    .X(_06518_));
 sky130_fd_sc_hd__clkbuf_2 _14285_ (.A(net2915),
    .X(_06519_));
 sky130_fd_sc_hd__a22o_1 _14286_ (.A1(net75),
    .A2(_06518_),
    .B1(_06519_),
    .B2(net7820),
    .X(_00055_));
 sky130_fd_sc_hd__a22o_1 _14287_ (.A1(net76),
    .A2(_06518_),
    .B1(_06519_),
    .B2(net7819),
    .X(_00056_));
 sky130_fd_sc_hd__a22o_1 _14288_ (.A1(net77),
    .A2(_06518_),
    .B1(_06519_),
    .B2(net7791),
    .X(_00057_));
 sky130_fd_sc_hd__a22o_1 _14289_ (.A1(net78),
    .A2(net2901),
    .B1(net2264),
    .B2(net7771),
    .X(_00058_));
 sky130_fd_sc_hd__a22o_1 _14290_ (.A1(net79),
    .A2(net2901),
    .B1(net2264),
    .B2(net7734),
    .X(_00059_));
 sky130_fd_sc_hd__a22o_1 _14291_ (.A1(net80),
    .A2(_06518_),
    .B1(_06519_),
    .B2(net7724),
    .X(_00060_));
 sky130_fd_sc_hd__a22o_1 _14292_ (.A1(net66),
    .A2(_06518_),
    .B1(_06519_),
    .B2(net7711),
    .X(_00061_));
 sky130_fd_sc_hd__a22o_1 _14293_ (.A1(net67),
    .A2(net2901),
    .B1(net2264),
    .B2(net7684),
    .X(_00062_));
 sky130_fd_sc_hd__a22o_1 _14294_ (.A1(net68),
    .A2(net2901),
    .B1(net2264),
    .B2(net7670),
    .X(_00063_));
 sky130_fd_sc_hd__a22o_1 _14295_ (.A1(net69),
    .A2(net2901),
    .B1(net2264),
    .B2(net7649),
    .X(_00064_));
 sky130_fd_sc_hd__a22o_1 _14296_ (.A1(net70),
    .A2(net3649),
    .B1(net2915),
    .B2(net7634),
    .X(_00065_));
 sky130_fd_sc_hd__a22o_1 _14297_ (.A1(net71),
    .A2(net3649),
    .B1(net2915),
    .B2(net7614),
    .X(_00066_));
 sky130_fd_sc_hd__xor2_1 _14298_ (.A(net6455),
    .B(net6445),
    .X(_06520_));
 sky130_fd_sc_hd__and3_1 _14299_ (.A(net4236),
    .B(net1991),
    .C(_06520_),
    .X(_06521_));
 sky130_fd_sc_hd__buf_1 _14300_ (.A(net1549),
    .X(_06522_));
 sky130_fd_sc_hd__nand2_1 _14301_ (.A(net6451),
    .B(net6456),
    .Y(_06523_));
 sky130_fd_sc_hd__nor2_1 _14302_ (.A(net6446),
    .B(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__buf_1 _14303_ (.A(_06524_),
    .X(_06525_));
 sky130_fd_sc_hd__nor3_1 _14304_ (.A(net6448),
    .B(net6454),
    .C(net6444),
    .Y(_06526_));
 sky130_fd_sc_hd__clkbuf_1 _14305_ (.A(_06526_),
    .X(_06527_));
 sky130_fd_sc_hd__and2_1 _14306_ (.A(net8312),
    .B(net3645),
    .X(_06528_));
 sky130_fd_sc_hd__a221o_1 _14307_ (.A1(\matmul0.alpha_pass[0] ),
    .A2(net1302),
    .B1(net2898),
    .B2(net5367),
    .C1(_06528_),
    .X(_06529_));
 sky130_fd_sc_hd__inv_2 _14308_ (.A(net6453),
    .Y(_06530_));
 sky130_fd_sc_hd__nor2_1 _14309_ (.A(net6450),
    .B(_06513_),
    .Y(_06531_));
 sky130_fd_sc_hd__nand2_1 _14310_ (.A(net6750),
    .B(net6604),
    .Y(_06532_));
 sky130_fd_sc_hd__buf_1 _14311_ (.A(_06532_),
    .X(_06533_));
 sky130_fd_sc_hd__or3_1 _14312_ (.A(net6451),
    .B(net6456),
    .C(net8319),
    .X(_06534_));
 sky130_fd_sc_hd__o21a_1 _14313_ (.A1(net5370),
    .A2(_06523_),
    .B1(_06534_),
    .X(_06535_));
 sky130_fd_sc_hd__nor2_1 _14314_ (.A(net6443),
    .B(_06535_),
    .Y(_06536_));
 sky130_fd_sc_hd__a31o_1 _14315_ (.A1(\matmul0.state[1] ),
    .A2(net6597),
    .A3(cordic_done),
    .B1(net6432),
    .X(_06537_));
 sky130_fd_sc_hd__o21a_1 _14316_ (.A1(clarke_done),
    .A2(net2386),
    .B1(_06537_),
    .X(_06538_));
 sky130_fd_sc_hd__or4_1 _14317_ (.A(net6448),
    .B(_06530_),
    .C(net6443),
    .D(_06538_),
    .X(_06539_));
 sky130_fd_sc_hd__inv_2 _14318_ (.A(_06539_),
    .Y(_06540_));
 sky130_fd_sc_hd__a311o_2 _14319_ (.A1(net4235),
    .A2(net6443),
    .A3(net3638),
    .B1(_06536_),
    .C1(_06540_),
    .X(_06541_));
 sky130_fd_sc_hd__a211o_1 _14320_ (.A1(net6447),
    .A2(_06530_),
    .B1(_06531_),
    .C1(_06541_),
    .X(_06542_));
 sky130_fd_sc_hd__buf_1 _14321_ (.A(_06542_),
    .X(_06543_));
 sky130_fd_sc_hd__mux2_1 _14322_ (.A0(_06529_),
    .A1(\matmul0.a_in[0] ),
    .S(net904),
    .X(_06544_));
 sky130_fd_sc_hd__clkbuf_1 _14323_ (.A(_06544_),
    .X(_00067_));
 sky130_fd_sc_hd__and2_1 _14324_ (.A(net8271),
    .B(net3642),
    .X(_06545_));
 sky130_fd_sc_hd__a221o_1 _14325_ (.A1(net7356),
    .A2(net1299),
    .B1(net2896),
    .B2(\pid_d.out[1] ),
    .C1(_06545_),
    .X(_06546_));
 sky130_fd_sc_hd__mux2_1 _14326_ (.A0(_06546_),
    .A1(\matmul0.a_in[1] ),
    .S(net902),
    .X(_06547_));
 sky130_fd_sc_hd__clkbuf_1 _14327_ (.A(_06547_),
    .X(_00068_));
 sky130_fd_sc_hd__and2_1 _14328_ (.A(net8262),
    .B(net3642),
    .X(_06548_));
 sky130_fd_sc_hd__a221o_1 _14329_ (.A1(net7346),
    .A2(net1299),
    .B1(net2896),
    .B2(\pid_d.out[2] ),
    .C1(_06548_),
    .X(_06549_));
 sky130_fd_sc_hd__mux2_1 _14330_ (.A0(_06549_),
    .A1(\matmul0.a_in[2] ),
    .S(net902),
    .X(_06550_));
 sky130_fd_sc_hd__clkbuf_1 _14331_ (.A(_06550_),
    .X(_00069_));
 sky130_fd_sc_hd__and2_1 _14332_ (.A(net8253),
    .B(net3642),
    .X(_06551_));
 sky130_fd_sc_hd__a221o_1 _14333_ (.A1(net7332),
    .A2(net1299),
    .B1(net2896),
    .B2(\pid_d.out[3] ),
    .C1(_06551_),
    .X(_06552_));
 sky130_fd_sc_hd__mux2_1 _14334_ (.A0(_06552_),
    .A1(\matmul0.a_in[3] ),
    .S(net902),
    .X(_06553_));
 sky130_fd_sc_hd__clkbuf_1 _14335_ (.A(_06553_),
    .X(_00070_));
 sky130_fd_sc_hd__and2_1 _14336_ (.A(net8243),
    .B(net3642),
    .X(_06554_));
 sky130_fd_sc_hd__a221o_1 _14337_ (.A1(net7320),
    .A2(net1299),
    .B1(net2896),
    .B2(\pid_d.out[4] ),
    .C1(_06554_),
    .X(_06555_));
 sky130_fd_sc_hd__mux2_1 _14338_ (.A0(_06555_),
    .A1(\matmul0.a_in[4] ),
    .S(net902),
    .X(_06556_));
 sky130_fd_sc_hd__clkbuf_1 _14339_ (.A(_06556_),
    .X(_00071_));
 sky130_fd_sc_hd__and2_1 _14340_ (.A(net8233),
    .B(net3643),
    .X(_06557_));
 sky130_fd_sc_hd__a221o_1 _14341_ (.A1(net7309),
    .A2(net1299),
    .B1(net2896),
    .B2(\pid_d.out[5] ),
    .C1(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__mux2_1 _14342_ (.A0(_06558_),
    .A1(\matmul0.a_in[5] ),
    .S(net902),
    .X(_06559_));
 sky130_fd_sc_hd__clkbuf_1 _14343_ (.A(_06559_),
    .X(_00072_));
 sky130_fd_sc_hd__and2_1 _14344_ (.A(net8225),
    .B(net3645),
    .X(_06560_));
 sky130_fd_sc_hd__a221o_1 _14345_ (.A1(net7299),
    .A2(net1301),
    .B1(net2898),
    .B2(net5361),
    .C1(_06560_),
    .X(_06561_));
 sky130_fd_sc_hd__mux2_1 _14346_ (.A0(_06561_),
    .A1(\matmul0.a_in[6] ),
    .S(net904),
    .X(_06562_));
 sky130_fd_sc_hd__clkbuf_1 _14347_ (.A(_06562_),
    .X(_00073_));
 sky130_fd_sc_hd__and2_1 _14348_ (.A(net8217),
    .B(net3646),
    .X(_06563_));
 sky130_fd_sc_hd__a221o_1 _14349_ (.A1(net7291),
    .A2(net1301),
    .B1(net2899),
    .B2(net5358),
    .C1(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__mux2_1 _14350_ (.A0(_06564_),
    .A1(\matmul0.a_in[7] ),
    .S(net903),
    .X(_06565_));
 sky130_fd_sc_hd__clkbuf_1 _14351_ (.A(_06565_),
    .X(_00074_));
 sky130_fd_sc_hd__and2_1 _14352_ (.A(net8210),
    .B(net3646),
    .X(_06566_));
 sky130_fd_sc_hd__a221o_1 _14353_ (.A1(net7280),
    .A2(_06522_),
    .B1(net2900),
    .B2(net5355),
    .C1(_06566_),
    .X(_06567_));
 sky130_fd_sc_hd__mux2_1 _14354_ (.A0(_06567_),
    .A1(\matmul0.a_in[8] ),
    .S(net905),
    .X(_06568_));
 sky130_fd_sc_hd__clkbuf_1 _14355_ (.A(_06568_),
    .X(_00075_));
 sky130_fd_sc_hd__buf_1 _14356_ (.A(net3647),
    .X(_06569_));
 sky130_fd_sc_hd__and2_1 _14357_ (.A(net8204),
    .B(_06527_),
    .X(_06570_));
 sky130_fd_sc_hd__a221o_1 _14358_ (.A1(net7271),
    .A2(net1303),
    .B1(net2895),
    .B2(net5351),
    .C1(_06570_),
    .X(_06571_));
 sky130_fd_sc_hd__buf_1 _14359_ (.A(net994),
    .X(_06572_));
 sky130_fd_sc_hd__mux2_1 _14360_ (.A0(_06571_),
    .A1(\matmul0.a_in[9] ),
    .S(net901),
    .X(_06573_));
 sky130_fd_sc_hd__clkbuf_1 _14361_ (.A(_06573_),
    .X(_00076_));
 sky130_fd_sc_hd__buf_1 _14362_ (.A(net1548),
    .X(_06574_));
 sky130_fd_sc_hd__buf_1 _14363_ (.A(net4233),
    .X(_06575_));
 sky130_fd_sc_hd__and2_1 _14364_ (.A(net8305),
    .B(net3636),
    .X(_06576_));
 sky130_fd_sc_hd__a221o_1 _14365_ (.A1(net7259),
    .A2(_06574_),
    .B1(_06569_),
    .B2(net5346),
    .C1(_06576_),
    .X(_06577_));
 sky130_fd_sc_hd__mux2_1 _14366_ (.A0(_06577_),
    .A1(\matmul0.a_in[10] ),
    .S(_06572_),
    .X(_06578_));
 sky130_fd_sc_hd__clkbuf_1 _14367_ (.A(_06578_),
    .X(_00077_));
 sky130_fd_sc_hd__and2_1 _14368_ (.A(net8300),
    .B(net3637),
    .X(_06579_));
 sky130_fd_sc_hd__a221o_1 _14369_ (.A1(net7247),
    .A2(net1296),
    .B1(net2893),
    .B2(net5341),
    .C1(_06579_),
    .X(_06580_));
 sky130_fd_sc_hd__mux2_1 _14370_ (.A0(_06580_),
    .A1(\matmul0.a_in[11] ),
    .S(net899),
    .X(_06581_));
 sky130_fd_sc_hd__clkbuf_1 _14371_ (.A(_06581_),
    .X(_00078_));
 sky130_fd_sc_hd__and2_1 _14372_ (.A(net8295),
    .B(_06575_),
    .X(_06582_));
 sky130_fd_sc_hd__a221o_1 _14373_ (.A1(net7225),
    .A2(net1297),
    .B1(net2894),
    .B2(net5333),
    .C1(_06582_),
    .X(_06583_));
 sky130_fd_sc_hd__mux2_1 _14374_ (.A0(_06583_),
    .A1(\matmul0.a_in[12] ),
    .S(net900),
    .X(_06584_));
 sky130_fd_sc_hd__clkbuf_1 _14375_ (.A(_06584_),
    .X(_00079_));
 sky130_fd_sc_hd__and2_1 _14376_ (.A(net8290),
    .B(net3637),
    .X(_06585_));
 sky130_fd_sc_hd__a221o_1 _14377_ (.A1(net7217),
    .A2(net1296),
    .B1(net2893),
    .B2(net5328),
    .C1(_06585_),
    .X(_06586_));
 sky130_fd_sc_hd__mux2_1 _14378_ (.A0(_06586_),
    .A1(\matmul0.a_in[13] ),
    .S(net899),
    .X(_06587_));
 sky130_fd_sc_hd__clkbuf_1 _14379_ (.A(_06587_),
    .X(_00080_));
 sky130_fd_sc_hd__and2_1 _14380_ (.A(net8285),
    .B(net3637),
    .X(_06588_));
 sky130_fd_sc_hd__a221o_1 _14381_ (.A1(net7210),
    .A2(net1296),
    .B1(net2893),
    .B2(net5320),
    .C1(_06588_),
    .X(_06589_));
 sky130_fd_sc_hd__mux2_1 _14382_ (.A0(_06589_),
    .A1(net7584),
    .S(net899),
    .X(_06590_));
 sky130_fd_sc_hd__clkbuf_1 _14383_ (.A(_06590_),
    .X(_00081_));
 sky130_fd_sc_hd__and2_1 _14384_ (.A(net8280),
    .B(net3637),
    .X(_06591_));
 sky130_fd_sc_hd__a221o_1 _14385_ (.A1(net7198),
    .A2(net1296),
    .B1(net2893),
    .B2(net5315),
    .C1(_06591_),
    .X(_06592_));
 sky130_fd_sc_hd__mux2_1 _14386_ (.A0(_06592_),
    .A1(net7580),
    .S(net899),
    .X(_06593_));
 sky130_fd_sc_hd__clkbuf_1 _14387_ (.A(_06593_),
    .X(_00082_));
 sky130_fd_sc_hd__and2_1 _14388_ (.A(net8198),
    .B(net3636),
    .X(_06594_));
 sky130_fd_sc_hd__a221o_1 _14389_ (.A1(net5312),
    .A2(net1297),
    .B1(net2895),
    .B2(net4471),
    .C1(_06594_),
    .X(_06595_));
 sky130_fd_sc_hd__mux2_1 _14390_ (.A0(_06595_),
    .A1(\matmul0.b_in[0] ),
    .S(net900),
    .X(_06596_));
 sky130_fd_sc_hd__clkbuf_1 _14391_ (.A(_06596_),
    .X(_00083_));
 sky130_fd_sc_hd__and2_1 _14392_ (.A(net8163),
    .B(net3635),
    .X(_06597_));
 sky130_fd_sc_hd__a221o_1 _14393_ (.A1(net5306),
    .A2(net1297),
    .B1(net2894),
    .B2(net4467),
    .C1(_06597_),
    .X(_06598_));
 sky130_fd_sc_hd__mux2_1 _14394_ (.A0(_06598_),
    .A1(\matmul0.b_in[1] ),
    .S(net900),
    .X(_06599_));
 sky130_fd_sc_hd__clkbuf_1 _14395_ (.A(_06599_),
    .X(_00084_));
 sky130_fd_sc_hd__and2_1 _14396_ (.A(net8157),
    .B(net3635),
    .X(_06600_));
 sky130_fd_sc_hd__a221o_1 _14397_ (.A1(net5297),
    .A2(net1298),
    .B1(net2895),
    .B2(net4463),
    .C1(_06600_),
    .X(_06601_));
 sky130_fd_sc_hd__mux2_1 _14398_ (.A0(_06601_),
    .A1(\matmul0.b_in[2] ),
    .S(net901),
    .X(_06602_));
 sky130_fd_sc_hd__clkbuf_1 _14399_ (.A(_06602_),
    .X(_00085_));
 sky130_fd_sc_hd__buf_1 _14400_ (.A(net3647),
    .X(_06603_));
 sky130_fd_sc_hd__and2_1 _14401_ (.A(net8151),
    .B(net3635),
    .X(_06604_));
 sky130_fd_sc_hd__a221o_1 _14402_ (.A1(net5289),
    .A2(net1298),
    .B1(net2892),
    .B2(net4458),
    .C1(_06604_),
    .X(_06605_));
 sky130_fd_sc_hd__buf_1 _14403_ (.A(net994),
    .X(_06606_));
 sky130_fd_sc_hd__mux2_1 _14404_ (.A0(_06605_),
    .A1(\matmul0.b_in[3] ),
    .S(net898),
    .X(_06607_));
 sky130_fd_sc_hd__clkbuf_1 _14405_ (.A(_06607_),
    .X(_00086_));
 sky130_fd_sc_hd__buf_1 _14406_ (.A(net1548),
    .X(_06608_));
 sky130_fd_sc_hd__clkbuf_1 _14407_ (.A(net4233),
    .X(_06609_));
 sky130_fd_sc_hd__and2_1 _14408_ (.A(net8146),
    .B(net3633),
    .X(_06610_));
 sky130_fd_sc_hd__a221o_1 _14409_ (.A1(net5282),
    .A2(net1295),
    .B1(net2891),
    .B2(net4452),
    .C1(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__mux2_1 _14410_ (.A0(_06611_),
    .A1(\matmul0.b_in[4] ),
    .S(net897),
    .X(_06612_));
 sky130_fd_sc_hd__clkbuf_1 _14411_ (.A(_06612_),
    .X(_00087_));
 sky130_fd_sc_hd__and2_1 _14412_ (.A(net8141),
    .B(net3634),
    .X(_06613_));
 sky130_fd_sc_hd__a221o_1 _14413_ (.A1(net5272),
    .A2(_06608_),
    .B1(_06603_),
    .B2(net4448),
    .C1(_06613_),
    .X(_06614_));
 sky130_fd_sc_hd__mux2_1 _14414_ (.A0(_06614_),
    .A1(\matmul0.b_in[5] ),
    .S(_06606_),
    .X(_06615_));
 sky130_fd_sc_hd__clkbuf_1 _14415_ (.A(_06615_),
    .X(_00088_));
 sky130_fd_sc_hd__and2_1 _14416_ (.A(net8136),
    .B(net3632),
    .X(_06616_));
 sky130_fd_sc_hd__a221o_1 _14417_ (.A1(\matmul0.beta_pass[6] ),
    .A2(net1294),
    .B1(net2890),
    .B2(net4443),
    .C1(_06616_),
    .X(_06617_));
 sky130_fd_sc_hd__mux2_1 _14418_ (.A0(_06617_),
    .A1(\matmul0.b_in[6] ),
    .S(net896),
    .X(_06618_));
 sky130_fd_sc_hd__clkbuf_1 _14419_ (.A(_06618_),
    .X(_00089_));
 sky130_fd_sc_hd__and2_1 _14420_ (.A(net8132),
    .B(net3631),
    .X(_06619_));
 sky130_fd_sc_hd__a221o_1 _14421_ (.A1(\matmul0.beta_pass[7] ),
    .A2(net1293),
    .B1(net2889),
    .B2(net4436),
    .C1(_06619_),
    .X(_06620_));
 sky130_fd_sc_hd__mux2_1 _14422_ (.A0(_06620_),
    .A1(\matmul0.b_in[7] ),
    .S(net895),
    .X(_06621_));
 sky130_fd_sc_hd__clkbuf_1 _14423_ (.A(_06621_),
    .X(_00090_));
 sky130_fd_sc_hd__and2_1 _14424_ (.A(net8127),
    .B(net3633),
    .X(_06622_));
 sky130_fd_sc_hd__a221o_1 _14425_ (.A1(net5243),
    .A2(net1295),
    .B1(net2891),
    .B2(net4431),
    .C1(_06622_),
    .X(_06623_));
 sky130_fd_sc_hd__mux2_1 _14426_ (.A0(_06623_),
    .A1(\matmul0.b_in[8] ),
    .S(net897),
    .X(_06624_));
 sky130_fd_sc_hd__clkbuf_1 _14427_ (.A(_06624_),
    .X(_00091_));
 sky130_fd_sc_hd__and2_1 _14428_ (.A(net8123),
    .B(net3631),
    .X(_06625_));
 sky130_fd_sc_hd__a221o_1 _14429_ (.A1(\matmul0.beta_pass[9] ),
    .A2(net1293),
    .B1(net2889),
    .B2(net4425),
    .C1(_06625_),
    .X(_06626_));
 sky130_fd_sc_hd__mux2_1 _14430_ (.A0(_06626_),
    .A1(\matmul0.b_in[9] ),
    .S(net895),
    .X(_06627_));
 sky130_fd_sc_hd__clkbuf_1 _14431_ (.A(_06627_),
    .X(_00092_));
 sky130_fd_sc_hd__and2_1 _14432_ (.A(net8194),
    .B(net3632),
    .X(_06628_));
 sky130_fd_sc_hd__a221o_1 _14433_ (.A1(net5219),
    .A2(net1294),
    .B1(net2890),
    .B2(net4419),
    .C1(_06628_),
    .X(_06629_));
 sky130_fd_sc_hd__mux2_1 _14434_ (.A0(_06629_),
    .A1(\matmul0.b_in[10] ),
    .S(net896),
    .X(_06630_));
 sky130_fd_sc_hd__clkbuf_1 _14435_ (.A(_06630_),
    .X(_00093_));
 sky130_fd_sc_hd__and2_1 _14436_ (.A(net8190),
    .B(net3632),
    .X(_06631_));
 sky130_fd_sc_hd__a221o_1 _14437_ (.A1(\matmul0.beta_pass[11] ),
    .A2(net1294),
    .B1(net2890),
    .B2(net4413),
    .C1(_06631_),
    .X(_06632_));
 sky130_fd_sc_hd__mux2_1 _14438_ (.A0(_06632_),
    .A1(\matmul0.b_in[11] ),
    .S(net896),
    .X(_06633_));
 sky130_fd_sc_hd__clkbuf_1 _14439_ (.A(_06633_),
    .X(_00094_));
 sky130_fd_sc_hd__and2_1 _14440_ (.A(net8186),
    .B(net3631),
    .X(_06634_));
 sky130_fd_sc_hd__a221o_1 _14441_ (.A1(net5210),
    .A2(net1293),
    .B1(net2889),
    .B2(net4407),
    .C1(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__mux2_1 _14442_ (.A0(_06635_),
    .A1(\matmul0.b_in[12] ),
    .S(net895),
    .X(_06636_));
 sky130_fd_sc_hd__clkbuf_1 _14443_ (.A(_06636_),
    .X(_00095_));
 sky130_fd_sc_hd__and2_1 _14444_ (.A(net8180),
    .B(net3634),
    .X(_06637_));
 sky130_fd_sc_hd__a221o_1 _14445_ (.A1(net5202),
    .A2(_06608_),
    .B1(net3647),
    .B2(net4402),
    .C1(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__mux2_1 _14446_ (.A0(_06638_),
    .A1(\matmul0.b_in[13] ),
    .S(net994),
    .X(_06639_));
 sky130_fd_sc_hd__clkbuf_1 _14447_ (.A(_06639_),
    .X(_00096_));
 sky130_fd_sc_hd__and2_1 _14448_ (.A(net8174),
    .B(net4233),
    .X(_06640_));
 sky130_fd_sc_hd__a221o_1 _14449_ (.A1(net5197),
    .A2(net1548),
    .B1(net3647),
    .B2(net4397),
    .C1(_06640_),
    .X(_06641_));
 sky130_fd_sc_hd__mux2_1 _14450_ (.A0(_06641_),
    .A1(\matmul0.b_in[14] ),
    .S(net994),
    .X(_06642_));
 sky130_fd_sc_hd__clkbuf_1 _14451_ (.A(_06642_),
    .X(_00097_));
 sky130_fd_sc_hd__and2_1 _14452_ (.A(net8168),
    .B(net4234),
    .X(_06643_));
 sky130_fd_sc_hd__a221o_1 _14453_ (.A1(net5192),
    .A2(net1550),
    .B1(net3648),
    .B2(net4394),
    .C1(_06643_),
    .X(_06644_));
 sky130_fd_sc_hd__mux2_1 _14454_ (.A0(_06644_),
    .A1(\matmul0.b_in[15] ),
    .S(net995),
    .X(_06645_));
 sky130_fd_sc_hd__clkbuf_1 _14455_ (.A(_06645_),
    .X(_00098_));
 sky130_fd_sc_hd__inv_2 _14456_ (.A(_06541_),
    .Y(_06646_));
 sky130_fd_sc_hd__o211a_1 _14457_ (.A1(net6454),
    .A2(\matmul0.op_in[0] ),
    .B1(_06513_),
    .C1(net6447),
    .X(_06647_));
 sky130_fd_sc_hd__o221a_1 _14458_ (.A1(_06530_),
    .A2(\matmul0.op_in[0] ),
    .B1(_06541_),
    .B2(net6443),
    .C1(net4235),
    .X(_06648_));
 sky130_fd_sc_hd__o22a_1 _14459_ (.A1(net9192),
    .A2(_06646_),
    .B1(_06647_),
    .B2(_06648_),
    .X(_00099_));
 sky130_fd_sc_hd__nor2_1 _14460_ (.A(net6443),
    .B(_06541_),
    .Y(_06649_));
 sky130_fd_sc_hd__a22o_1 _14461_ (.A1(net9086),
    .A2(_06543_),
    .B1(_06649_),
    .B2(net6453),
    .X(_00100_));
 sky130_fd_sc_hd__or2_1 _14462_ (.A(_06513_),
    .B(_06541_),
    .X(_06650_));
 sky130_fd_sc_hd__buf_1 _14463_ (.A(_06650_),
    .X(_06651_));
 sky130_fd_sc_hd__buf_1 _14464_ (.A(net892),
    .X(_06652_));
 sky130_fd_sc_hd__buf_1 _14465_ (.A(_06531_),
    .X(_06653_));
 sky130_fd_sc_hd__and2_1 _14466_ (.A(net1990),
    .B(net2887),
    .X(_06654_));
 sky130_fd_sc_hd__buf_1 _14467_ (.A(_06654_),
    .X(_06655_));
 sky130_fd_sc_hd__xor2_1 _14468_ (.A(net7364),
    .B(net5311),
    .X(_06656_));
 sky130_fd_sc_hd__a22o_1 _14469_ (.A1(net9072),
    .A2(net831),
    .B1(net1292),
    .B2(_06656_),
    .X(_00101_));
 sky130_fd_sc_hd__or2_1 _14470_ (.A(net7361),
    .B(net5305),
    .X(_06657_));
 sky130_fd_sc_hd__nand2_1 _14471_ (.A(net7361),
    .B(net5305),
    .Y(_06658_));
 sky130_fd_sc_hd__nor2_1 _14472_ (.A(net7365),
    .B(net5311),
    .Y(_06659_));
 sky130_fd_sc_hd__a21oi_1 _14473_ (.A1(_06657_),
    .A2(_06658_),
    .B1(_06659_),
    .Y(_06660_));
 sky130_fd_sc_hd__and3_1 _14474_ (.A(_06659_),
    .B(_06657_),
    .C(_06658_),
    .X(_06661_));
 sky130_fd_sc_hd__or2_1 _14475_ (.A(_06660_),
    .B(_06661_),
    .X(_06662_));
 sky130_fd_sc_hd__a22o_1 _14476_ (.A1(net9070),
    .A2(net831),
    .B1(net1292),
    .B2(_06662_),
    .X(_00102_));
 sky130_fd_sc_hd__xnor2_1 _14477_ (.A(net7340),
    .B(net5296),
    .Y(_06663_));
 sky130_fd_sc_hd__mux2_1 _14478_ (.A0(_06658_),
    .A1(_06657_),
    .S(_06659_),
    .X(_06664_));
 sky130_fd_sc_hd__xnor2_1 _14479_ (.A(_06663_),
    .B(_06664_),
    .Y(_06665_));
 sky130_fd_sc_hd__a22o_1 _14480_ (.A1(net9095),
    .A2(net831),
    .B1(net1292),
    .B2(_06665_),
    .X(_00103_));
 sky130_fd_sc_hd__a21oi_1 _14481_ (.A1(net7361),
    .A2(net5305),
    .B1(_06663_),
    .Y(_06666_));
 sky130_fd_sc_hd__o2bb2a_1 _14482_ (.A1_N(_06657_),
    .A2_N(_06663_),
    .B1(_06666_),
    .B2(_06659_),
    .X(_06667_));
 sky130_fd_sc_hd__nor2_1 _14483_ (.A(net7340),
    .B(net5294),
    .Y(_06668_));
 sky130_fd_sc_hd__xor2_2 _14484_ (.A(net7336),
    .B(net5287),
    .X(_06669_));
 sky130_fd_sc_hd__xnor2_1 _14485_ (.A(_06668_),
    .B(_06669_),
    .Y(_06670_));
 sky130_fd_sc_hd__xnor2_1 _14486_ (.A(_06667_),
    .B(_06670_),
    .Y(_06671_));
 sky130_fd_sc_hd__a22o_1 _14487_ (.A1(net9051),
    .A2(net832),
    .B1(net1292),
    .B2(_06671_),
    .X(_00104_));
 sky130_fd_sc_hd__a21o_1 _14488_ (.A1(_06667_),
    .A2(_06669_),
    .B1(_06668_),
    .X(_06672_));
 sky130_fd_sc_hd__o21ai_2 _14489_ (.A1(_06667_),
    .A2(_06669_),
    .B1(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__nor2_1 _14490_ (.A(net7336),
    .B(net5286),
    .Y(_06674_));
 sky130_fd_sc_hd__xnor2_2 _14491_ (.A(net7324),
    .B(net5279),
    .Y(_06675_));
 sky130_fd_sc_hd__xnor2_1 _14492_ (.A(_06674_),
    .B(_06675_),
    .Y(_06676_));
 sky130_fd_sc_hd__xnor2_1 _14493_ (.A(_06673_),
    .B(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__a22o_1 _14494_ (.A1(net9047),
    .A2(net831),
    .B1(net1292),
    .B2(_06677_),
    .X(_00105_));
 sky130_fd_sc_hd__o21ba_1 _14495_ (.A1(_06673_),
    .A2(_06675_),
    .B1_N(_06674_),
    .X(_06678_));
 sky130_fd_sc_hd__a21o_1 _14496_ (.A1(_06673_),
    .A2(_06675_),
    .B1(_06678_),
    .X(_06679_));
 sky130_fd_sc_hd__nor2_1 _14497_ (.A(net7324),
    .B(net5278),
    .Y(_06680_));
 sky130_fd_sc_hd__xnor2_2 _14498_ (.A(net7313),
    .B(net5270),
    .Y(_06681_));
 sky130_fd_sc_hd__xnor2_1 _14499_ (.A(_06680_),
    .B(_06681_),
    .Y(_06682_));
 sky130_fd_sc_hd__xnor2_1 _14500_ (.A(_06679_),
    .B(_06682_),
    .Y(_06683_));
 sky130_fd_sc_hd__a22o_1 _14501_ (.A1(net9058),
    .A2(net832),
    .B1(net1292),
    .B2(_06683_),
    .X(_00106_));
 sky130_fd_sc_hd__o21ba_1 _14502_ (.A1(_06679_),
    .A2(_06681_),
    .B1_N(_06680_),
    .X(_06684_));
 sky130_fd_sc_hd__a21o_1 _14503_ (.A1(_06679_),
    .A2(_06681_),
    .B1(_06684_),
    .X(_06685_));
 sky130_fd_sc_hd__or2_1 _14504_ (.A(net7313),
    .B(net5269),
    .X(_06686_));
 sky130_fd_sc_hd__xnor2_1 _14505_ (.A(net7302),
    .B(net5262),
    .Y(_06687_));
 sky130_fd_sc_hd__xnor2_1 _14506_ (.A(_06686_),
    .B(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__nand2_1 _14507_ (.A(_06685_),
    .B(_06688_),
    .Y(_06689_));
 sky130_fd_sc_hd__or2_1 _14508_ (.A(_06685_),
    .B(_06688_),
    .X(_06690_));
 sky130_fd_sc_hd__a32o_1 _14509_ (.A1(_06655_),
    .A2(_06689_),
    .A3(_06690_),
    .B1(net893),
    .B2(net9005),
    .X(_00107_));
 sky130_fd_sc_hd__xor2_1 _14510_ (.A(net7282),
    .B(net5254),
    .X(_06691_));
 sky130_fd_sc_hd__nand2_1 _14511_ (.A(net3032),
    .B(_06691_),
    .Y(_06692_));
 sky130_fd_sc_hd__o21a_1 _14512_ (.A1(net7313),
    .A2(net5269),
    .B1(_06685_),
    .X(_06693_));
 sky130_fd_sc_hd__or3_1 _14513_ (.A(net7313),
    .B(net5267),
    .C(_06685_),
    .X(_06694_));
 sky130_fd_sc_hd__o21a_1 _14514_ (.A1(net5262),
    .A2(_06693_),
    .B1(_06694_),
    .X(_06695_));
 sky130_fd_sc_hd__nand2_1 _14515_ (.A(net5262),
    .B(_06693_),
    .Y(_06696_));
 sky130_fd_sc_hd__o311a_1 _14516_ (.A1(net7302),
    .A2(net5262),
    .A3(_06694_),
    .B1(_06696_),
    .C1(net1990),
    .X(_06697_));
 sky130_fd_sc_hd__a21bo_1 _14517_ (.A1(net7302),
    .A2(_06695_),
    .B1_N(_06697_),
    .X(_06698_));
 sky130_fd_sc_hd__xor2_1 _14518_ (.A(_06692_),
    .B(_06698_),
    .X(_06699_));
 sky130_fd_sc_hd__a22o_1 _14519_ (.A1(net9068),
    .A2(net832),
    .B1(_06699_),
    .B2(net2886),
    .X(_00108_));
 sky130_fd_sc_hd__a21o_1 _14520_ (.A1(_06692_),
    .A2(_06694_),
    .B1(net5262),
    .X(_06700_));
 sky130_fd_sc_hd__o21a_1 _14521_ (.A1(_06692_),
    .A2(_06693_),
    .B1(_06700_),
    .X(_06701_));
 sky130_fd_sc_hd__o221a_1 _14522_ (.A1(_06692_),
    .A2(_06695_),
    .B1(_06701_),
    .B2(net7302),
    .C1(net2389),
    .X(_06702_));
 sky130_fd_sc_hd__or2_1 _14523_ (.A(net7282),
    .B(net5253),
    .X(_06703_));
 sky130_fd_sc_hd__xnor2_1 _14524_ (.A(net7278),
    .B(net5246),
    .Y(_06704_));
 sky130_fd_sc_hd__xnor2_1 _14525_ (.A(_06703_),
    .B(_06704_),
    .Y(_06705_));
 sky130_fd_sc_hd__nand2_1 _14526_ (.A(net1625),
    .B(_06705_),
    .Y(_06706_));
 sky130_fd_sc_hd__xnor2_1 _14527_ (.A(net726),
    .B(_06706_),
    .Y(_06707_));
 sky130_fd_sc_hd__a22o_1 _14528_ (.A1(net9030),
    .A2(_06652_),
    .B1(net676),
    .B2(net2886),
    .X(_00109_));
 sky130_fd_sc_hd__inv_2 _14529_ (.A(net7279),
    .Y(_06708_));
 sky130_fd_sc_hd__and2_1 _14530_ (.A(net726),
    .B(_06703_),
    .X(_06709_));
 sky130_fd_sc_hd__clkbuf_2 _14531_ (.A(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__xor2_4 _14532_ (.A(net7264),
    .B(net5239),
    .X(_06711_));
 sky130_fd_sc_hd__a21o_1 _14533_ (.A1(net2388),
    .A2(_06703_),
    .B1(net726),
    .X(_06712_));
 sky130_fd_sc_hd__a21o_1 _14534_ (.A1(_06711_),
    .A2(_06712_),
    .B1(net5247),
    .X(_06713_));
 sky130_fd_sc_hd__o21ai_1 _14535_ (.A1(_06710_),
    .A2(_06711_),
    .B1(_06713_),
    .Y(_06714_));
 sky130_fd_sc_hd__o21a_1 _14536_ (.A1(net5247),
    .A2(_06710_),
    .B1(net7278),
    .X(_06715_));
 sky130_fd_sc_hd__a21o_1 _14537_ (.A1(net5247),
    .A2(_06710_),
    .B1(_06715_),
    .X(_06716_));
 sky130_fd_sc_hd__nor2_1 _14538_ (.A(net726),
    .B(_06703_),
    .Y(_06717_));
 sky130_fd_sc_hd__nor3_1 _14539_ (.A(net5247),
    .B(_06710_),
    .C(_06711_),
    .Y(_06718_));
 sky130_fd_sc_hd__clkbuf_1 _14540_ (.A(net3639),
    .X(_06719_));
 sky130_fd_sc_hd__a311o_1 _14541_ (.A1(net7278),
    .A2(net5247),
    .A3(_06717_),
    .B1(_06718_),
    .C1(net2885),
    .X(_06720_));
 sky130_fd_sc_hd__a221o_1 _14542_ (.A1(net4225),
    .A2(_06714_),
    .B1(_06716_),
    .B2(_06711_),
    .C1(_06720_),
    .X(_06721_));
 sky130_fd_sc_hd__nand2_1 _14543_ (.A(net7278),
    .B(_06711_),
    .Y(_06722_));
 sky130_fd_sc_hd__or3_1 _14544_ (.A(net7278),
    .B(net5250),
    .C(_06711_),
    .X(_06723_));
 sky130_fd_sc_hd__a31o_1 _14545_ (.A1(net1624),
    .A2(_06722_),
    .A3(_06723_),
    .B1(_06712_),
    .X(_06724_));
 sky130_fd_sc_hd__a32o_1 _14546_ (.A1(_06653_),
    .A2(_06721_),
    .A3(_06724_),
    .B1(_06651_),
    .B2(net8964),
    .X(_00110_));
 sky130_fd_sc_hd__inv_2 _14547_ (.A(_06711_),
    .Y(_06725_));
 sky130_fd_sc_hd__nor2_1 _14548_ (.A(_06711_),
    .B(_06717_),
    .Y(_06726_));
 sky130_fd_sc_hd__o22a_1 _14549_ (.A1(_06710_),
    .A2(_06725_),
    .B1(_06726_),
    .B2(net5250),
    .X(_06727_));
 sky130_fd_sc_hd__o21ai_1 _14550_ (.A1(net5250),
    .A2(_06710_),
    .B1(_06712_),
    .Y(_06728_));
 sky130_fd_sc_hd__a21oi_1 _14551_ (.A1(_06711_),
    .A2(_06728_),
    .B1(net3639),
    .Y(_06729_));
 sky130_fd_sc_hd__o21a_2 _14552_ (.A1(net7278),
    .A2(_06727_),
    .B1(_06729_),
    .X(_06730_));
 sky130_fd_sc_hd__or2_2 _14553_ (.A(net7264),
    .B(net5238),
    .X(_06731_));
 sky130_fd_sc_hd__xnor2_1 _14554_ (.A(net7257),
    .B(net5223),
    .Y(_06732_));
 sky130_fd_sc_hd__nor2_1 _14555_ (.A(_06731_),
    .B(_06732_),
    .Y(_06733_));
 sky130_fd_sc_hd__and2_1 _14556_ (.A(_06731_),
    .B(_06732_),
    .X(_06734_));
 sky130_fd_sc_hd__o21ai_1 _14557_ (.A1(_06733_),
    .A2(_06734_),
    .B1(net1625),
    .Y(_06735_));
 sky130_fd_sc_hd__xnor2_1 _14558_ (.A(_06730_),
    .B(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__a22o_1 _14559_ (.A1(net9056),
    .A2(net832),
    .B1(net448),
    .B2(net2886),
    .X(_00111_));
 sky130_fd_sc_hd__or3_1 _14560_ (.A(net7257),
    .B(net5222),
    .C(_06731_),
    .X(_06737_));
 sky130_fd_sc_hd__and2_1 _14561_ (.A(net5223),
    .B(_06731_),
    .X(_06738_));
 sky130_fd_sc_hd__nor2_1 _14562_ (.A(net7257),
    .B(net5223),
    .Y(_06739_));
 sky130_fd_sc_hd__a21o_1 _14563_ (.A1(net7257),
    .A2(_06738_),
    .B1(_06739_),
    .X(_06740_));
 sky130_fd_sc_hd__xor2_2 _14564_ (.A(net7244),
    .B(net5213),
    .X(_06741_));
 sky130_fd_sc_hd__mux2_1 _14565_ (.A0(_06737_),
    .A1(_06740_),
    .S(_06741_),
    .X(_06742_));
 sky130_fd_sc_hd__a21o_1 _14566_ (.A1(net1625),
    .A2(_06742_),
    .B1(_06730_),
    .X(_06743_));
 sky130_fd_sc_hd__o21a_1 _14567_ (.A1(net7260),
    .A2(net3640),
    .B1(_06730_),
    .X(_06744_));
 sky130_fd_sc_hd__o32a_1 _14568_ (.A1(net5223),
    .A2(net3640),
    .A3(_06731_),
    .B1(_06730_),
    .B2(net7260),
    .X(_06745_));
 sky130_fd_sc_hd__o21ai_1 _14569_ (.A1(_06738_),
    .A2(_06744_),
    .B1(_06745_),
    .Y(_06746_));
 sky130_fd_sc_hd__o21a_1 _14570_ (.A1(_06730_),
    .A2(_06731_),
    .B1(_06739_),
    .X(_06747_));
 sky130_fd_sc_hd__nor2_1 _14571_ (.A(_06733_),
    .B(_06747_),
    .Y(_06748_));
 sky130_fd_sc_hd__mux2_1 _14572_ (.A0(_06746_),
    .A1(_06748_),
    .S(_06741_),
    .X(_06749_));
 sky130_fd_sc_hd__or2_1 _14573_ (.A(net2884),
    .B(_06749_),
    .X(_06750_));
 sky130_fd_sc_hd__a32o_1 _14574_ (.A1(net2888),
    .A2(_06743_),
    .A3(_06750_),
    .B1(net894),
    .B2(net8967),
    .X(_00112_));
 sky130_fd_sc_hd__a21oi_1 _14575_ (.A1(net2389),
    .A2(_06737_),
    .B1(_06730_),
    .Y(_06751_));
 sky130_fd_sc_hd__a21oi_2 _14576_ (.A1(_06741_),
    .A2(_06746_),
    .B1(_06751_),
    .Y(_06752_));
 sky130_fd_sc_hd__nor2_1 _14577_ (.A(net7244),
    .B(net5213),
    .Y(_06753_));
 sky130_fd_sc_hd__xnor2_2 _14578_ (.A(net7234),
    .B(net5207),
    .Y(_06754_));
 sky130_fd_sc_hd__xor2_1 _14579_ (.A(_06753_),
    .B(_06754_),
    .X(_06755_));
 sky130_fd_sc_hd__nand2_1 _14580_ (.A(_04860_),
    .B(_06755_),
    .Y(_06756_));
 sky130_fd_sc_hd__xnor2_1 _14581_ (.A(_06752_),
    .B(_06756_),
    .Y(_06757_));
 sky130_fd_sc_hd__a22o_1 _14582_ (.A1(net9115),
    .A2(_06652_),
    .B1(net318),
    .B2(net2886),
    .X(_00113_));
 sky130_fd_sc_hd__a21oi_1 _14583_ (.A1(net2390),
    .A2(_06754_),
    .B1(_06752_),
    .Y(_06758_));
 sky130_fd_sc_hd__o21ai_1 _14584_ (.A1(net3640),
    .A2(_06754_),
    .B1(_06752_),
    .Y(_06759_));
 sky130_fd_sc_hd__o21a_1 _14585_ (.A1(_06753_),
    .A2(_06758_),
    .B1(_06759_),
    .X(_06760_));
 sky130_fd_sc_hd__nor2_1 _14586_ (.A(net7233),
    .B(net5207),
    .Y(_06761_));
 sky130_fd_sc_hd__xnor2_2 _14587_ (.A(net7214),
    .B(net5198),
    .Y(_06762_));
 sky130_fd_sc_hd__xnor2_1 _14588_ (.A(_06761_),
    .B(_06762_),
    .Y(_06763_));
 sky130_fd_sc_hd__or3_1 _14589_ (.A(net2882),
    .B(net281),
    .C(_06763_),
    .X(_06764_));
 sky130_fd_sc_hd__o21ai_1 _14590_ (.A1(net2882),
    .A2(_06763_),
    .B1(net281),
    .Y(_06765_));
 sky130_fd_sc_hd__a32o_1 _14591_ (.A1(net2887),
    .A2(_06764_),
    .A3(_06765_),
    .B1(net892),
    .B2(net8995),
    .X(_00114_));
 sky130_fd_sc_hd__a21boi_1 _14592_ (.A1(net1989),
    .A2(_06762_),
    .B1_N(net281),
    .Y(_06766_));
 sky130_fd_sc_hd__nor2_1 _14593_ (.A(net3641),
    .B(_06762_),
    .Y(_06767_));
 sky130_fd_sc_hd__o22a_1 _14594_ (.A1(_06761_),
    .A2(_06766_),
    .B1(_06767_),
    .B2(net281),
    .X(_06768_));
 sky130_fd_sc_hd__xnor2_1 _14595_ (.A(net7209),
    .B(net5195),
    .Y(_06769_));
 sky130_fd_sc_hd__or3_1 _14596_ (.A(net7214),
    .B(net5200),
    .C(_06769_),
    .X(_06770_));
 sky130_fd_sc_hd__o21ai_1 _14597_ (.A1(net7214),
    .A2(net5200),
    .B1(_06769_),
    .Y(_06771_));
 sky130_fd_sc_hd__a21oi_1 _14598_ (.A1(_06770_),
    .A2(_06771_),
    .B1(net2882),
    .Y(_06772_));
 sky130_fd_sc_hd__xnor2_1 _14599_ (.A(_06768_),
    .B(_06772_),
    .Y(_06773_));
 sky130_fd_sc_hd__a22o_1 _14600_ (.A1(net9084),
    .A2(net892),
    .B1(_06773_),
    .B2(net2887),
    .X(_00115_));
 sky130_fd_sc_hd__xnor2_1 _14601_ (.A(net7199),
    .B(net5190),
    .Y(_06774_));
 sky130_fd_sc_hd__nor2_1 _14602_ (.A(net7209),
    .B(net5194),
    .Y(_06775_));
 sky130_fd_sc_hd__xnor2_1 _14603_ (.A(_06774_),
    .B(_06775_),
    .Y(_06776_));
 sky130_fd_sc_hd__nor2_1 _14604_ (.A(net3641),
    .B(_06776_),
    .Y(_06777_));
 sky130_fd_sc_hd__mux2_1 _14605_ (.A0(_06771_),
    .A1(_06770_),
    .S(_06777_),
    .X(_06778_));
 sky130_fd_sc_hd__inv_2 _14606_ (.A(_06778_),
    .Y(_06779_));
 sky130_fd_sc_hd__mux2_1 _14607_ (.A0(_06770_),
    .A1(_06771_),
    .S(_06777_),
    .X(_06780_));
 sky130_fd_sc_hd__and2_1 _14608_ (.A(_06768_),
    .B(_06777_),
    .X(_06781_));
 sky130_fd_sc_hd__nor2_1 _14609_ (.A(_06768_),
    .B(_06777_),
    .Y(_06782_));
 sky130_fd_sc_hd__o221a_1 _14610_ (.A1(net2882),
    .A2(_06780_),
    .B1(_06781_),
    .B2(_06782_),
    .C1(net2887),
    .X(_06783_));
 sky130_fd_sc_hd__a221o_1 _14611_ (.A1(net9097),
    .A2(net892),
    .B1(_06655_),
    .B2(_06779_),
    .C1(_06783_),
    .X(_00116_));
 sky130_fd_sc_hd__nand2_1 _14612_ (.A(_06512_),
    .B(net6443),
    .Y(_06784_));
 sky130_fd_sc_hd__or2_1 _14613_ (.A(_06512_),
    .B(net6443),
    .X(_06785_));
 sky130_fd_sc_hd__and3_1 _14614_ (.A(net6453),
    .B(_06784_),
    .C(_06785_),
    .X(_06786_));
 sky130_fd_sc_hd__a21o_1 _14615_ (.A1(net6432),
    .A2(_06786_),
    .B1(cordic_done),
    .X(_06787_));
 sky130_fd_sc_hd__nand2_1 _14616_ (.A(_06539_),
    .B(_06786_),
    .Y(_06788_));
 sky130_fd_sc_hd__and2_1 _14617_ (.A(_06787_),
    .B(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__clkbuf_1 _14618_ (.A(_06789_),
    .X(_00117_));
 sky130_fd_sc_hd__a21o_1 _14619_ (.A1(net1622),
    .A2(_06786_),
    .B1(clarke_done),
    .X(_06790_));
 sky130_fd_sc_hd__and2_1 _14620_ (.A(_06788_),
    .B(_06790_),
    .X(_06791_));
 sky130_fd_sc_hd__clkbuf_1 _14621_ (.A(_06791_),
    .X(_00118_));
 sky130_fd_sc_hd__a21bo_1 _14622_ (.A1(net6446),
    .A2(\cordic0.in_valid ),
    .B1_N(_06497_),
    .X(_06792_));
 sky130_fd_sc_hd__nand2_1 _14623_ (.A(net6456),
    .B(_06785_),
    .Y(_06793_));
 sky130_fd_sc_hd__a22o_1 _14624_ (.A1(_06512_),
    .A2(_06792_),
    .B1(_06793_),
    .B2(net9102),
    .X(_00119_));
 sky130_fd_sc_hd__nor2_1 _14625_ (.A(net6448),
    .B(_06541_),
    .Y(_06794_));
 sky130_fd_sc_hd__a31o_1 _14626_ (.A1(net6448),
    .A2(net6443),
    .A3(\matmul0.start ),
    .B1(_06794_),
    .X(_06795_));
 sky130_fd_sc_hd__a22o_1 _14627_ (.A1(\matmul0.start ),
    .A2(_06536_),
    .B1(_06649_),
    .B2(net6453),
    .X(_06796_));
 sky130_fd_sc_hd__a21o_1 _14628_ (.A1(_06530_),
    .A2(_06795_),
    .B1(_06796_),
    .X(_00120_));
 sky130_fd_sc_hd__nor2_1 _14629_ (.A(net2881),
    .B(_06785_),
    .Y(_06797_));
 sky130_fd_sc_hd__o21a_1 _14630_ (.A1(net8992),
    .A2(_06797_),
    .B1(_06523_),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _14631_ (.A0(net7551),
    .A1(net7461),
    .S(_04877_),
    .X(_06798_));
 sky130_fd_sc_hd__clkbuf_1 _14632_ (.A(_06798_),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _14633_ (.A0(net7550),
    .A1(\matmul0.op[1] ),
    .S(net3704),
    .X(_06799_));
 sky130_fd_sc_hd__clkbuf_1 _14634_ (.A(_06799_),
    .X(_00123_));
 sky130_fd_sc_hd__clkbuf_1 _14635_ (.A(net4282),
    .X(_06800_));
 sky130_fd_sc_hd__clkbuf_2 _14636_ (.A(net3629),
    .X(_06801_));
 sky130_fd_sc_hd__buf_1 _14637_ (.A(net3697),
    .X(_06802_));
 sky130_fd_sc_hd__and3_1 _14638_ (.A(net7437),
    .B(\matmul0.cos[0] ),
    .C(net2878),
    .X(_06803_));
 sky130_fd_sc_hd__a21o_1 _14639_ (.A1(net8960),
    .A2(net2879),
    .B1(_06803_),
    .X(_00124_));
 sky130_fd_sc_hd__and3_1 _14640_ (.A(net7437),
    .B(net7182),
    .C(net2878),
    .X(_06804_));
 sky130_fd_sc_hd__a21o_1 _14641_ (.A1(net8979),
    .A2(net2879),
    .B1(_06804_),
    .X(_00125_));
 sky130_fd_sc_hd__clkbuf_1 _14642_ (.A(net3697),
    .X(_06805_));
 sky130_fd_sc_hd__and3_1 _14643_ (.A(net7439),
    .B(net7181),
    .C(net2875),
    .X(_06806_));
 sky130_fd_sc_hd__a21o_1 _14644_ (.A1(net8959),
    .A2(net2880),
    .B1(_06806_),
    .X(_00126_));
 sky130_fd_sc_hd__and3_1 _14645_ (.A(net7437),
    .B(\matmul0.cos[4] ),
    .C(_06805_),
    .X(_06807_));
 sky130_fd_sc_hd__a21o_1 _14646_ (.A1(net8969),
    .A2(net2879),
    .B1(_06807_),
    .X(_00127_));
 sky130_fd_sc_hd__and3_1 _14647_ (.A(net7440),
    .B(net7178),
    .C(net2874),
    .X(_06808_));
 sky130_fd_sc_hd__a21o_1 _14648_ (.A1(net8961),
    .A2(_06801_),
    .B1(_06808_),
    .X(_00128_));
 sky130_fd_sc_hd__and3_1 _14649_ (.A(net7437),
    .B(\matmul0.cos[6] ),
    .C(net2875),
    .X(_06809_));
 sky130_fd_sc_hd__a21o_1 _14650_ (.A1(net8989),
    .A2(net2880),
    .B1(_06809_),
    .X(_00129_));
 sky130_fd_sc_hd__and3_1 _14651_ (.A(net7440),
    .B(net7175),
    .C(net2874),
    .X(_06810_));
 sky130_fd_sc_hd__a21o_1 _14652_ (.A1(net8958),
    .A2(_06801_),
    .B1(_06810_),
    .X(_00130_));
 sky130_fd_sc_hd__and3_1 _14653_ (.A(net7440),
    .B(net7172),
    .C(net2874),
    .X(_06811_));
 sky130_fd_sc_hd__a21o_1 _14654_ (.A1(net8970),
    .A2(_06801_),
    .B1(_06811_),
    .X(_00131_));
 sky130_fd_sc_hd__and3_1 _14655_ (.A(net7439),
    .B(net7170),
    .C(net2874),
    .X(_06812_));
 sky130_fd_sc_hd__a21o_1 _14656_ (.A1(net8965),
    .A2(_06801_),
    .B1(_06812_),
    .X(_00132_));
 sky130_fd_sc_hd__and3_1 _14657_ (.A(net7439),
    .B(net7169),
    .C(net2875),
    .X(_06813_));
 sky130_fd_sc_hd__a21o_1 _14658_ (.A1(net8956),
    .A2(net2880),
    .B1(_06813_),
    .X(_00133_));
 sky130_fd_sc_hd__buf_1 _14659_ (.A(net3628),
    .X(_06814_));
 sky130_fd_sc_hd__and3_1 _14660_ (.A(net7446),
    .B(net7168),
    .C(net2873),
    .X(_06815_));
 sky130_fd_sc_hd__a21o_1 _14661_ (.A1(net9021),
    .A2(net2872),
    .B1(_06815_),
    .X(_00134_));
 sky130_fd_sc_hd__and3_1 _14662_ (.A(net7442),
    .B(net7167),
    .C(net2873),
    .X(_06816_));
 sky130_fd_sc_hd__a21o_1 _14663_ (.A1(net8982),
    .A2(_06814_),
    .B1(_06816_),
    .X(_00135_));
 sky130_fd_sc_hd__inv_2 _14664_ (.A(net7441),
    .Y(_06817_));
 sky130_fd_sc_hd__buf_1 _14665_ (.A(_06817_),
    .X(_06818_));
 sky130_fd_sc_hd__o21a_1 _14666_ (.A1(net3625),
    .A2(net7166),
    .B1(net2876),
    .X(_06819_));
 sky130_fd_sc_hd__a21o_1 _14667_ (.A1(net9024),
    .A2(net2872),
    .B1(_06819_),
    .X(_00136_));
 sky130_fd_sc_hd__buf_1 _14668_ (.A(net3630),
    .X(_06820_));
 sky130_fd_sc_hd__nand2_1 _14669_ (.A(net7455),
    .B(net7163),
    .Y(_06821_));
 sky130_fd_sc_hd__xnor2_1 _14670_ (.A(net7160),
    .B(_06821_),
    .Y(_06822_));
 sky130_fd_sc_hd__buf_1 _14671_ (.A(net4281),
    .X(_06823_));
 sky130_fd_sc_hd__nor2_1 _14672_ (.A(_06817_),
    .B(net3620),
    .Y(_06824_));
 sky130_fd_sc_hd__a22o_1 _14673_ (.A1(net9081),
    .A2(net2869),
    .B1(_06822_),
    .B2(net2865),
    .X(_00137_));
 sky130_fd_sc_hd__buf_1 _14674_ (.A(net2865),
    .X(_06825_));
 sky130_fd_sc_hd__inv_2 _14675_ (.A(net7454),
    .Y(_06826_));
 sky130_fd_sc_hd__nor2_1 _14676_ (.A(net7160),
    .B(net7164),
    .Y(_06827_));
 sky130_fd_sc_hd__or2_1 _14677_ (.A(net4223),
    .B(_06827_),
    .X(_06828_));
 sky130_fd_sc_hd__xnor2_1 _14678_ (.A(net7158),
    .B(_06828_),
    .Y(_06829_));
 sky130_fd_sc_hd__a22o_1 _14679_ (.A1(net7433),
    .A2(net2869),
    .B1(net2263),
    .B2(net2864),
    .X(_00138_));
 sky130_fd_sc_hd__o31a_1 _14680_ (.A1(net7160),
    .A2(net7164),
    .A3(net7158),
    .B1(net7453),
    .X(_06830_));
 sky130_fd_sc_hd__xor2_1 _14681_ (.A(net7156),
    .B(_06830_),
    .X(_06831_));
 sky130_fd_sc_hd__a22o_1 _14682_ (.A1(net9033),
    .A2(net2868),
    .B1(_06825_),
    .B2(net3617),
    .X(_00139_));
 sky130_fd_sc_hd__or4_2 _14683_ (.A(net7161),
    .B(net7165),
    .C(net7159),
    .D(net7157),
    .X(_06832_));
 sky130_fd_sc_hd__nand2_1 _14684_ (.A(net7454),
    .B(_06832_),
    .Y(_06833_));
 sky130_fd_sc_hd__xnor2_1 _14685_ (.A(\matmul0.sin[4] ),
    .B(_06833_),
    .Y(_06834_));
 sky130_fd_sc_hd__a22o_1 _14686_ (.A1(net9031),
    .A2(net2868),
    .B1(net2262),
    .B2(net2863),
    .X(_00140_));
 sky130_fd_sc_hd__nor2_1 _14687_ (.A(\matmul0.sin[4] ),
    .B(_06832_),
    .Y(_06835_));
 sky130_fd_sc_hd__or2_1 _14688_ (.A(_06826_),
    .B(_06835_),
    .X(_06836_));
 sky130_fd_sc_hd__xnor2_1 _14689_ (.A(net7155),
    .B(_06836_),
    .Y(_06837_));
 sky130_fd_sc_hd__a22o_1 _14690_ (.A1(net8994),
    .A2(net2868),
    .B1(net2262),
    .B2(net2261),
    .X(_00141_));
 sky130_fd_sc_hd__clkbuf_1 _14691_ (.A(net3630),
    .X(_06838_));
 sky130_fd_sc_hd__or3_1 _14692_ (.A(\matmul0.sin[4] ),
    .B(net7155),
    .C(_06832_),
    .X(_06839_));
 sky130_fd_sc_hd__nand2_1 _14693_ (.A(net7454),
    .B(_06839_),
    .Y(_06840_));
 sky130_fd_sc_hd__xnor2_1 _14694_ (.A(net7153),
    .B(_06840_),
    .Y(_06841_));
 sky130_fd_sc_hd__a22o_1 _14695_ (.A1(net9036),
    .A2(net2862),
    .B1(net2262),
    .B2(net2260),
    .X(_00142_));
 sky130_fd_sc_hd__or2_2 _14696_ (.A(net7153),
    .B(_06839_),
    .X(_06842_));
 sky130_fd_sc_hd__nand2_1 _14697_ (.A(net7453),
    .B(_06842_),
    .Y(_06843_));
 sky130_fd_sc_hd__xnor2_1 _14698_ (.A(net7152),
    .B(_06843_),
    .Y(_06844_));
 sky130_fd_sc_hd__a22o_1 _14699_ (.A1(net9094),
    .A2(net2862),
    .B1(net2262),
    .B2(net1910),
    .X(_00143_));
 sky130_fd_sc_hd__o21ai_1 _14700_ (.A1(net7152),
    .A2(_06842_),
    .B1(net7459),
    .Y(_06845_));
 sky130_fd_sc_hd__xnor2_1 _14701_ (.A(net7151),
    .B(_06845_),
    .Y(_06846_));
 sky130_fd_sc_hd__a22o_1 _14702_ (.A1(net9113),
    .A2(net2862),
    .B1(net2262),
    .B2(net1909),
    .X(_00144_));
 sky130_fd_sc_hd__or3_1 _14703_ (.A(net7152),
    .B(net7151),
    .C(_06842_),
    .X(_06847_));
 sky130_fd_sc_hd__nand2_1 _14704_ (.A(net7459),
    .B(_06847_),
    .Y(_06848_));
 sky130_fd_sc_hd__xnor2_1 _14705_ (.A(net7149),
    .B(_06848_),
    .Y(_06849_));
 sky130_fd_sc_hd__a22o_1 _14706_ (.A1(net9039),
    .A2(net2862),
    .B1(net2262),
    .B2(net1547),
    .X(_00145_));
 sky130_fd_sc_hd__or2_1 _14707_ (.A(net7149),
    .B(_06847_),
    .X(_06850_));
 sky130_fd_sc_hd__nand2_1 _14708_ (.A(net7456),
    .B(net1908),
    .Y(_06851_));
 sky130_fd_sc_hd__xnor2_1 _14709_ (.A(\matmul0.sin[10] ),
    .B(_06851_),
    .Y(_06852_));
 sky130_fd_sc_hd__a22o_1 _14710_ (.A1(net9082),
    .A2(net2861),
    .B1(net2263),
    .B2(net1290),
    .X(_00146_));
 sky130_fd_sc_hd__o21ai_1 _14711_ (.A1(\matmul0.sin[10] ),
    .A2(net1908),
    .B1(net7456),
    .Y(_06853_));
 sky130_fd_sc_hd__xnor2_1 _14712_ (.A(\matmul0.sin[11] ),
    .B(_06853_),
    .Y(_06854_));
 sky130_fd_sc_hd__a22o_1 _14713_ (.A1(net9130),
    .A2(net2861),
    .B1(net2263),
    .B2(net1288),
    .X(_00147_));
 sky130_fd_sc_hd__or3_1 _14714_ (.A(\matmul0.sin[10] ),
    .B(\matmul0.sin[11] ),
    .C(net1908),
    .X(_06855_));
 sky130_fd_sc_hd__nand2_1 _14715_ (.A(net7456),
    .B(_06855_),
    .Y(_06856_));
 sky130_fd_sc_hd__xnor2_1 _14716_ (.A(\matmul0.sin[12] ),
    .B(_06856_),
    .Y(_06857_));
 sky130_fd_sc_hd__a22o_1 _14717_ (.A1(net9092),
    .A2(net2861),
    .B1(net2865),
    .B2(net1118),
    .X(_00148_));
 sky130_fd_sc_hd__or2_1 _14718_ (.A(\matmul0.sin[12] ),
    .B(_06855_),
    .X(_06858_));
 sky130_fd_sc_hd__a21boi_1 _14719_ (.A1(net7457),
    .A2(_06858_),
    .B1_N(net7148),
    .Y(_06859_));
 sky130_fd_sc_hd__and3b_1 _14720_ (.A_N(net7148),
    .B(_06858_),
    .C(net7457),
    .X(_06860_));
 sky130_fd_sc_hd__o211a_1 _14721_ (.A1(_06859_),
    .A2(_06860_),
    .B1(net7441),
    .C1(net2876),
    .X(_06861_));
 sky130_fd_sc_hd__a21o_1 _14722_ (.A1(net8991),
    .A2(_06814_),
    .B1(_06861_),
    .X(_00149_));
 sky130_fd_sc_hd__clkbuf_1 _14723_ (.A(net4224),
    .X(_06862_));
 sky130_fd_sc_hd__a21o_1 _14724_ (.A1(net3613),
    .A2(net7148),
    .B1(_06860_),
    .X(_06863_));
 sky130_fd_sc_hd__nand2_1 _14725_ (.A(_06824_),
    .B(_06863_),
    .Y(_06864_));
 sky130_fd_sc_hd__a21bo_1 _14726_ (.A1(net9120),
    .A2(_06820_),
    .B1_N(net890),
    .X(_00150_));
 sky130_fd_sc_hd__a21bo_1 _14727_ (.A1(net8973),
    .A2(_06820_),
    .B1_N(net890),
    .X(_00151_));
 sky130_fd_sc_hd__and3_1 _14728_ (.A(net7437),
    .B(net7162),
    .C(net3697),
    .X(_06865_));
 sky130_fd_sc_hd__a21o_1 _14729_ (.A1(net8980),
    .A2(net2872),
    .B1(_06865_),
    .X(_00152_));
 sky130_fd_sc_hd__and3_1 _14730_ (.A(net3613),
    .B(net7160),
    .C(net7163),
    .X(_06866_));
 sky130_fd_sc_hd__o21ai_1 _14731_ (.A1(_06827_),
    .A2(_06866_),
    .B1(net7444),
    .Y(_06867_));
 sky130_fd_sc_hd__nand2_1 _14732_ (.A(net7444),
    .B(net7160),
    .Y(_06868_));
 sky130_fd_sc_hd__buf_1 _14733_ (.A(net3619),
    .X(_06869_));
 sky130_fd_sc_hd__a21oi_1 _14734_ (.A1(net7455),
    .A2(_06868_),
    .B1(net2859),
    .Y(_06870_));
 sky130_fd_sc_hd__a22o_1 _14735_ (.A1(net9071),
    .A2(net2860),
    .B1(_06867_),
    .B2(_06870_),
    .X(_00153_));
 sky130_fd_sc_hd__or2_1 _14736_ (.A(net7455),
    .B(_06827_),
    .X(_06871_));
 sky130_fd_sc_hd__xnor2_1 _14737_ (.A(net7158),
    .B(_06871_),
    .Y(_06872_));
 sky130_fd_sc_hd__a22o_1 _14738_ (.A1(net9104),
    .A2(net2861),
    .B1(net2865),
    .B2(_06872_),
    .X(_00154_));
 sky130_fd_sc_hd__inv_2 _14739_ (.A(_06832_),
    .Y(_06873_));
 sky130_fd_sc_hd__o311a_1 _14740_ (.A1(net7161),
    .A2(net7164),
    .A3(net7158),
    .B1(net7156),
    .C1(net3614),
    .X(_06874_));
 sky130_fd_sc_hd__o21ai_1 _14741_ (.A1(_06873_),
    .A2(_06874_),
    .B1(net7448),
    .Y(_06875_));
 sky130_fd_sc_hd__nand2_1 _14742_ (.A(net7448),
    .B(net7156),
    .Y(_06876_));
 sky130_fd_sc_hd__a21oi_1 _14743_ (.A1(net7453),
    .A2(_06876_),
    .B1(net2858),
    .Y(_06877_));
 sky130_fd_sc_hd__a22o_1 _14744_ (.A1(net9063),
    .A2(net2860),
    .B1(net2259),
    .B2(_06877_),
    .X(_00155_));
 sky130_fd_sc_hd__and3_1 _14745_ (.A(net3616),
    .B(\matmul0.sin[4] ),
    .C(_06832_),
    .X(_06878_));
 sky130_fd_sc_hd__o21ai_1 _14746_ (.A1(_06835_),
    .A2(_06878_),
    .B1(net7448),
    .Y(_06879_));
 sky130_fd_sc_hd__nand2_1 _14747_ (.A(net7448),
    .B(\matmul0.sin[4] ),
    .Y(_06880_));
 sky130_fd_sc_hd__a21oi_1 _14748_ (.A1(net7454),
    .A2(_06880_),
    .B1(net2857),
    .Y(_06881_));
 sky130_fd_sc_hd__a22o_1 _14749_ (.A1(net9017),
    .A2(net2857),
    .B1(_06879_),
    .B2(_06881_),
    .X(_00156_));
 sky130_fd_sc_hd__or3b_1 _14750_ (.A(net7454),
    .B(_06835_),
    .C_N(net7155),
    .X(_06882_));
 sky130_fd_sc_hd__nand2_1 _14751_ (.A(_06839_),
    .B(_06882_),
    .Y(_06883_));
 sky130_fd_sc_hd__nand2_1 _14752_ (.A(net7448),
    .B(net7155),
    .Y(_06884_));
 sky130_fd_sc_hd__a221o_1 _14753_ (.A1(net7448),
    .A2(_06883_),
    .B1(_06884_),
    .B2(net7454),
    .C1(net3621),
    .X(_06885_));
 sky130_fd_sc_hd__a21bo_1 _14754_ (.A1(net8974),
    .A2(net2870),
    .B1_N(net1906),
    .X(_00157_));
 sky130_fd_sc_hd__nand3_1 _14755_ (.A(_06826_),
    .B(net7153),
    .C(_06839_),
    .Y(_06886_));
 sky130_fd_sc_hd__nand2_1 _14756_ (.A(_06842_),
    .B(_06886_),
    .Y(_06887_));
 sky130_fd_sc_hd__nand2_1 _14757_ (.A(net7448),
    .B(net7153),
    .Y(_06888_));
 sky130_fd_sc_hd__a221o_1 _14758_ (.A1(net7448),
    .A2(_06887_),
    .B1(_06888_),
    .B2(net7454),
    .C1(net3621),
    .X(_06889_));
 sky130_fd_sc_hd__a21bo_1 _14759_ (.A1(net8955),
    .A2(net2867),
    .B1_N(_06889_),
    .X(_00158_));
 sky130_fd_sc_hd__and2_1 _14760_ (.A(net3615),
    .B(_06842_),
    .X(_06890_));
 sky130_fd_sc_hd__xor2_1 _14761_ (.A(net7152),
    .B(_06890_),
    .X(_06891_));
 sky130_fd_sc_hd__a22o_1 _14762_ (.A1(net9128),
    .A2(net2858),
    .B1(net2865),
    .B2(_06891_),
    .X(_00159_));
 sky130_fd_sc_hd__o21a_1 _14763_ (.A1(net7152),
    .A2(_06842_),
    .B1(net3615),
    .X(_06892_));
 sky130_fd_sc_hd__xor2_1 _14764_ (.A(net7151),
    .B(_06892_),
    .X(_06893_));
 sky130_fd_sc_hd__a22o_1 _14765_ (.A1(net9034),
    .A2(net2858),
    .B1(net2865),
    .B2(_06893_),
    .X(_00160_));
 sky130_fd_sc_hd__nand3_1 _14766_ (.A(_06826_),
    .B(net7149),
    .C(_06847_),
    .Y(_06894_));
 sky130_fd_sc_hd__nand2_1 _14767_ (.A(_06850_),
    .B(_06894_),
    .Y(_06895_));
 sky130_fd_sc_hd__nand2_1 _14768_ (.A(net7448),
    .B(net7149),
    .Y(_06896_));
 sky130_fd_sc_hd__a221o_1 _14769_ (.A1(net7448),
    .A2(_06895_),
    .B1(_06896_),
    .B2(net7459),
    .C1(net3621),
    .X(_06897_));
 sky130_fd_sc_hd__a21bo_1 _14770_ (.A1(net8954),
    .A2(net2867),
    .B1_N(_06897_),
    .X(_00161_));
 sky130_fd_sc_hd__and2_1 _14771_ (.A(net4224),
    .B(net1908),
    .X(_06898_));
 sky130_fd_sc_hd__xor2_1 _14772_ (.A(\matmul0.sin[10] ),
    .B(_06898_),
    .X(_06899_));
 sky130_fd_sc_hd__a22o_1 _14773_ (.A1(net9003),
    .A2(net2857),
    .B1(net2866),
    .B2(_06899_),
    .X(_00162_));
 sky130_fd_sc_hd__o21a_1 _14774_ (.A1(\matmul0.sin[10] ),
    .A2(net1908),
    .B1(net3616),
    .X(_06900_));
 sky130_fd_sc_hd__xor2_1 _14775_ (.A(\matmul0.sin[11] ),
    .B(_06900_),
    .X(_06901_));
 sky130_fd_sc_hd__a22o_1 _14776_ (.A1(net9040),
    .A2(net2857),
    .B1(net2866),
    .B2(_06901_),
    .X(_00163_));
 sky130_fd_sc_hd__and2_1 _14777_ (.A(net3616),
    .B(_06855_),
    .X(_06902_));
 sky130_fd_sc_hd__xnor2_1 _14778_ (.A(\matmul0.sin[12] ),
    .B(_06902_),
    .Y(_06903_));
 sky130_fd_sc_hd__o2bb2a_1 _14779_ (.A1_N(net2866),
    .A2_N(_06903_),
    .B1(net9116),
    .B2(net3001),
    .X(_00164_));
 sky130_fd_sc_hd__and2_1 _14780_ (.A(net4223),
    .B(_06858_),
    .X(_06904_));
 sky130_fd_sc_hd__a21oi_1 _14781_ (.A1(net7148),
    .A2(_06858_),
    .B1(_06817_),
    .Y(_06905_));
 sky130_fd_sc_hd__o32a_1 _14782_ (.A1(_06817_),
    .A2(net7148),
    .A3(_06904_),
    .B1(_06905_),
    .B2(net7457),
    .X(_06906_));
 sky130_fd_sc_hd__mux2_1 _14783_ (.A0(\matmul0.matmul_stage_inst.c[13] ),
    .A1(_06906_),
    .S(net3698),
    .X(_06907_));
 sky130_fd_sc_hd__clkbuf_1 _14784_ (.A(_06907_),
    .X(_00165_));
 sky130_fd_sc_hd__nor2_1 _14785_ (.A(_06818_),
    .B(net7148),
    .Y(_06908_));
 sky130_fd_sc_hd__nor2_1 _14786_ (.A(net3613),
    .B(_06908_),
    .Y(_06909_));
 sky130_fd_sc_hd__a211o_1 _14787_ (.A1(_06904_),
    .A2(_06908_),
    .B1(_06909_),
    .C1(net3627),
    .X(_06910_));
 sky130_fd_sc_hd__o21a_1 _14788_ (.A1(net9146),
    .A2(net3003),
    .B1(net992),
    .X(_00166_));
 sky130_fd_sc_hd__o21a_1 _14789_ (.A1(net9057),
    .A2(net3003),
    .B1(net992),
    .X(_00167_));
 sky130_fd_sc_hd__nand2_1 _14790_ (.A(_06818_),
    .B(net7457),
    .Y(_06911_));
 sky130_fd_sc_hd__o211a_1 _14791_ (.A1(net3624),
    .A2(\matmul0.cos[0] ),
    .B1(net2878),
    .C1(net2855),
    .X(_06912_));
 sky130_fd_sc_hd__a21o_1 _14792_ (.A1(net9007),
    .A2(net2871),
    .B1(_06912_),
    .X(_00168_));
 sky130_fd_sc_hd__or3_1 _14793_ (.A(net3624),
    .B(net7182),
    .C(net3618),
    .X(_06913_));
 sky130_fd_sc_hd__o21a_1 _14794_ (.A1(net9052),
    .A2(net3006),
    .B1(_06913_),
    .X(_00169_));
 sky130_fd_sc_hd__nor2_1 _14795_ (.A(net7441),
    .B(net3614),
    .Y(_06914_));
 sky130_fd_sc_hd__a21o_1 _14796_ (.A1(net7438),
    .A2(net7181),
    .B1(net2856),
    .X(_06915_));
 sky130_fd_sc_hd__o22a_1 _14797_ (.A1(net9069),
    .A2(net3005),
    .B1(net2853),
    .B2(_06915_),
    .X(_00170_));
 sky130_fd_sc_hd__and3_1 _14798_ (.A(net7445),
    .B(\matmul0.cos[3] ),
    .C(net3697),
    .X(_06916_));
 sky130_fd_sc_hd__a21o_1 _14799_ (.A1(net8981),
    .A2(net2871),
    .B1(_06916_),
    .X(_00171_));
 sky130_fd_sc_hd__or3_1 _14800_ (.A(net3624),
    .B(net7180),
    .C(net3618),
    .X(_06917_));
 sky130_fd_sc_hd__o21a_1 _14801_ (.A1(net9019),
    .A2(net3006),
    .B1(_06917_),
    .X(_00172_));
 sky130_fd_sc_hd__or3_1 _14802_ (.A(net3626),
    .B(net7178),
    .C(net3622),
    .X(_06918_));
 sky130_fd_sc_hd__o21a_1 _14803_ (.A1(net9020),
    .A2(net3004),
    .B1(_06918_),
    .X(_00173_));
 sky130_fd_sc_hd__o211a_1 _14804_ (.A1(net3625),
    .A2(\matmul0.cos[6] ),
    .B1(_06802_),
    .C1(net2855),
    .X(_06919_));
 sky130_fd_sc_hd__a21o_1 _14805_ (.A1(net9002),
    .A2(net2871),
    .B1(_06919_),
    .X(_00174_));
 sky130_fd_sc_hd__or3_1 _14806_ (.A(net3626),
    .B(net7175),
    .C(net3622),
    .X(_06920_));
 sky130_fd_sc_hd__o21a_1 _14807_ (.A1(net9008),
    .A2(net3004),
    .B1(_06920_),
    .X(_00175_));
 sky130_fd_sc_hd__a21o_1 _14808_ (.A1(net7442),
    .A2(net7172),
    .B1(net3628),
    .X(_06921_));
 sky130_fd_sc_hd__o22a_1 _14809_ (.A1(net9045),
    .A2(net3005),
    .B1(net2853),
    .B2(_06921_),
    .X(_00176_));
 sky130_fd_sc_hd__a21o_1 _14810_ (.A1(net7442),
    .A2(net7170),
    .B1(net3628),
    .X(_06922_));
 sky130_fd_sc_hd__o22a_1 _14811_ (.A1(net9065),
    .A2(net2876),
    .B1(net2854),
    .B2(_06922_),
    .X(_00177_));
 sky130_fd_sc_hd__o211a_1 _14812_ (.A1(net3625),
    .A2(net7169),
    .B1(_06802_),
    .C1(net2855),
    .X(_06923_));
 sky130_fd_sc_hd__a21o_1 _14813_ (.A1(net8978),
    .A2(net2871),
    .B1(_06923_),
    .X(_00178_));
 sky130_fd_sc_hd__a21o_1 _14814_ (.A1(net7446),
    .A2(net7168),
    .B1(net3627),
    .X(_06924_));
 sky130_fd_sc_hd__o22a_1 _14815_ (.A1(net9044),
    .A2(net2877),
    .B1(net2854),
    .B2(_06924_),
    .X(_00179_));
 sky130_fd_sc_hd__a21o_1 _14816_ (.A1(net7441),
    .A2(net7167),
    .B1(net3627),
    .X(_06925_));
 sky130_fd_sc_hd__o22a_1 _14817_ (.A1(net9026),
    .A2(net2877),
    .B1(net2854),
    .B2(_06925_),
    .X(_00180_));
 sky130_fd_sc_hd__a22o_1 _14818_ (.A1(net9087),
    .A2(_06869_),
    .B1(_06819_),
    .B2(_06911_),
    .X(_00181_));
 sky130_fd_sc_hd__and3_1 _14819_ (.A(net7438),
    .B(net7166),
    .C(_04884_),
    .X(_06926_));
 sky130_fd_sc_hd__a21o_1 _14820_ (.A1(net8984),
    .A2(net2872),
    .B1(_06926_),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _14821_ (.A0(net7183),
    .A1(\matmul0.matmul_stage_inst.e[0] ),
    .S(net3630),
    .X(_06927_));
 sky130_fd_sc_hd__clkbuf_1 _14822_ (.A(_06927_),
    .X(_00183_));
 sky130_fd_sc_hd__buf_1 _14823_ (.A(net4285),
    .X(_06928_));
 sky130_fd_sc_hd__mux2_1 _14824_ (.A0(\matmul0.a[1] ),
    .A1(\matmul0.matmul_stage_inst.e[1] ),
    .S(net3610),
    .X(_06929_));
 sky130_fd_sc_hd__clkbuf_1 _14825_ (.A(_06929_),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _14826_ (.A0(\matmul0.a[2] ),
    .A1(\matmul0.matmul_stage_inst.e[2] ),
    .S(net3610),
    .X(_06930_));
 sky130_fd_sc_hd__clkbuf_1 _14827_ (.A(_06930_),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _14828_ (.A0(\matmul0.a[3] ),
    .A1(\matmul0.matmul_stage_inst.e[3] ),
    .S(net3610),
    .X(_06931_));
 sky130_fd_sc_hd__clkbuf_1 _14829_ (.A(_06931_),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _14830_ (.A0(net9231),
    .A1(\matmul0.matmul_stage_inst.e[4] ),
    .S(net3610),
    .X(_06932_));
 sky130_fd_sc_hd__clkbuf_1 _14831_ (.A(_06932_),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _14832_ (.A0(\matmul0.a[5] ),
    .A1(\matmul0.matmul_stage_inst.e[5] ),
    .S(net3610),
    .X(_06933_));
 sky130_fd_sc_hd__clkbuf_1 _14833_ (.A(_06933_),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _14834_ (.A0(\matmul0.a[6] ),
    .A1(\matmul0.matmul_stage_inst.e[6] ),
    .S(net3611),
    .X(_06934_));
 sky130_fd_sc_hd__clkbuf_1 _14835_ (.A(_06934_),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _14836_ (.A0(\matmul0.a[7] ),
    .A1(\matmul0.matmul_stage_inst.e[7] ),
    .S(net3611),
    .X(_06935_));
 sky130_fd_sc_hd__clkbuf_1 _14837_ (.A(_06935_),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _14838_ (.A0(\matmul0.a[8] ),
    .A1(\matmul0.matmul_stage_inst.e[8] ),
    .S(_06928_),
    .X(_06936_));
 sky130_fd_sc_hd__clkbuf_1 _14839_ (.A(_06936_),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _14840_ (.A0(net9227),
    .A1(\matmul0.matmul_stage_inst.e[9] ),
    .S(net3612),
    .X(_06937_));
 sky130_fd_sc_hd__clkbuf_1 _14841_ (.A(_06937_),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _14842_ (.A0(\matmul0.a[10] ),
    .A1(\matmul0.matmul_stage_inst.e[10] ),
    .S(net3612),
    .X(_06938_));
 sky130_fd_sc_hd__clkbuf_1 _14843_ (.A(_06938_),
    .X(_00193_));
 sky130_fd_sc_hd__buf_1 _14844_ (.A(net4283),
    .X(_06939_));
 sky130_fd_sc_hd__mux2_1 _14845_ (.A0(\matmul0.a[11] ),
    .A1(\matmul0.matmul_stage_inst.e[11] ),
    .S(net3607),
    .X(_06940_));
 sky130_fd_sc_hd__clkbuf_1 _14846_ (.A(_06940_),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _14847_ (.A0(\matmul0.a[12] ),
    .A1(\matmul0.matmul_stage_inst.e[12] ),
    .S(net3607),
    .X(_06941_));
 sky130_fd_sc_hd__clkbuf_1 _14848_ (.A(_06941_),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _14849_ (.A0(net9183),
    .A1(\matmul0.matmul_stage_inst.e[13] ),
    .S(net3608),
    .X(_06942_));
 sky130_fd_sc_hd__clkbuf_1 _14850_ (.A(_06942_),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _14851_ (.A0(\matmul0.a[14] ),
    .A1(\matmul0.matmul_stage_inst.e[14] ),
    .S(net3607),
    .X(_06943_));
 sky130_fd_sc_hd__clkbuf_1 _14852_ (.A(_06943_),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _14853_ (.A0(\matmul0.a[15] ),
    .A1(\matmul0.matmul_stage_inst.e[15] ),
    .S(net3607),
    .X(_06944_));
 sky130_fd_sc_hd__clkbuf_1 _14854_ (.A(_06944_),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _14855_ (.A0(\matmul0.b[0] ),
    .A1(\matmul0.matmul_stage_inst.f[0] ),
    .S(net3609),
    .X(_06945_));
 sky130_fd_sc_hd__clkbuf_1 _14856_ (.A(_06945_),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _14857_ (.A0(net7190),
    .A1(\matmul0.matmul_stage_inst.f[1] ),
    .S(net3608),
    .X(_06946_));
 sky130_fd_sc_hd__clkbuf_1 _14858_ (.A(_06946_),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _14859_ (.A0(net7188),
    .A1(\matmul0.matmul_stage_inst.f[2] ),
    .S(_06939_),
    .X(_06947_));
 sky130_fd_sc_hd__clkbuf_1 _14860_ (.A(_06947_),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _14861_ (.A0(net7187),
    .A1(\matmul0.matmul_stage_inst.f[3] ),
    .S(net3609),
    .X(_06948_));
 sky130_fd_sc_hd__clkbuf_1 _14862_ (.A(_06948_),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _14863_ (.A0(net7186),
    .A1(\matmul0.matmul_stage_inst.f[4] ),
    .S(_06939_),
    .X(_06949_));
 sky130_fd_sc_hd__clkbuf_1 _14864_ (.A(_06949_),
    .X(_00203_));
 sky130_fd_sc_hd__buf_1 _14865_ (.A(net4284),
    .X(_06950_));
 sky130_fd_sc_hd__mux2_1 _14866_ (.A0(\matmul0.b[5] ),
    .A1(\matmul0.matmul_stage_inst.f[5] ),
    .S(net3606),
    .X(_06951_));
 sky130_fd_sc_hd__clkbuf_1 _14867_ (.A(_06951_),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _14868_ (.A0(\matmul0.b[6] ),
    .A1(\matmul0.matmul_stage_inst.f[6] ),
    .S(_06950_),
    .X(_06952_));
 sky130_fd_sc_hd__clkbuf_1 _14869_ (.A(_06952_),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _14870_ (.A0(net7185),
    .A1(\matmul0.matmul_stage_inst.f[7] ),
    .S(net3606),
    .X(_06953_));
 sky130_fd_sc_hd__clkbuf_1 _14871_ (.A(_06953_),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _14872_ (.A0(net7184),
    .A1(\matmul0.matmul_stage_inst.f[8] ),
    .S(net3606),
    .X(_06954_));
 sky130_fd_sc_hd__clkbuf_1 _14873_ (.A(_06954_),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _14874_ (.A0(\matmul0.b[9] ),
    .A1(\matmul0.matmul_stage_inst.f[9] ),
    .S(net3604),
    .X(_06955_));
 sky130_fd_sc_hd__clkbuf_1 _14875_ (.A(_06955_),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _14876_ (.A0(\matmul0.b[10] ),
    .A1(\matmul0.matmul_stage_inst.f[10] ),
    .S(net3604),
    .X(_06956_));
 sky130_fd_sc_hd__clkbuf_1 _14877_ (.A(_06956_),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _14878_ (.A0(net9225),
    .A1(\matmul0.matmul_stage_inst.f[11] ),
    .S(net3604),
    .X(_06957_));
 sky130_fd_sc_hd__clkbuf_1 _14879_ (.A(_06957_),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _14880_ (.A0(\matmul0.b[12] ),
    .A1(\matmul0.matmul_stage_inst.f[12] ),
    .S(net3604),
    .X(_06958_));
 sky130_fd_sc_hd__clkbuf_1 _14881_ (.A(_06958_),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _14882_ (.A0(net9237),
    .A1(\matmul0.matmul_stage_inst.f[13] ),
    .S(net3606),
    .X(_06959_));
 sky130_fd_sc_hd__clkbuf_1 _14883_ (.A(_06959_),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _14884_ (.A0(\matmul0.b[14] ),
    .A1(\matmul0.matmul_stage_inst.f[14] ),
    .S(net3605),
    .X(_06960_));
 sky130_fd_sc_hd__clkbuf_1 _14885_ (.A(_06960_),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _14886_ (.A0(\matmul0.b[15] ),
    .A1(\matmul0.matmul_stage_inst.f[15] ),
    .S(net3623),
    .X(_06961_));
 sky130_fd_sc_hd__clkbuf_1 _14887_ (.A(_06961_),
    .X(_00214_));
 sky130_fd_sc_hd__o21a_1 _14888_ (.A1(net6620),
    .A2(net6638),
    .B1(\matmul0.matmul_stage_inst.f[0] ),
    .X(_06962_));
 sky130_fd_sc_hd__o21a_1 _14889_ (.A1(net6539),
    .A2(net6590),
    .B1(\matmul0.matmul_stage_inst.e[0] ),
    .X(_06963_));
 sky130_fd_sc_hd__nor2_1 _14890_ (.A(net4221),
    .B(net4219),
    .Y(_06964_));
 sky130_fd_sc_hd__a22o_1 _14891_ (.A1(net6631),
    .A2(\matmul0.matmul_stage_inst.d[11] ),
    .B1(net7405),
    .B2(net6533),
    .X(_06965_));
 sky130_fd_sc_hd__a22o_1 _14892_ (.A1(net6611),
    .A2(\matmul0.matmul_stage_inst.b[11] ),
    .B1(\matmul0.matmul_stage_inst.a[11] ),
    .B2(net6581),
    .X(_06966_));
 sky130_fd_sc_hd__nor2_1 _14893_ (.A(net4216),
    .B(net4214),
    .Y(_06967_));
 sky130_fd_sc_hd__nor2_1 _14894_ (.A(net3602),
    .B(net3601),
    .Y(_06968_));
 sky130_fd_sc_hd__o21a_1 _14895_ (.A1(net6615),
    .A2(net6638),
    .B1(\matmul0.matmul_stage_inst.f[2] ),
    .X(_06969_));
 sky130_fd_sc_hd__o21a_1 _14896_ (.A1(net6543),
    .A2(net6588),
    .B1(net7396),
    .X(_06970_));
 sky130_fd_sc_hd__a22o_1 _14897_ (.A1(net6612),
    .A2(net7421),
    .B1(\matmul0.matmul_stage_inst.a[9] ),
    .B2(net6580),
    .X(_06971_));
 sky130_fd_sc_hd__a22o_1 _14898_ (.A1(net6631),
    .A2(\matmul0.matmul_stage_inst.d[9] ),
    .B1(net7408),
    .B2(net6533),
    .X(_06972_));
 sky130_fd_sc_hd__o22a_1 _14899_ (.A1(net4213),
    .A2(net4211),
    .B1(net4210),
    .B2(net4208),
    .X(_06973_));
 sky130_fd_sc_hd__o21a_1 _14900_ (.A1(net6620),
    .A2(net6644),
    .B1(\matmul0.matmul_stage_inst.f[1] ),
    .X(_06974_));
 sky130_fd_sc_hd__o21a_1 _14901_ (.A1(net6542),
    .A2(net6586),
    .B1(net7398),
    .X(_06975_));
 sky130_fd_sc_hd__a22o_1 _14902_ (.A1(net6630),
    .A2(\matmul0.matmul_stage_inst.d[10] ),
    .B1(net7406),
    .B2(net6532),
    .X(_06976_));
 sky130_fd_sc_hd__a22o_1 _14903_ (.A1(net6612),
    .A2(net7420),
    .B1(\matmul0.matmul_stage_inst.a[10] ),
    .B2(net6583),
    .X(_06977_));
 sky130_fd_sc_hd__o22a_1 _14904_ (.A1(net4207),
    .A2(net4203),
    .B1(net4198),
    .B2(net4197),
    .X(_06978_));
 sky130_fd_sc_hd__xnor2_1 _14905_ (.A(net3598),
    .B(_06978_),
    .Y(_06979_));
 sky130_fd_sc_hd__xnor2_1 _14906_ (.A(_06968_),
    .B(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__o22a_1 _14907_ (.A1(net4206),
    .A2(net4202),
    .B1(net4210),
    .B2(net4208),
    .X(_06981_));
 sky130_fd_sc_hd__a22o_1 _14908_ (.A1(net6636),
    .A2(\matmul0.matmul_stage_inst.d[8] ),
    .B1(net7410),
    .B2(net6531),
    .X(_06982_));
 sky130_fd_sc_hd__a22o_1 _14909_ (.A1(net6614),
    .A2(net7423),
    .B1(\matmul0.matmul_stage_inst.a[8] ),
    .B2(net6585),
    .X(_06983_));
 sky130_fd_sc_hd__clkbuf_1 _14910_ (.A(_06969_),
    .X(_06984_));
 sky130_fd_sc_hd__clkbuf_1 _14911_ (.A(net4212),
    .X(_06985_));
 sky130_fd_sc_hd__o22a_1 _14912_ (.A1(net4196),
    .A2(net4194),
    .B1(net3595),
    .B2(net3593),
    .X(_06986_));
 sky130_fd_sc_hd__or2_1 _14913_ (.A(net4222),
    .B(net4220),
    .X(_06987_));
 sky130_fd_sc_hd__buf_1 _14914_ (.A(_06987_),
    .X(_06988_));
 sky130_fd_sc_hd__or2_1 _14915_ (.A(net4198),
    .B(net4197),
    .X(_06989_));
 sky130_fd_sc_hd__a22o_1 _14916_ (.A1(_06988_),
    .A2(_06989_),
    .B1(_06981_),
    .B2(_06986_),
    .X(_06990_));
 sky130_fd_sc_hd__o21a_1 _14917_ (.A1(_06981_),
    .A2(_06986_),
    .B1(_06990_),
    .X(_06991_));
 sky130_fd_sc_hd__o21a_1 _14918_ (.A1(net6619),
    .A2(net6644),
    .B1(net7385),
    .X(_06992_));
 sky130_fd_sc_hd__o21a_1 _14919_ (.A1(net6556),
    .A2(net6587),
    .B1(\matmul0.matmul_stage_inst.e[5] ),
    .X(_06993_));
 sky130_fd_sc_hd__a22o_1 _14920_ (.A1(net6630),
    .A2(\matmul0.matmul_stage_inst.d[6] ),
    .B1(net7411),
    .B2(net6532),
    .X(_06994_));
 sky130_fd_sc_hd__a22o_1 _14921_ (.A1(net6610),
    .A2(net7425),
    .B1(\matmul0.matmul_stage_inst.a[6] ),
    .B2(net6583),
    .X(_06995_));
 sky130_fd_sc_hd__o22a_1 _14922_ (.A1(net4192),
    .A2(net4187),
    .B1(net4182),
    .B2(net4180),
    .X(_06996_));
 sky130_fd_sc_hd__o21a_1 _14923_ (.A1(net6613),
    .A2(net6638),
    .B1(\matmul0.matmul_stage_inst.f[4] ),
    .X(_06997_));
 sky130_fd_sc_hd__o21a_1 _14924_ (.A1(net6545),
    .A2(net6585),
    .B1(net7392),
    .X(_06998_));
 sky130_fd_sc_hd__a22o_1 _14925_ (.A1(net6627),
    .A2(\matmul0.matmul_stage_inst.d[7] ),
    .B1(\matmul0.matmul_stage_inst.c[7] ),
    .B2(net6535),
    .X(_06999_));
 sky130_fd_sc_hd__a22o_1 _14926_ (.A1(net6609),
    .A2(net7424),
    .B1(\matmul0.matmul_stage_inst.a[7] ),
    .B2(net6585),
    .X(_07000_));
 sky130_fd_sc_hd__o22a_1 _14927_ (.A1(net4178),
    .A2(_06998_),
    .B1(net4177),
    .B2(_07000_),
    .X(_07001_));
 sky130_fd_sc_hd__o21a_1 _14928_ (.A1(net6619),
    .A2(net6644),
    .B1(\matmul0.matmul_stage_inst.f[3] ),
    .X(_07002_));
 sky130_fd_sc_hd__o21a_1 _14929_ (.A1(net6559),
    .A2(net6587),
    .B1(\matmul0.matmul_stage_inst.e[3] ),
    .X(_07003_));
 sky130_fd_sc_hd__o22a_1 _14930_ (.A1(net4171),
    .A2(net4167),
    .B1(net4196),
    .B2(net4194),
    .X(_07004_));
 sky130_fd_sc_hd__xnor2_1 _14931_ (.A(_07001_),
    .B(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__xnor2_1 _14932_ (.A(_06996_),
    .B(_07005_),
    .Y(_07006_));
 sky130_fd_sc_hd__xnor2_1 _14933_ (.A(net1902),
    .B(net2252),
    .Y(_07007_));
 sky130_fd_sc_hd__xnor2_2 _14934_ (.A(net2256),
    .B(_07007_),
    .Y(_07008_));
 sky130_fd_sc_hd__a22o_1 _14935_ (.A1(net6635),
    .A2(\matmul0.matmul_stage_inst.d[5] ),
    .B1(net7413),
    .B2(net6535),
    .X(_07009_));
 sky130_fd_sc_hd__a22o_1 _14936_ (.A1(net6611),
    .A2(net7427),
    .B1(\matmul0.matmul_stage_inst.a[5] ),
    .B2(net6585),
    .X(_07010_));
 sky130_fd_sc_hd__or2_1 _14937_ (.A(net4161),
    .B(net4157),
    .X(_07011_));
 sky130_fd_sc_hd__buf_1 _14938_ (.A(_07011_),
    .X(_07012_));
 sky130_fd_sc_hd__o21a_1 _14939_ (.A1(net6619),
    .A2(net6644),
    .B1(net7384),
    .X(_07013_));
 sky130_fd_sc_hd__o21a_1 _14940_ (.A1(net6536),
    .A2(net6588),
    .B1(\matmul0.matmul_stage_inst.e[6] ),
    .X(_07014_));
 sky130_fd_sc_hd__or2_1 _14941_ (.A(net4153),
    .B(net4148),
    .X(_07015_));
 sky130_fd_sc_hd__buf_1 _14942_ (.A(_07015_),
    .X(_07016_));
 sky130_fd_sc_hd__nand2_1 _14943_ (.A(_07012_),
    .B(_07016_),
    .Y(_07017_));
 sky130_fd_sc_hd__o21a_1 _14944_ (.A1(net6634),
    .A2(net6582),
    .B1(net7404),
    .X(_07018_));
 sky130_fd_sc_hd__buf_1 _14945_ (.A(_07018_),
    .X(_07019_));
 sky130_fd_sc_hd__a22o_1 _14946_ (.A1(net6537),
    .A2(\matmul0.matmul_stage_inst.c[3] ),
    .B1(\matmul0.matmul_stage_inst.b[3] ),
    .B2(net6617),
    .X(_07020_));
 sky130_fd_sc_hd__clkbuf_1 _14947_ (.A(net4146),
    .X(_07021_));
 sky130_fd_sc_hd__o21a_1 _14948_ (.A1(net6620),
    .A2(net6640),
    .B1(\matmul0.matmul_stage_inst.f[8] ),
    .X(_07022_));
 sky130_fd_sc_hd__o21a_1 _14949_ (.A1(net6543),
    .A2(net6588),
    .B1(net7391),
    .X(_07023_));
 sky130_fd_sc_hd__o22a_1 _14950_ (.A1(net3582),
    .A2(net3580),
    .B1(net4143),
    .B2(net4140),
    .X(_07024_));
 sky130_fd_sc_hd__a22o_1 _14951_ (.A1(net6630),
    .A2(\matmul0.matmul_stage_inst.d[4] ),
    .B1(net7414),
    .B2(net6532),
    .X(_07025_));
 sky130_fd_sc_hd__buf_1 _14952_ (.A(net4139),
    .X(_07026_));
 sky130_fd_sc_hd__a22o_1 _14953_ (.A1(net6610),
    .A2(net7429),
    .B1(\matmul0.matmul_stage_inst.a[4] ),
    .B2(net6582),
    .X(_07027_));
 sky130_fd_sc_hd__buf_1 _14954_ (.A(_07027_),
    .X(_07028_));
 sky130_fd_sc_hd__o21a_1 _14955_ (.A1(net6620),
    .A2(net6640),
    .B1(\matmul0.matmul_stage_inst.f[7] ),
    .X(_07029_));
 sky130_fd_sc_hd__o21a_1 _14956_ (.A1(net6559),
    .A2(net6587),
    .B1(\matmul0.matmul_stage_inst.e[7] ),
    .X(_07030_));
 sky130_fd_sc_hd__o22a_1 _14957_ (.A1(net3575),
    .A2(net3571),
    .B1(net4137),
    .B2(net4130),
    .X(_07031_));
 sky130_fd_sc_hd__xnor2_1 _14958_ (.A(_07024_),
    .B(_07031_),
    .Y(_07032_));
 sky130_fd_sc_hd__xnor2_1 _14959_ (.A(_07017_),
    .B(_07032_),
    .Y(_07033_));
 sky130_fd_sc_hd__o22a_1 _14960_ (.A1(_07018_),
    .A2(net4146),
    .B1(net4139),
    .B2(_07027_),
    .X(_07034_));
 sky130_fd_sc_hd__o22a_1 _14961_ (.A1(_07029_),
    .A2(net4132),
    .B1(_07013_),
    .B2(net4151),
    .X(_07035_));
 sky130_fd_sc_hd__a22o_1 _14962_ (.A1(net6634),
    .A2(\matmul0.matmul_stage_inst.d[2] ),
    .B1(net7417),
    .B2(net6538),
    .X(_07036_));
 sky130_fd_sc_hd__a22o_1 _14963_ (.A1(net6612),
    .A2(net7432),
    .B1(\matmul0.matmul_stage_inst.a[2] ),
    .B2(net6583),
    .X(_07037_));
 sky130_fd_sc_hd__nor2_1 _14964_ (.A(net4126),
    .B(net4124),
    .Y(_07038_));
 sky130_fd_sc_hd__nor2_1 _14965_ (.A(net4143),
    .B(net4140),
    .Y(_07039_));
 sky130_fd_sc_hd__o2bb2a_1 _14966_ (.A1_N(net3567),
    .A2_N(net3562),
    .B1(net3560),
    .B2(net3558),
    .X(_07040_));
 sky130_fd_sc_hd__nor2_1 _14967_ (.A(net3584),
    .B(net3577),
    .Y(_07041_));
 sky130_fd_sc_hd__nor2_1 _14968_ (.A(net4136),
    .B(net4129),
    .Y(_07042_));
 sky130_fd_sc_hd__nor2_1 _14969_ (.A(net4154),
    .B(net4149),
    .Y(_07043_));
 sky130_fd_sc_hd__nor2_1 _14970_ (.A(net4139),
    .B(_07027_),
    .Y(_07044_));
 sky130_fd_sc_hd__o22a_1 _14971_ (.A1(net2834),
    .A2(net3555),
    .B1(net3553),
    .B2(net3545),
    .X(_07045_));
 sky130_fd_sc_hd__nor2_1 _14972_ (.A(net2839),
    .B(_07045_),
    .Y(_07046_));
 sky130_fd_sc_hd__o22a_1 _14973_ (.A1(net4191),
    .A2(net4185),
    .B1(net4162),
    .B2(net4158),
    .X(_07047_));
 sky130_fd_sc_hd__o22a_1 _14974_ (.A1(net4178),
    .A2(_06998_),
    .B1(net4182),
    .B2(net4180),
    .X(_07048_));
 sky130_fd_sc_hd__o22a_1 _14975_ (.A1(net4170),
    .A2(net4165),
    .B1(net4175),
    .B2(net4173),
    .X(_07049_));
 sky130_fd_sc_hd__a21oi_1 _14976_ (.A1(net3544),
    .A2(net3541),
    .B1(net3539),
    .Y(_07050_));
 sky130_fd_sc_hd__nor2_1 _14977_ (.A(net3544),
    .B(net3541),
    .Y(_07051_));
 sky130_fd_sc_hd__nor2_1 _14978_ (.A(_07050_),
    .B(_07051_),
    .Y(_07052_));
 sky130_fd_sc_hd__xnor2_1 _14979_ (.A(_07046_),
    .B(_07052_),
    .Y(_07053_));
 sky130_fd_sc_hd__xnor2_1 _14980_ (.A(net1901),
    .B(_07053_),
    .Y(_07054_));
 sky130_fd_sc_hd__nor2_1 _14981_ (.A(net4198),
    .B(net4197),
    .Y(_07055_));
 sky130_fd_sc_hd__nor2_1 _14982_ (.A(net3603),
    .B(_07055_),
    .Y(_07056_));
 sky130_fd_sc_hd__xnor2_1 _14983_ (.A(_06981_),
    .B(_06986_),
    .Y(_07057_));
 sky130_fd_sc_hd__xnor2_1 _14984_ (.A(_07056_),
    .B(_07057_),
    .Y(_07058_));
 sky130_fd_sc_hd__xnor2_1 _14985_ (.A(net3539),
    .B(net3541),
    .Y(_07059_));
 sky130_fd_sc_hd__xnor2_2 _14986_ (.A(net3544),
    .B(_07059_),
    .Y(_07060_));
 sky130_fd_sc_hd__nor2_1 _14987_ (.A(net4195),
    .B(net4193),
    .Y(_07061_));
 sky130_fd_sc_hd__nor2_1 _14988_ (.A(net4206),
    .B(net4202),
    .Y(_07062_));
 sky130_fd_sc_hd__or2_1 _14989_ (.A(net4210),
    .B(net4208),
    .X(_07063_));
 sky130_fd_sc_hd__o22a_1 _14990_ (.A1(net4213),
    .A2(net4211),
    .B1(net4175),
    .B2(net4173),
    .X(_07064_));
 sky130_fd_sc_hd__a21oi_1 _14991_ (.A1(net2850),
    .A2(net3525),
    .B1(_07064_),
    .Y(_07065_));
 sky130_fd_sc_hd__nor2_1 _14992_ (.A(net4210),
    .B(net4208),
    .Y(_07066_));
 sky130_fd_sc_hd__or3b_1 _14993_ (.A(net3603),
    .B(net3521),
    .C_N(_07064_),
    .X(_07067_));
 sky130_fd_sc_hd__o31a_1 _14994_ (.A1(net3536),
    .A2(net3529),
    .A3(_07065_),
    .B1(_07067_),
    .X(_07068_));
 sky130_fd_sc_hd__o21bai_1 _14995_ (.A1(net1898),
    .A2(_07060_),
    .B1_N(net1896),
    .Y(_07069_));
 sky130_fd_sc_hd__a21bo_1 _14996_ (.A1(net1898),
    .A2(_07060_),
    .B1_N(_07069_),
    .X(_07070_));
 sky130_fd_sc_hd__xnor2_1 _14997_ (.A(net1287),
    .B(net1286),
    .Y(_07071_));
 sky130_fd_sc_hd__xnor2_1 _14998_ (.A(_07008_),
    .B(_07071_),
    .Y(_07072_));
 sky130_fd_sc_hd__inv_2 _14999_ (.A(_07072_),
    .Y(_07073_));
 sky130_fd_sc_hd__xor2_1 _15000_ (.A(net1896),
    .B(_07060_),
    .X(_07074_));
 sky130_fd_sc_hd__xnor2_2 _15001_ (.A(net1898),
    .B(_07074_),
    .Y(_07075_));
 sky130_fd_sc_hd__nor2_1 _15002_ (.A(_07038_),
    .B(net3558),
    .Y(_07076_));
 sky130_fd_sc_hd__or2_1 _15003_ (.A(net3584),
    .B(net3577),
    .X(_07077_));
 sky130_fd_sc_hd__or2_1 _15004_ (.A(net4136),
    .B(net4129),
    .X(_07078_));
 sky130_fd_sc_hd__a211o_1 _15005_ (.A1(net2831),
    .A2(_07078_),
    .B1(net3553),
    .C1(net3545),
    .X(_07079_));
 sky130_fd_sc_hd__or2_1 _15006_ (.A(net3573),
    .B(net3569),
    .X(_07080_));
 sky130_fd_sc_hd__a211o_1 _15007_ (.A1(net2827),
    .A2(_07015_),
    .B1(net3555),
    .C1(net2834),
    .X(_07081_));
 sky130_fd_sc_hd__and3_1 _15008_ (.A(_07076_),
    .B(_07079_),
    .C(_07081_),
    .X(_07082_));
 sky130_fd_sc_hd__a21oi_1 _15009_ (.A1(_07079_),
    .A2(_07081_),
    .B1(_07076_),
    .Y(_07083_));
 sky130_fd_sc_hd__or2_1 _15010_ (.A(_07082_),
    .B(_07083_),
    .X(_07084_));
 sky130_fd_sc_hd__o22a_1 _15011_ (.A1(net3582),
    .A2(net3580),
    .B1(net4153),
    .B2(net4148),
    .X(_07085_));
 sky130_fd_sc_hd__or2_1 _15012_ (.A(net4126),
    .B(net4124),
    .X(_07086_));
 sky130_fd_sc_hd__buf_1 _15013_ (.A(_07086_),
    .X(_07087_));
 sky130_fd_sc_hd__a22o_1 _15014_ (.A1(net6629),
    .A2(\matmul0.matmul_stage_inst.d[1] ),
    .B1(net7418),
    .B2(net6534),
    .X(_07088_));
 sky130_fd_sc_hd__a22o_1 _15015_ (.A1(net6610),
    .A2(net7434),
    .B1(\matmul0.matmul_stage_inst.a[1] ),
    .B2(net6582),
    .X(_07089_));
 sky130_fd_sc_hd__o22a_1 _15016_ (.A1(net4143),
    .A2(net4140),
    .B1(net4122),
    .B2(net4117),
    .X(_07090_));
 sky130_fd_sc_hd__a21o_1 _15017_ (.A1(net2826),
    .A2(_07078_),
    .B1(_07090_),
    .X(_07091_));
 sky130_fd_sc_hd__clkbuf_1 _15018_ (.A(_07078_),
    .X(_07092_));
 sky130_fd_sc_hd__and3_1 _15019_ (.A(net2826),
    .B(_07092_),
    .C(_07090_),
    .X(_07093_));
 sky130_fd_sc_hd__a21o_1 _15020_ (.A1(_07085_),
    .A2(_07091_),
    .B1(_07093_),
    .X(_07094_));
 sky130_fd_sc_hd__buf_1 _15021_ (.A(net4178),
    .X(_07095_));
 sky130_fd_sc_hd__buf_1 _15022_ (.A(_06998_),
    .X(_07096_));
 sky130_fd_sc_hd__o22a_1 _15023_ (.A1(net3511),
    .A2(net3506),
    .B1(net4163),
    .B2(net4159),
    .X(_07097_));
 sky130_fd_sc_hd__o22a_1 _15024_ (.A1(net4190),
    .A2(net4184),
    .B1(_07026_),
    .B2(_07028_),
    .X(_07098_));
 sky130_fd_sc_hd__or2_1 _15025_ (.A(net4171),
    .B(net4167),
    .X(_07099_));
 sky130_fd_sc_hd__clkbuf_1 _15026_ (.A(_07099_),
    .X(_07100_));
 sky130_fd_sc_hd__or2_1 _15027_ (.A(net4181),
    .B(net4179),
    .X(_07101_));
 sky130_fd_sc_hd__o211a_1 _15028_ (.A1(_07097_),
    .A2(_07098_),
    .B1(net2809),
    .C1(_07101_),
    .X(_07102_));
 sky130_fd_sc_hd__a21o_1 _15029_ (.A1(_07097_),
    .A2(_07098_),
    .B1(_07102_),
    .X(_07103_));
 sky130_fd_sc_hd__xnor2_1 _15030_ (.A(_07094_),
    .B(net1895),
    .Y(_07104_));
 sky130_fd_sc_hd__xnor2_1 _15031_ (.A(_07084_),
    .B(_07104_),
    .Y(_07105_));
 sky130_fd_sc_hd__nor2_1 _15032_ (.A(net4171),
    .B(net4166),
    .Y(_07106_));
 sky130_fd_sc_hd__nor2_1 _15033_ (.A(net4181),
    .B(net4179),
    .Y(_07107_));
 sky130_fd_sc_hd__clkbuf_1 _15034_ (.A(net3495),
    .X(_07108_));
 sky130_fd_sc_hd__nor2_1 _15035_ (.A(net3496),
    .B(net2808),
    .Y(_07109_));
 sky130_fd_sc_hd__xnor2_1 _15036_ (.A(_07097_),
    .B(_07098_),
    .Y(_07110_));
 sky130_fd_sc_hd__xnor2_2 _15037_ (.A(_07109_),
    .B(_07110_),
    .Y(_07111_));
 sky130_fd_sc_hd__nor2_1 _15038_ (.A(_06964_),
    .B(net3521),
    .Y(_07112_));
 sky130_fd_sc_hd__o22a_1 _15039_ (.A1(net4195),
    .A2(net4193),
    .B1(net4205),
    .B2(net4204),
    .X(_07113_));
 sky130_fd_sc_hd__xnor2_1 _15040_ (.A(_07064_),
    .B(_07113_),
    .Y(_07114_));
 sky130_fd_sc_hd__xnor2_1 _15041_ (.A(_07112_),
    .B(_07114_),
    .Y(_07115_));
 sky130_fd_sc_hd__o22a_1 _15042_ (.A1(net4181),
    .A2(net4180),
    .B1(net3595),
    .B2(net3593),
    .X(_07116_));
 sky130_fd_sc_hd__o22a_1 _15043_ (.A1(net4176),
    .A2(net4174),
    .B1(net4205),
    .B2(net4204),
    .X(_07117_));
 sky130_fd_sc_hd__or2_1 _15044_ (.A(net4195),
    .B(net4193),
    .X(_07118_));
 sky130_fd_sc_hd__a22o_1 _15045_ (.A1(net2850),
    .A2(_07118_),
    .B1(_07116_),
    .B2(_07117_),
    .X(_07119_));
 sky130_fd_sc_hd__o21a_1 _15046_ (.A1(_07116_),
    .A2(_07117_),
    .B1(_07119_),
    .X(_07120_));
 sky130_fd_sc_hd__o21a_1 _15047_ (.A1(_07111_),
    .A2(_07115_),
    .B1(_07120_),
    .X(_07121_));
 sky130_fd_sc_hd__a21oi_1 _15048_ (.A1(_07111_),
    .A2(_07115_),
    .B1(_07121_),
    .Y(_07122_));
 sky130_fd_sc_hd__o21ba_1 _15049_ (.A1(_07075_),
    .A2(net1285),
    .B1_N(net1283),
    .X(_07123_));
 sky130_fd_sc_hd__a21o_1 _15050_ (.A1(_07075_),
    .A2(net1285),
    .B1(_07123_),
    .X(_07124_));
 sky130_fd_sc_hd__buf_1 _15051_ (.A(net3560),
    .X(_07125_));
 sky130_fd_sc_hd__a22o_1 _15052_ (.A1(net6629),
    .A2(\matmul0.matmul_stage_inst.d[0] ),
    .B1(\matmul0.matmul_stage_inst.a[0] ),
    .B2(net6582),
    .X(_07126_));
 sky130_fd_sc_hd__o21a_1 _15053_ (.A1(net6610),
    .A2(net6534),
    .B1(\matmul0.matmul_stage_inst.b[0] ),
    .X(_07127_));
 sky130_fd_sc_hd__or2_1 _15054_ (.A(_07126_),
    .B(_07127_),
    .X(_07128_));
 sky130_fd_sc_hd__buf_1 _15055_ (.A(_07128_),
    .X(_07129_));
 sky130_fd_sc_hd__clkbuf_1 _15056_ (.A(net2794),
    .X(_07130_));
 sky130_fd_sc_hd__o21a_1 _15057_ (.A1(net6622),
    .A2(net6639),
    .B1(\matmul0.matmul_stage_inst.f[9] ),
    .X(_07131_));
 sky130_fd_sc_hd__o21a_1 _15058_ (.A1(net6547),
    .A2(net6592),
    .B1(net7389),
    .X(_07132_));
 sky130_fd_sc_hd__or2_1 _15059_ (.A(net4105),
    .B(net4101),
    .X(_07133_));
 sky130_fd_sc_hd__buf_1 _15060_ (.A(_07133_),
    .X(_07134_));
 sky130_fd_sc_hd__or2_1 _15061_ (.A(net6540),
    .B(net6592),
    .X(_07135_));
 sky130_fd_sc_hd__or2_1 _15062_ (.A(net6618),
    .B(net6639),
    .X(_07136_));
 sky130_fd_sc_hd__a22o_1 _15063_ (.A1(\matmul0.matmul_stage_inst.e[11] ),
    .A2(_07135_),
    .B1(_07136_),
    .B2(net7382),
    .X(_07137_));
 sky130_fd_sc_hd__clkbuf_1 _15064_ (.A(net3488),
    .X(_07138_));
 sky130_fd_sc_hd__or2_1 _15065_ (.A(net4120),
    .B(net4115),
    .X(_07139_));
 sky130_fd_sc_hd__buf_1 _15066_ (.A(_07139_),
    .X(_07140_));
 sky130_fd_sc_hd__nor2_1 _15067_ (.A(net4111),
    .B(net4108),
    .Y(_07141_));
 sky130_fd_sc_hd__buf_1 _15068_ (.A(net3486),
    .X(_07142_));
 sky130_fd_sc_hd__o21a_1 _15069_ (.A1(net6622),
    .A2(net6639),
    .B1(net7383),
    .X(_07143_));
 sky130_fd_sc_hd__o21a_1 _15070_ (.A1(net6546),
    .A2(net6594),
    .B1(net7386),
    .X(_07144_));
 sky130_fd_sc_hd__or2_1 _15071_ (.A(net4098),
    .B(net4096),
    .X(_07145_));
 sky130_fd_sc_hd__buf_1 _15072_ (.A(_07145_),
    .X(_07146_));
 sky130_fd_sc_hd__and3_1 _15073_ (.A(net2780),
    .B(net2776),
    .C(_07146_),
    .X(_07147_));
 sky130_fd_sc_hd__a31o_1 _15074_ (.A1(net2251),
    .A2(net2790),
    .A3(net2789),
    .B1(_07147_),
    .X(_07148_));
 sky130_fd_sc_hd__nor2_1 _15075_ (.A(net4120),
    .B(net4115),
    .Y(_07149_));
 sky130_fd_sc_hd__nor2_1 _15076_ (.A(net4099),
    .B(net4096),
    .Y(_07150_));
 sky130_fd_sc_hd__clkbuf_2 _15077_ (.A(_07135_),
    .X(_07151_));
 sky130_fd_sc_hd__clkbuf_2 _15078_ (.A(_07136_),
    .X(_07152_));
 sky130_fd_sc_hd__a22oi_1 _15079_ (.A1(\matmul0.matmul_stage_inst.e[11] ),
    .A2(_07151_),
    .B1(_07152_),
    .B2(net7382),
    .Y(_07153_));
 sky130_fd_sc_hd__o22a_1 _15080_ (.A1(_07149_),
    .A2(net3483),
    .B1(net2768),
    .B2(net3486),
    .X(_07154_));
 sky130_fd_sc_hd__and4_1 _15081_ (.A(net2781),
    .B(net2795),
    .C(_07145_),
    .D(net3489),
    .X(_07155_));
 sky130_fd_sc_hd__buf_1 _15082_ (.A(net2765),
    .X(_07156_));
 sky130_fd_sc_hd__nor2_1 _15083_ (.A(net4105),
    .B(net4101),
    .Y(_07157_));
 sky130_fd_sc_hd__nor2_1 _15084_ (.A(net3559),
    .B(_07157_),
    .Y(_07158_));
 sky130_fd_sc_hd__o21ai_1 _15085_ (.A1(net2778),
    .A2(net2243),
    .B1(_07158_),
    .Y(_07159_));
 sky130_fd_sc_hd__o32a_1 _15086_ (.A1(net2790),
    .A2(_07154_),
    .A3(_07155_),
    .B1(_07147_),
    .B2(_07159_),
    .X(_07160_));
 sky130_fd_sc_hd__a21bo_1 _15087_ (.A1(net2800),
    .A2(_07148_),
    .B1_N(_07160_),
    .X(_07161_));
 sky130_fd_sc_hd__o21a_1 _15088_ (.A1(_07094_),
    .A2(net1895),
    .B1(_07084_),
    .X(_07162_));
 sky130_fd_sc_hd__a21o_1 _15089_ (.A1(_07094_),
    .A2(net1895),
    .B1(_07162_),
    .X(_07163_));
 sky130_fd_sc_hd__xnor2_1 _15090_ (.A(net1280),
    .B(net1117),
    .Y(_07164_));
 sky130_fd_sc_hd__xnor2_1 _15091_ (.A(_07124_),
    .B(_07164_),
    .Y(_07165_));
 sky130_fd_sc_hd__xnor2_1 _15092_ (.A(_07073_),
    .B(_07165_),
    .Y(_07166_));
 sky130_fd_sc_hd__xnor2_1 _15093_ (.A(net1285),
    .B(net1283),
    .Y(_07167_));
 sky130_fd_sc_hd__xnor2_1 _15094_ (.A(_07075_),
    .B(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__nor2_1 _15095_ (.A(_07125_),
    .B(_07042_),
    .Y(_07169_));
 sky130_fd_sc_hd__xnor2_1 _15096_ (.A(_07085_),
    .B(_07090_),
    .Y(_07170_));
 sky130_fd_sc_hd__xnor2_1 _15097_ (.A(_07169_),
    .B(_07170_),
    .Y(_07171_));
 sky130_fd_sc_hd__o22a_1 _15098_ (.A1(net3511),
    .A2(net3506),
    .B1(_07026_),
    .B2(_07028_),
    .X(_07172_));
 sky130_fd_sc_hd__o22a_1 _15099_ (.A1(net4163),
    .A2(net4159),
    .B1(net4169),
    .B2(net4164),
    .X(_07173_));
 sky130_fd_sc_hd__o22a_1 _15100_ (.A1(net4190),
    .A2(net4184),
    .B1(net3583),
    .B2(net3581),
    .X(_07174_));
 sky130_fd_sc_hd__a21o_1 _15101_ (.A1(_07172_),
    .A2(_07173_),
    .B1(_07174_),
    .X(_07175_));
 sky130_fd_sc_hd__o21ai_1 _15102_ (.A1(_07172_),
    .A2(_07173_),
    .B1(_07175_),
    .Y(_07176_));
 sky130_fd_sc_hd__o22a_1 _15103_ (.A1(net4135),
    .A2(net4128),
    .B1(net4123),
    .B2(net4118),
    .X(_07177_));
 sky130_fd_sc_hd__o22a_1 _15104_ (.A1(net4126),
    .A2(net4124),
    .B1(net4153),
    .B2(net4148),
    .X(_07178_));
 sky130_fd_sc_hd__or2_1 _15105_ (.A(net4143),
    .B(net4140),
    .X(_07179_));
 sky130_fd_sc_hd__o211a_1 _15106_ (.A1(_07177_),
    .A2(_07178_),
    .B1(_07129_),
    .C1(net3464),
    .X(_07180_));
 sky130_fd_sc_hd__a21o_1 _15107_ (.A1(_07177_),
    .A2(_07178_),
    .B1(_07180_),
    .X(_07181_));
 sky130_fd_sc_hd__xor2_1 _15108_ (.A(_07176_),
    .B(_07181_),
    .X(_07182_));
 sky130_fd_sc_hd__xnor2_2 _15109_ (.A(net1894),
    .B(_07182_),
    .Y(_07183_));
 sky130_fd_sc_hd__xnor2_1 _15110_ (.A(_07120_),
    .B(_07115_),
    .Y(_07184_));
 sky130_fd_sc_hd__xnor2_1 _15111_ (.A(_07111_),
    .B(_07184_),
    .Y(_07185_));
 sky130_fd_sc_hd__nor2_1 _15112_ (.A(_06964_),
    .B(_07061_),
    .Y(_07186_));
 sky130_fd_sc_hd__xnor2_1 _15113_ (.A(_07116_),
    .B(_07117_),
    .Y(_07187_));
 sky130_fd_sc_hd__xnor2_1 _15114_ (.A(_07186_),
    .B(_07187_),
    .Y(_07188_));
 sky130_fd_sc_hd__nor2_1 _15115_ (.A(net4160),
    .B(net4156),
    .Y(_07189_));
 sky130_fd_sc_hd__nor2_1 _15116_ (.A(net3597),
    .B(net3591),
    .Y(_07190_));
 sky130_fd_sc_hd__nor2_1 _15117_ (.A(net3462),
    .B(net2760),
    .Y(_07191_));
 sky130_fd_sc_hd__nor2_1 _15118_ (.A(net4175),
    .B(net4173),
    .Y(_07192_));
 sky130_fd_sc_hd__nor2_1 _15119_ (.A(net3603),
    .B(_07192_),
    .Y(_07193_));
 sky130_fd_sc_hd__or2_1 _15120_ (.A(net4206),
    .B(net4203),
    .X(_07194_));
 sky130_fd_sc_hd__o22a_1 _15121_ (.A1(net4162),
    .A2(net4158),
    .B1(net4221),
    .B2(net4219),
    .X(_07195_));
 sky130_fd_sc_hd__a22o_1 _15122_ (.A1(net3503),
    .A2(net3453),
    .B1(_07064_),
    .B2(_07195_),
    .X(_07196_));
 sky130_fd_sc_hd__o21a_1 _15123_ (.A1(_07191_),
    .A2(_07193_),
    .B1(_07196_),
    .X(_07197_));
 sky130_fd_sc_hd__xnor2_1 _15124_ (.A(_07172_),
    .B(_07173_),
    .Y(_07198_));
 sky130_fd_sc_hd__xnor2_1 _15125_ (.A(_07174_),
    .B(_07198_),
    .Y(_07199_));
 sky130_fd_sc_hd__a21o_1 _15126_ (.A1(net1893),
    .A2(net1892),
    .B1(_07199_),
    .X(_07200_));
 sky130_fd_sc_hd__o21a_1 _15127_ (.A1(net1893),
    .A2(net1892),
    .B1(_07200_),
    .X(_07201_));
 sky130_fd_sc_hd__a21oi_1 _15128_ (.A1(_07183_),
    .A2(net1278),
    .B1(net1277),
    .Y(_07202_));
 sky130_fd_sc_hd__nor2_1 _15129_ (.A(_07183_),
    .B(net1278),
    .Y(_07203_));
 sky130_fd_sc_hd__clkbuf_1 _15130_ (.A(_07149_),
    .X(_07204_));
 sky130_fd_sc_hd__clkbuf_1 _15131_ (.A(net3465),
    .X(_07205_));
 sky130_fd_sc_hd__nor2_1 _15132_ (.A(net2759),
    .B(net2749),
    .Y(_07206_));
 sky130_fd_sc_hd__clkbuf_1 _15133_ (.A(net3481),
    .X(_07207_));
 sky130_fd_sc_hd__nor2_1 _15134_ (.A(net2777),
    .B(net2743),
    .Y(_07208_));
 sky130_fd_sc_hd__xnor2_1 _15135_ (.A(_07206_),
    .B(_07208_),
    .Y(_07209_));
 sky130_fd_sc_hd__o21ba_1 _15136_ (.A1(net1894),
    .A2(_07181_),
    .B1_N(_07176_),
    .X(_07210_));
 sky130_fd_sc_hd__a21o_1 _15137_ (.A1(net1894),
    .A2(_07181_),
    .B1(_07210_),
    .X(_07211_));
 sky130_fd_sc_hd__or2b_1 _15138_ (.A(net1889),
    .B_N(_07211_),
    .X(_07212_));
 sky130_fd_sc_hd__or3_1 _15139_ (.A(_07202_),
    .B(_07203_),
    .C(_07212_),
    .X(_07213_));
 sky130_fd_sc_hd__xor2_1 _15140_ (.A(net1889),
    .B(_07211_),
    .X(_07214_));
 sky130_fd_sc_hd__o21a_1 _15141_ (.A1(_07202_),
    .A2(_07203_),
    .B1(_07214_),
    .X(_07215_));
 sky130_fd_sc_hd__or3_1 _15142_ (.A(_07202_),
    .B(_07203_),
    .C(_07214_),
    .X(_07216_));
 sky130_fd_sc_hd__o211a_1 _15143_ (.A1(net991),
    .A2(_07215_),
    .B1(_07216_),
    .C1(_07212_),
    .X(_07217_));
 sky130_fd_sc_hd__o21ba_1 _15144_ (.A1(net991),
    .A2(_07213_),
    .B1_N(_07217_),
    .X(_07218_));
 sky130_fd_sc_hd__xnor2_2 _15145_ (.A(net830),
    .B(_07218_),
    .Y(_07219_));
 sky130_fd_sc_hd__nand2_1 _15146_ (.A(net2251),
    .B(net2790),
    .Y(_07220_));
 sky130_fd_sc_hd__nand2_1 _15147_ (.A(net3464),
    .B(_07129_),
    .Y(_07221_));
 sky130_fd_sc_hd__xnor2_1 _15148_ (.A(_07177_),
    .B(_07178_),
    .Y(_07222_));
 sky130_fd_sc_hd__xnor2_2 _15149_ (.A(_07221_),
    .B(_07222_),
    .Y(_07223_));
 sky130_fd_sc_hd__nor2_1 _15150_ (.A(net2757),
    .B(_07142_),
    .Y(_07224_));
 sky130_fd_sc_hd__nand2_1 _15151_ (.A(net3562),
    .B(_07224_),
    .Y(_07225_));
 sky130_fd_sc_hd__o22a_1 _15152_ (.A1(net3512),
    .A2(net3507),
    .B1(net4170),
    .B2(net4165),
    .X(_07226_));
 sky130_fd_sc_hd__o22a_1 _15153_ (.A1(net3583),
    .A2(net3581),
    .B1(net3511),
    .B2(net3506),
    .X(_07227_));
 sky130_fd_sc_hd__o22a_1 _15154_ (.A1(_07026_),
    .A2(_07028_),
    .B1(net4169),
    .B2(net4164),
    .X(_07228_));
 sky130_fd_sc_hd__xor2_2 _15155_ (.A(_07227_),
    .B(_07228_),
    .X(_07229_));
 sky130_fd_sc_hd__nor2_1 _15156_ (.A(_06992_),
    .B(net4186),
    .Y(_07230_));
 sky130_fd_sc_hd__nor2_1 _15157_ (.A(net3451),
    .B(_07125_),
    .Y(_07231_));
 sky130_fd_sc_hd__a22o_1 _15158_ (.A1(net3568),
    .A2(net2742),
    .B1(_07229_),
    .B2(net2242),
    .X(_07232_));
 sky130_fd_sc_hd__a21bo_1 _15159_ (.A1(_07223_),
    .A2(net1884),
    .B1_N(_07232_),
    .X(_07233_));
 sky130_fd_sc_hd__o21a_1 _15160_ (.A1(_07223_),
    .A2(net1884),
    .B1(_07233_),
    .X(_07234_));
 sky130_fd_sc_hd__or2_1 _15161_ (.A(net1886),
    .B(_07234_),
    .X(_07235_));
 sky130_fd_sc_hd__xnor2_1 _15162_ (.A(_07223_),
    .B(net1884),
    .Y(_07236_));
 sky130_fd_sc_hd__xnor2_2 _15163_ (.A(_07232_),
    .B(_07236_),
    .Y(_07237_));
 sky130_fd_sc_hd__xnor2_1 _15164_ (.A(_07199_),
    .B(net1892),
    .Y(_07238_));
 sky130_fd_sc_hd__xnor2_2 _15165_ (.A(net1893),
    .B(_07238_),
    .Y(_07239_));
 sky130_fd_sc_hd__clkbuf_1 _15166_ (.A(net3502),
    .X(_07240_));
 sky130_fd_sc_hd__clkbuf_1 _15167_ (.A(_07194_),
    .X(_07241_));
 sky130_fd_sc_hd__nand2_1 _15168_ (.A(net2730),
    .B(net2729),
    .Y(_07242_));
 sky130_fd_sc_hd__xnor2_1 _15169_ (.A(_07193_),
    .B(_07242_),
    .Y(_07243_));
 sky130_fd_sc_hd__xnor2_1 _15170_ (.A(_07191_),
    .B(_07243_),
    .Y(_07244_));
 sky130_fd_sc_hd__o22a_1 _15171_ (.A1(net4222),
    .A2(net4220),
    .B1(net4206),
    .B2(net4202),
    .X(_07245_));
 sky130_fd_sc_hd__o22a_1 _15172_ (.A1(net3576),
    .A2(net3572),
    .B1(net4213),
    .B2(net4211),
    .X(_07246_));
 sky130_fd_sc_hd__o22a_1 _15173_ (.A1(net4221),
    .A2(net4219),
    .B1(net4181),
    .B2(net4179),
    .X(_07247_));
 sky130_fd_sc_hd__a21o_1 _15174_ (.A1(net2849),
    .A2(net3453),
    .B1(_07247_),
    .X(_07248_));
 sky130_fd_sc_hd__a32o_1 _15175_ (.A1(net2849),
    .A2(net2730),
    .A3(net3446),
    .B1(_07246_),
    .B2(_07248_),
    .X(_07249_));
 sky130_fd_sc_hd__xor2_2 _15176_ (.A(_07229_),
    .B(net2242),
    .X(_07250_));
 sky130_fd_sc_hd__nand2_1 _15177_ (.A(net1883),
    .B(_07250_),
    .Y(_07251_));
 sky130_fd_sc_hd__nor2_1 _15178_ (.A(net1883),
    .B(_07250_),
    .Y(_07252_));
 sky130_fd_sc_hd__a21oi_2 _15179_ (.A1(net1545),
    .A2(_07251_),
    .B1(_07252_),
    .Y(_07253_));
 sky130_fd_sc_hd__a21o_1 _15180_ (.A1(_07237_),
    .A2(_07239_),
    .B1(_07253_),
    .X(_07254_));
 sky130_fd_sc_hd__o21ai_2 _15181_ (.A1(_07237_),
    .A2(_07239_),
    .B1(_07254_),
    .Y(_07255_));
 sky130_fd_sc_hd__nand2_1 _15182_ (.A(net1886),
    .B(_07234_),
    .Y(_07256_));
 sky130_fd_sc_hd__nand2_1 _15183_ (.A(_07235_),
    .B(_07256_),
    .Y(_07257_));
 sky130_fd_sc_hd__xor2_1 _15184_ (.A(net1277),
    .B(_07183_),
    .X(_07258_));
 sky130_fd_sc_hd__xnor2_2 _15185_ (.A(net1278),
    .B(_07258_),
    .Y(_07259_));
 sky130_fd_sc_hd__o21a_1 _15186_ (.A1(_07255_),
    .A2(_07257_),
    .B1(_07259_),
    .X(_07260_));
 sky130_fd_sc_hd__a21o_1 _15187_ (.A1(_07255_),
    .A2(_07257_),
    .B1(_07260_),
    .X(_07261_));
 sky130_fd_sc_hd__nor3_1 _15188_ (.A(_07259_),
    .B(_07255_),
    .C(_07235_),
    .Y(_07262_));
 sky130_fd_sc_hd__and2b_1 _15189_ (.A_N(_07215_),
    .B(_07216_),
    .X(_07263_));
 sky130_fd_sc_hd__xnor2_1 _15190_ (.A(net991),
    .B(_07263_),
    .Y(_07264_));
 sky130_fd_sc_hd__o2bb2a_1 _15191_ (.A1_N(_07235_),
    .A2_N(_07261_),
    .B1(_07262_),
    .B2(_07264_),
    .X(_07265_));
 sky130_fd_sc_hd__xnor2_1 _15192_ (.A(_07259_),
    .B(_07257_),
    .Y(_07266_));
 sky130_fd_sc_hd__xnor2_1 _15193_ (.A(_07255_),
    .B(_07266_),
    .Y(_07267_));
 sky130_fd_sc_hd__clkbuf_1 _15194_ (.A(net3554),
    .X(_07268_));
 sky130_fd_sc_hd__o211a_1 _15195_ (.A1(_07268_),
    .A2(net3486),
    .B1(_07140_),
    .C1(net2845),
    .X(_07269_));
 sky130_fd_sc_hd__o211a_1 _15196_ (.A1(net3552),
    .A2(net2757),
    .B1(net2794),
    .C1(net2819),
    .X(_07270_));
 sky130_fd_sc_hd__nor2_1 _15197_ (.A(_07269_),
    .B(_07270_),
    .Y(_07271_));
 sky130_fd_sc_hd__o22a_1 _15198_ (.A1(net3583),
    .A2(net3581),
    .B1(net4169),
    .B2(net4164),
    .X(_07272_));
 sky130_fd_sc_hd__o22a_1 _15199_ (.A1(net4190),
    .A2(net4184),
    .B1(net4121),
    .B2(net4116),
    .X(_07273_));
 sky130_fd_sc_hd__or2_1 _15200_ (.A(_07095_),
    .B(net3508),
    .X(_07274_));
 sky130_fd_sc_hd__clkbuf_1 _15201_ (.A(_07274_),
    .X(_07275_));
 sky130_fd_sc_hd__a22o_1 _15202_ (.A1(net2238),
    .A2(_07087_),
    .B1(_07272_),
    .B2(_07273_),
    .X(_07276_));
 sky130_fd_sc_hd__o21a_1 _15203_ (.A1(_07272_),
    .A2(_07273_),
    .B1(_07276_),
    .X(_07277_));
 sky130_fd_sc_hd__or2b_1 _15204_ (.A(net1882),
    .B_N(net1544),
    .X(_07278_));
 sky130_fd_sc_hd__xor2_1 _15205_ (.A(_07237_),
    .B(_07239_),
    .X(_07279_));
 sky130_fd_sc_hd__xnor2_2 _15206_ (.A(_07253_),
    .B(_07279_),
    .Y(_07280_));
 sky130_fd_sc_hd__nor2_1 _15207_ (.A(net3462),
    .B(net3529),
    .Y(_07281_));
 sky130_fd_sc_hd__xnor2_1 _15208_ (.A(_07246_),
    .B(_07247_),
    .Y(_07282_));
 sky130_fd_sc_hd__xnor2_1 _15209_ (.A(_07281_),
    .B(_07282_),
    .Y(_07283_));
 sky130_fd_sc_hd__o22a_1 _15210_ (.A1(net3586),
    .A2(net3579),
    .B1(net3594),
    .B2(net3592),
    .X(_07284_));
 sky130_fd_sc_hd__a22o_1 _15211_ (.A1(net2828),
    .A2(net3453),
    .B1(_07195_),
    .B2(_07284_),
    .X(_07285_));
 sky130_fd_sc_hd__o21a_1 _15212_ (.A1(_07195_),
    .A2(_07284_),
    .B1(_07285_),
    .X(_07286_));
 sky130_fd_sc_hd__nor2_1 _15213_ (.A(net3513),
    .B(net3505),
    .Y(_07287_));
 sky130_fd_sc_hd__nor2_1 _15214_ (.A(net2715),
    .B(_07125_),
    .Y(_07288_));
 sky130_fd_sc_hd__xnor2_1 _15215_ (.A(_07272_),
    .B(_07273_),
    .Y(_07289_));
 sky130_fd_sc_hd__xnor2_1 _15216_ (.A(_07288_),
    .B(_07289_),
    .Y(_07290_));
 sky130_fd_sc_hd__o21a_1 _15217_ (.A1(net1881),
    .A2(net1880),
    .B1(net1879),
    .X(_07291_));
 sky130_fd_sc_hd__a21o_1 _15218_ (.A1(net1881),
    .A2(net1880),
    .B1(_07291_),
    .X(_07292_));
 sky130_fd_sc_hd__xor2_1 _15219_ (.A(net1883),
    .B(_07250_),
    .X(_07293_));
 sky130_fd_sc_hd__xnor2_1 _15220_ (.A(net1545),
    .B(_07293_),
    .Y(_07294_));
 sky130_fd_sc_hd__nand2_1 _15221_ (.A(_07292_),
    .B(net1276),
    .Y(_07295_));
 sky130_fd_sc_hd__xnor2_1 _15222_ (.A(net1882),
    .B(net1544),
    .Y(_07296_));
 sky130_fd_sc_hd__o21ai_1 _15223_ (.A1(_07292_),
    .A2(net1276),
    .B1(_07296_),
    .Y(_07297_));
 sky130_fd_sc_hd__a22o_1 _15224_ (.A1(_07278_),
    .A2(_07280_),
    .B1(_07295_),
    .B2(_07297_),
    .X(_07298_));
 sky130_fd_sc_hd__o21a_1 _15225_ (.A1(_07278_),
    .A2(_07280_),
    .B1(_07298_),
    .X(_07299_));
 sky130_fd_sc_hd__xor2_1 _15226_ (.A(_07292_),
    .B(_07296_),
    .X(_07300_));
 sky130_fd_sc_hd__xnor2_1 _15227_ (.A(net1276),
    .B(_07300_),
    .Y(_07301_));
 sky130_fd_sc_hd__nor2_1 _15228_ (.A(net3451),
    .B(net3487),
    .Y(_07302_));
 sky130_fd_sc_hd__o22a_1 _15229_ (.A1(net4169),
    .A2(net4164),
    .B1(net4127),
    .B2(net4124),
    .X(_07303_));
 sky130_fd_sc_hd__or2_1 _15230_ (.A(_06992_),
    .B(net4186),
    .X(_07304_));
 sky130_fd_sc_hd__clkbuf_1 _15231_ (.A(_07304_),
    .X(_07305_));
 sky130_fd_sc_hd__o22a_1 _15232_ (.A1(net3509),
    .A2(net3504),
    .B1(net4121),
    .B2(net4116),
    .X(_07306_));
 sky130_fd_sc_hd__a31o_1 _15233_ (.A1(net2711),
    .A2(net2797),
    .A3(net3443),
    .B1(_07306_),
    .X(_07307_));
 sky130_fd_sc_hd__o21a_1 _15234_ (.A1(_07302_),
    .A2(net3443),
    .B1(_07307_),
    .X(_07308_));
 sky130_fd_sc_hd__clkbuf_1 _15235_ (.A(net3551),
    .X(_07309_));
 sky130_fd_sc_hd__nor2_1 _15236_ (.A(net2705),
    .B(net2779),
    .Y(_07310_));
 sky130_fd_sc_hd__xnor2_1 _15237_ (.A(net1881),
    .B(net1879),
    .Y(_07311_));
 sky130_fd_sc_hd__xnor2_2 _15238_ (.A(net1880),
    .B(_07311_),
    .Y(_07312_));
 sky130_fd_sc_hd__or2_1 _15239_ (.A(_07310_),
    .B(_07312_),
    .X(_07313_));
 sky130_fd_sc_hd__xnor2_1 _15240_ (.A(_07306_),
    .B(net3443),
    .Y(_07314_));
 sky130_fd_sc_hd__xnor2_2 _15241_ (.A(_07302_),
    .B(_07314_),
    .Y(_07315_));
 sky130_fd_sc_hd__nor2_1 _15242_ (.A(net3549),
    .B(net3528),
    .Y(_07316_));
 sky130_fd_sc_hd__xnor2_1 _15243_ (.A(_07195_),
    .B(_07284_),
    .Y(_07317_));
 sky130_fd_sc_hd__xnor2_2 _15244_ (.A(_07316_),
    .B(_07317_),
    .Y(_07318_));
 sky130_fd_sc_hd__o22a_1 _15245_ (.A1(net3576),
    .A2(net3572),
    .B1(net4221),
    .B2(net4219),
    .X(_07319_));
 sky130_fd_sc_hd__o22a_1 _15246_ (.A1(net3594),
    .A2(net3592),
    .B1(net4127),
    .B2(net4125),
    .X(_07320_));
 sky130_fd_sc_hd__o211a_1 _15247_ (.A1(_07319_),
    .A2(_07320_),
    .B1(net2832),
    .C1(net3453),
    .X(_07321_));
 sky130_fd_sc_hd__a21o_1 _15248_ (.A1(_07319_),
    .A2(net2704),
    .B1(_07321_),
    .X(_07322_));
 sky130_fd_sc_hd__a21o_1 _15249_ (.A1(_07315_),
    .A2(_07318_),
    .B1(_07322_),
    .X(_07323_));
 sky130_fd_sc_hd__o21a_1 _15250_ (.A1(_07315_),
    .A2(_07318_),
    .B1(_07323_),
    .X(_07324_));
 sky130_fd_sc_hd__o21a_1 _15251_ (.A1(net1878),
    .A2(_07313_),
    .B1(net1275),
    .X(_07325_));
 sky130_fd_sc_hd__a21oi_1 _15252_ (.A1(net1878),
    .A2(_07313_),
    .B1(_07325_),
    .Y(_07326_));
 sky130_fd_sc_hd__nand2_1 _15253_ (.A(net1878),
    .B(net1275),
    .Y(_07327_));
 sky130_fd_sc_hd__inv_2 _15254_ (.A(_07312_),
    .Y(_07328_));
 sky130_fd_sc_hd__a2111o_1 _15255_ (.A1(_07327_),
    .A2(net990),
    .B1(_07328_),
    .C1(net2779),
    .D1(net2705),
    .X(_07329_));
 sky130_fd_sc_hd__o21ai_1 _15256_ (.A1(net990),
    .A2(_07326_),
    .B1(_07329_),
    .Y(_07330_));
 sky130_fd_sc_hd__o21a_1 _15257_ (.A1(net1276),
    .A2(_07296_),
    .B1(_07292_),
    .X(_07331_));
 sky130_fd_sc_hd__mux2_1 _15258_ (.A0(_07331_),
    .A1(_07295_),
    .S(_07278_),
    .X(_07332_));
 sky130_fd_sc_hd__and2_1 _15259_ (.A(_07297_),
    .B(_07332_),
    .X(_07333_));
 sky130_fd_sc_hd__xnor2_1 _15260_ (.A(_07280_),
    .B(_07333_),
    .Y(_07334_));
 sky130_fd_sc_hd__a21oi_1 _15261_ (.A1(_07267_),
    .A2(_07299_),
    .B1(_07334_),
    .Y(_07335_));
 sky130_fd_sc_hd__a2bb2o_1 _15262_ (.A1_N(_07267_),
    .A2_N(_07299_),
    .B1(net829),
    .B2(_07335_),
    .X(_07336_));
 sky130_fd_sc_hd__o211a_1 _15263_ (.A1(_07259_),
    .A2(_07257_),
    .B1(_07235_),
    .C1(_07255_),
    .X(_07337_));
 sky130_fd_sc_hd__a311o_1 _15264_ (.A1(net1886),
    .A2(_07234_),
    .A3(_07259_),
    .B1(_07262_),
    .C1(_07337_),
    .X(_07338_));
 sky130_fd_sc_hd__xnor2_1 _15265_ (.A(_07264_),
    .B(_07338_),
    .Y(_07339_));
 sky130_fd_sc_hd__and2_1 _15266_ (.A(_07219_),
    .B(_07339_),
    .X(_07340_));
 sky130_fd_sc_hd__a22oi_2 _15267_ (.A1(_07219_),
    .A2(_07265_),
    .B1(_07336_),
    .B2(_07340_),
    .Y(_07341_));
 sky130_fd_sc_hd__o22ai_2 _15268_ (.A1(net991),
    .A2(_07213_),
    .B1(net830),
    .B2(_07217_),
    .Y(_07342_));
 sky130_fd_sc_hd__nand2_1 _15269_ (.A(_07008_),
    .B(net1286),
    .Y(_07343_));
 sky130_fd_sc_hd__o21bai_2 _15270_ (.A1(_07008_),
    .A2(net1286),
    .B1_N(net1287),
    .Y(_07344_));
 sky130_fd_sc_hd__nor2_1 _15271_ (.A(net2838),
    .B(net3466),
    .Y(_07345_));
 sky130_fd_sc_hd__nor2_1 _15272_ (.A(_07149_),
    .B(net2768),
    .Y(_07346_));
 sky130_fd_sc_hd__nor2_1 _15273_ (.A(net3559),
    .B(net3482),
    .Y(_07347_));
 sky130_fd_sc_hd__xnor2_1 _15274_ (.A(_07346_),
    .B(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__xnor2_1 _15275_ (.A(_07345_),
    .B(_07348_),
    .Y(_07349_));
 sky130_fd_sc_hd__o21ba_1 _15276_ (.A1(_07155_),
    .A2(_07158_),
    .B1_N(_07154_),
    .X(_07350_));
 sky130_fd_sc_hd__o21a_1 _15277_ (.A1(net6622),
    .A2(net6639),
    .B1(net7381),
    .X(_07351_));
 sky130_fd_sc_hd__o21a_1 _15278_ (.A1(net6546),
    .A2(net6594),
    .B1(\matmul0.matmul_stage_inst.e[12] ),
    .X(_07352_));
 sky130_fd_sc_hd__nor2_1 _15279_ (.A(net4095),
    .B(net4094),
    .Y(_07353_));
 sky130_fd_sc_hd__nor2_1 _15280_ (.A(net3486),
    .B(net3441),
    .Y(_07354_));
 sky130_fd_sc_hd__xor2_1 _15281_ (.A(net1877),
    .B(net2703),
    .X(_07355_));
 sky130_fd_sc_hd__xnor2_1 _15282_ (.A(net1543),
    .B(_07355_),
    .Y(_07356_));
 sky130_fd_sc_hd__or4_1 _15283_ (.A(net2839),
    .B(_07045_),
    .C(_07050_),
    .D(_07051_),
    .X(_07357_));
 sky130_fd_sc_hd__o22a_1 _15284_ (.A1(net2839),
    .A2(_07045_),
    .B1(_07050_),
    .B2(_07051_),
    .X(_07358_));
 sky130_fd_sc_hd__a21o_1 _15285_ (.A1(net1901),
    .A2(_07357_),
    .B1(_07358_),
    .X(_07359_));
 sky130_fd_sc_hd__nor2_1 _15286_ (.A(net3559),
    .B(net2768),
    .Y(_07360_));
 sky130_fd_sc_hd__nor2_1 _15287_ (.A(net2822),
    .B(net2789),
    .Y(_07361_));
 sky130_fd_sc_hd__nor2_1 _15288_ (.A(net2757),
    .B(net3483),
    .Y(_07362_));
 sky130_fd_sc_hd__o2111ai_1 _15289_ (.A1(_07360_),
    .A2(_07361_),
    .B1(net2794),
    .C1(net2790),
    .D1(_07362_),
    .Y(_07363_));
 sky130_fd_sc_hd__xnor2_1 _15290_ (.A(net1542),
    .B(net1875),
    .Y(_07364_));
 sky130_fd_sc_hd__xnor2_1 _15291_ (.A(net1274),
    .B(_07364_),
    .Y(_07365_));
 sky130_fd_sc_hd__and3_1 _15292_ (.A(_07343_),
    .B(_07344_),
    .C(_07365_),
    .X(_07366_));
 sky130_fd_sc_hd__a21oi_1 _15293_ (.A1(_07343_),
    .A2(_07344_),
    .B1(_07365_),
    .Y(_07367_));
 sky130_fd_sc_hd__buf_1 _15294_ (.A(net3602),
    .X(_07368_));
 sky130_fd_sc_hd__a22o_1 _15295_ (.A1(net6616),
    .A2(\matmul0.matmul_stage_inst.b[12] ),
    .B1(\matmul0.matmul_stage_inst.a[12] ),
    .B2(net6589),
    .X(_07369_));
 sky130_fd_sc_hd__a22o_1 _15296_ (.A1(net6631),
    .A2(\matmul0.matmul_stage_inst.d[12] ),
    .B1(\matmul0.matmul_stage_inst.c[12] ),
    .B2(net6533),
    .X(_07370_));
 sky130_fd_sc_hd__nor2_1 _15297_ (.A(net4092),
    .B(net4089),
    .Y(_07371_));
 sky130_fd_sc_hd__nor2_1 _15298_ (.A(_07368_),
    .B(net3438),
    .Y(_07372_));
 sky130_fd_sc_hd__o22a_1 _15299_ (.A1(net3596),
    .A2(net3590),
    .B1(net4198),
    .B2(net4197),
    .X(_07373_));
 sky130_fd_sc_hd__o22a_1 _15300_ (.A1(net4207),
    .A2(net4201),
    .B1(net4216),
    .B2(net4214),
    .X(_07374_));
 sky130_fd_sc_hd__xnor2_1 _15301_ (.A(_07373_),
    .B(_07374_),
    .Y(_07375_));
 sky130_fd_sc_hd__xnor2_1 _15302_ (.A(_07372_),
    .B(_07375_),
    .Y(_07376_));
 sky130_fd_sc_hd__buf_1 _15303_ (.A(net2852),
    .X(_07377_));
 sky130_fd_sc_hd__or2_1 _15304_ (.A(net4216),
    .B(net4214),
    .X(_07378_));
 sky130_fd_sc_hd__a31o_1 _15305_ (.A1(net2233),
    .A2(_07378_),
    .A3(net3598),
    .B1(_06978_),
    .X(_07379_));
 sky130_fd_sc_hd__o21a_1 _15306_ (.A1(_06968_),
    .A2(net3598),
    .B1(_07379_),
    .X(_07380_));
 sky130_fd_sc_hd__nor2_1 _15307_ (.A(net3501),
    .B(_07066_),
    .Y(_07381_));
 sky130_fd_sc_hd__o22a_1 _15308_ (.A1(net4192),
    .A2(net4186),
    .B1(net4176),
    .B2(net4174),
    .X(_07382_));
 sky130_fd_sc_hd__o22a_1 _15309_ (.A1(net3510),
    .A2(net3505),
    .B1(net4196),
    .B2(net4194),
    .X(_07383_));
 sky130_fd_sc_hd__xnor2_1 _15310_ (.A(_07382_),
    .B(_07383_),
    .Y(_07384_));
 sky130_fd_sc_hd__xnor2_1 _15311_ (.A(_07381_),
    .B(_07384_),
    .Y(_07385_));
 sky130_fd_sc_hd__xnor2_2 _15312_ (.A(net1539),
    .B(net1869),
    .Y(_07386_));
 sky130_fd_sc_hd__xnor2_4 _15313_ (.A(net1872),
    .B(_07386_),
    .Y(_07387_));
 sky130_fd_sc_hd__nor2_1 _15314_ (.A(net3545),
    .B(net3558),
    .Y(_07388_));
 sky130_fd_sc_hd__nor2_1 _15315_ (.A(net3461),
    .B(net3555),
    .Y(_07389_));
 sky130_fd_sc_hd__nor2_1 _15316_ (.A(net3495),
    .B(net3553),
    .Y(_07390_));
 sky130_fd_sc_hd__xnor2_1 _15317_ (.A(_07389_),
    .B(_07390_),
    .Y(_07391_));
 sky130_fd_sc_hd__xnor2_1 _15318_ (.A(_07388_),
    .B(_07391_),
    .Y(_07392_));
 sky130_fd_sc_hd__a21o_1 _15319_ (.A1(_06996_),
    .A2(_07001_),
    .B1(_07004_),
    .X(_07393_));
 sky130_fd_sc_hd__o21a_1 _15320_ (.A1(_06996_),
    .A2(_07001_),
    .B1(_07393_),
    .X(_07394_));
 sky130_fd_sc_hd__a22o_1 _15321_ (.A1(_07011_),
    .A2(_07015_),
    .B1(_07024_),
    .B2(_07031_),
    .X(_07395_));
 sky130_fd_sc_hd__o21a_1 _15322_ (.A1(_07024_),
    .A2(_07031_),
    .B1(_07395_),
    .X(_07396_));
 sky130_fd_sc_hd__xnor2_1 _15323_ (.A(net2229),
    .B(net1866),
    .Y(_07397_));
 sky130_fd_sc_hd__xnor2_2 _15324_ (.A(net1868),
    .B(_07397_),
    .Y(_07398_));
 sky130_fd_sc_hd__o21a_1 _15325_ (.A1(net2256),
    .A2(net2252),
    .B1(net1902),
    .X(_07399_));
 sky130_fd_sc_hd__a21o_1 _15326_ (.A1(net2256),
    .A2(net2252),
    .B1(_07399_),
    .X(_07400_));
 sky130_fd_sc_hd__xor2_2 _15327_ (.A(_07398_),
    .B(_07400_),
    .X(_07401_));
 sky130_fd_sc_hd__xnor2_4 _15328_ (.A(_07387_),
    .B(_07401_),
    .Y(_07402_));
 sky130_fd_sc_hd__o21ai_1 _15329_ (.A1(_07366_),
    .A2(_07367_),
    .B1(_07402_),
    .Y(_07403_));
 sky130_fd_sc_hd__or3_1 _15330_ (.A(_07402_),
    .B(_07366_),
    .C(_07367_),
    .X(_07404_));
 sky130_fd_sc_hd__and2_1 _15331_ (.A(_07403_),
    .B(_07404_),
    .X(_07405_));
 sky130_fd_sc_hd__or2_1 _15332_ (.A(_07124_),
    .B(net1117),
    .X(_07406_));
 sky130_fd_sc_hd__and2_1 _15333_ (.A(_07124_),
    .B(net1117),
    .X(_07407_));
 sky130_fd_sc_hd__a21o_1 _15334_ (.A1(net1280),
    .A2(_07406_),
    .B1(_07407_),
    .X(_07408_));
 sky130_fd_sc_hd__nand3_1 _15335_ (.A(_07073_),
    .B(net1280),
    .C(_07407_),
    .Y(_07409_));
 sky130_fd_sc_hd__o221ai_2 _15336_ (.A1(net1280),
    .A2(_07406_),
    .B1(_07408_),
    .B2(_07073_),
    .C1(_07409_),
    .Y(_07410_));
 sky130_fd_sc_hd__xnor2_1 _15337_ (.A(_07405_),
    .B(_07410_),
    .Y(_07411_));
 sky130_fd_sc_hd__nand2_1 _15338_ (.A(net2740),
    .B(_07224_),
    .Y(_07412_));
 sky130_fd_sc_hd__xor2_1 _15339_ (.A(net1878),
    .B(net1275),
    .X(_07413_));
 sky130_fd_sc_hd__xnor2_1 _15340_ (.A(_07310_),
    .B(_07312_),
    .Y(_07414_));
 sky130_fd_sc_hd__xnor2_1 _15341_ (.A(_07413_),
    .B(_07414_),
    .Y(_07415_));
 sky130_fd_sc_hd__a211o_1 _15342_ (.A1(net2236),
    .A2(net2796),
    .B1(net2756),
    .C1(net3497),
    .X(_07416_));
 sky130_fd_sc_hd__a211o_1 _15343_ (.A1(net2811),
    .A2(net2782),
    .B1(net3487),
    .C1(net2716),
    .X(_07417_));
 sky130_fd_sc_hd__nand2_1 _15344_ (.A(_07416_),
    .B(_07417_),
    .Y(_07418_));
 sky130_fd_sc_hd__nor2_1 _15345_ (.A(net2760),
    .B(net2756),
    .Y(_07419_));
 sky130_fd_sc_hd__nor2_1 _15346_ (.A(net3528),
    .B(net2801),
    .Y(_07420_));
 sky130_fd_sc_hd__nor2_1 _15347_ (.A(net2835),
    .B(net2702),
    .Y(_07421_));
 sky130_fd_sc_hd__and3_1 _15348_ (.A(net2726),
    .B(net2782),
    .C(net2704),
    .X(_07422_));
 sky130_fd_sc_hd__o22a_1 _15349_ (.A1(_07419_),
    .A2(_07420_),
    .B1(_07421_),
    .B2(_07422_),
    .X(_07423_));
 sky130_fd_sc_hd__nand2_1 _15350_ (.A(net2832),
    .B(net2726),
    .Y(_07424_));
 sky130_fd_sc_hd__xnor2_1 _15351_ (.A(_07319_),
    .B(net2704),
    .Y(_07425_));
 sky130_fd_sc_hd__xnor2_1 _15352_ (.A(_07424_),
    .B(_07425_),
    .Y(_07426_));
 sky130_fd_sc_hd__o21ba_1 _15353_ (.A1(_07418_),
    .A2(_07423_),
    .B1_N(_07426_),
    .X(_07427_));
 sky130_fd_sc_hd__a21o_1 _15354_ (.A1(_07418_),
    .A2(_07423_),
    .B1(_07427_),
    .X(_07428_));
 sky130_fd_sc_hd__xnor2_1 _15355_ (.A(_07315_),
    .B(_07322_),
    .Y(_07429_));
 sky130_fd_sc_hd__xnor2_1 _15356_ (.A(_07318_),
    .B(_07429_),
    .Y(_07430_));
 sky130_fd_sc_hd__nand2_1 _15357_ (.A(net1116),
    .B(_07430_),
    .Y(_07431_));
 sky130_fd_sc_hd__or2_1 _15358_ (.A(net1116),
    .B(_07430_),
    .X(_07432_));
 sky130_fd_sc_hd__nand4_1 _15359_ (.A(_07412_),
    .B(_07415_),
    .C(_07431_),
    .D(_07432_),
    .Y(_07433_));
 sky130_fd_sc_hd__or3b_1 _15360_ (.A(_07412_),
    .B(_07432_),
    .C_N(_07415_),
    .X(_07434_));
 sky130_fd_sc_hd__o311a_1 _15361_ (.A1(_07412_),
    .A2(_07415_),
    .A3(_07431_),
    .B1(_07433_),
    .C1(_07434_),
    .X(_07435_));
 sky130_fd_sc_hd__xor2_1 _15362_ (.A(_07418_),
    .B(_07423_),
    .X(_07436_));
 sky130_fd_sc_hd__xnor2_1 _15363_ (.A(_07426_),
    .B(_07436_),
    .Y(_07437_));
 sky130_fd_sc_hd__or2_1 _15364_ (.A(net3596),
    .B(net3590),
    .X(_07438_));
 sky130_fd_sc_hd__a22o_1 _15365_ (.A1(net2233),
    .A2(net2824),
    .B1(net2249),
    .B2(_07438_),
    .X(_07439_));
 sky130_fd_sc_hd__and3_1 _15366_ (.A(net2233),
    .B(net2249),
    .C(net2704),
    .X(_07440_));
 sky130_fd_sc_hd__a31o_1 _15367_ (.A1(net2726),
    .A2(net2782),
    .A3(_07439_),
    .B1(_07440_),
    .X(_07441_));
 sky130_fd_sc_hd__xnor2_1 _15368_ (.A(_07420_),
    .B(_07421_),
    .Y(_07442_));
 sky130_fd_sc_hd__xnor2_1 _15369_ (.A(_07419_),
    .B(_07442_),
    .Y(_07443_));
 sky130_fd_sc_hd__nor2_1 _15370_ (.A(_07438_),
    .B(net2824),
    .Y(_07444_));
 sky130_fd_sc_hd__o211a_1 _15371_ (.A1(net2704),
    .A2(_07444_),
    .B1(_07224_),
    .C1(net3445),
    .X(_07445_));
 sky130_fd_sc_hd__or2_1 _15372_ (.A(_07443_),
    .B(_07445_),
    .X(_07446_));
 sky130_fd_sc_hd__and2_1 _15373_ (.A(_07443_),
    .B(_07445_),
    .X(_07447_));
 sky130_fd_sc_hd__a21o_1 _15374_ (.A1(_07441_),
    .A2(_07446_),
    .B1(_07447_),
    .X(_07448_));
 sky130_fd_sc_hd__or2_1 _15375_ (.A(_07437_),
    .B(_07447_),
    .X(_07449_));
 sky130_fd_sc_hd__a22o_1 _15376_ (.A1(_07437_),
    .A2(_07446_),
    .B1(_07449_),
    .B2(_07441_),
    .X(_07450_));
 sky130_fd_sc_hd__and3_1 _15377_ (.A(net2811),
    .B(net2249),
    .C(_07450_),
    .X(_07451_));
 sky130_fd_sc_hd__a21oi_1 _15378_ (.A1(_07437_),
    .A2(_07448_),
    .B1(_07451_),
    .Y(_07452_));
 sky130_fd_sc_hd__or2_1 _15379_ (.A(net1878),
    .B(net1275),
    .X(_07453_));
 sky130_fd_sc_hd__nand2_1 _15380_ (.A(_07310_),
    .B(_07312_),
    .Y(_07454_));
 sky130_fd_sc_hd__mux2_1 _15381_ (.A0(_07327_),
    .A1(_07453_),
    .S(_07454_),
    .X(_07455_));
 sky130_fd_sc_hd__a21o_1 _15382_ (.A1(net1878),
    .A2(net1275),
    .B1(_07313_),
    .X(_07456_));
 sky130_fd_sc_hd__nand2_1 _15383_ (.A(_07455_),
    .B(_07456_),
    .Y(_07457_));
 sky130_fd_sc_hd__xnor2_1 _15384_ (.A(net990),
    .B(_07457_),
    .Y(_07458_));
 sky130_fd_sc_hd__and3_1 _15385_ (.A(_07140_),
    .B(net2251),
    .C(net2740),
    .X(_07459_));
 sky130_fd_sc_hd__a21o_1 _15386_ (.A1(_07459_),
    .A2(net1116),
    .B1(_07430_),
    .X(_07460_));
 sky130_fd_sc_hd__o21ai_1 _15387_ (.A1(_07459_),
    .A2(net1116),
    .B1(_07460_),
    .Y(_07461_));
 sky130_fd_sc_hd__nand2_1 _15388_ (.A(_07327_),
    .B(_07453_),
    .Y(_07462_));
 sky130_fd_sc_hd__mux2_1 _15389_ (.A0(_07313_),
    .A1(_07454_),
    .S(net990),
    .X(_07463_));
 sky130_fd_sc_hd__mux2_1 _15390_ (.A0(_07453_),
    .A1(_07327_),
    .S(net990),
    .X(_07464_));
 sky130_fd_sc_hd__o22a_1 _15391_ (.A1(_07462_),
    .A2(_07463_),
    .B1(_07414_),
    .B2(_07464_),
    .X(_07465_));
 sky130_fd_sc_hd__o32ai_1 _15392_ (.A1(_07435_),
    .A2(net779),
    .A3(_07458_),
    .B1(_07461_),
    .B2(_07465_),
    .Y(_07466_));
 sky130_fd_sc_hd__xor2_1 _15393_ (.A(_07267_),
    .B(_07299_),
    .X(_07467_));
 sky130_fd_sc_hd__xnor2_1 _15394_ (.A(net829),
    .B(_07334_),
    .Y(_07468_));
 sky130_fd_sc_hd__and4_1 _15395_ (.A(_07339_),
    .B(net725),
    .C(_07467_),
    .D(_07468_),
    .X(_07469_));
 sky130_fd_sc_hd__xor2_1 _15396_ (.A(_07219_),
    .B(_07265_),
    .X(_07470_));
 sky130_fd_sc_hd__a22oi_2 _15397_ (.A1(_07342_),
    .A2(_07411_),
    .B1(_07469_),
    .B2(_07470_),
    .Y(_07471_));
 sky130_fd_sc_hd__nor2_1 _15398_ (.A(_07342_),
    .B(_07411_),
    .Y(_07472_));
 sky130_fd_sc_hd__a21o_1 _15399_ (.A1(_07403_),
    .A2(_07404_),
    .B1(_07407_),
    .X(_07473_));
 sky130_fd_sc_hd__a22oi_1 _15400_ (.A1(_07405_),
    .A2(_07406_),
    .B1(_07473_),
    .B2(net1280),
    .Y(_07474_));
 sky130_fd_sc_hd__o2bb2a_1 _15401_ (.A1_N(_07405_),
    .A2_N(_07408_),
    .B1(_07474_),
    .B2(_07072_),
    .X(_07475_));
 sky130_fd_sc_hd__nor2_1 _15402_ (.A(net2838),
    .B(net2768),
    .Y(_07476_));
 sky130_fd_sc_hd__and2_1 _15403_ (.A(_07206_),
    .B(_07476_),
    .X(_07477_));
 sky130_fd_sc_hd__o22a_2 _15404_ (.A1(_07345_),
    .A2(_07346_),
    .B1(_07347_),
    .B2(_07477_),
    .X(_07478_));
 sky130_fd_sc_hd__o22a_1 _15405_ (.A1(net3584),
    .A2(net3577),
    .B1(net4098),
    .B2(net4096),
    .X(_07479_));
 sky130_fd_sc_hd__o22a_1 _15406_ (.A1(net3573),
    .A2(net3569),
    .B1(net4105),
    .B2(net4101),
    .X(_07480_));
 sky130_fd_sc_hd__xor2_1 _15407_ (.A(_07479_),
    .B(_07480_),
    .X(_07481_));
 sky130_fd_sc_hd__xnor2_1 _15408_ (.A(_07360_),
    .B(_07481_),
    .Y(_07482_));
 sky130_fd_sc_hd__o21a_1 _15409_ (.A1(net6621),
    .A2(net6640),
    .B1(\matmul0.matmul_stage_inst.f[13] ),
    .X(_07483_));
 sky130_fd_sc_hd__o21a_1 _15410_ (.A1(net6541),
    .A2(net6594),
    .B1(\matmul0.matmul_stage_inst.e[13] ),
    .X(_07484_));
 sky130_fd_sc_hd__nor2_1 _15411_ (.A(net4087),
    .B(net4086),
    .Y(_07485_));
 sky130_fd_sc_hd__or2_1 _15412_ (.A(net4095),
    .B(net4094),
    .X(_07486_));
 sky130_fd_sc_hd__o211a_1 _15413_ (.A1(net2778),
    .A2(net3428),
    .B1(net3426),
    .C1(net2781),
    .X(_07487_));
 sky130_fd_sc_hd__or2_1 _15414_ (.A(net4087),
    .B(net4086),
    .X(_07488_));
 sky130_fd_sc_hd__clkbuf_1 _15415_ (.A(_07488_),
    .X(_07489_));
 sky130_fd_sc_hd__o211a_1 _15416_ (.A1(net2755),
    .A2(net3441),
    .B1(net2696),
    .C1(net2795),
    .X(_07490_));
 sky130_fd_sc_hd__nor2_1 _15417_ (.A(_07487_),
    .B(_07490_),
    .Y(_07491_));
 sky130_fd_sc_hd__nand2_1 _15418_ (.A(net1865),
    .B(net1864),
    .Y(_07492_));
 sky130_fd_sc_hd__inv_2 _15419_ (.A(_07492_),
    .Y(_07493_));
 sky130_fd_sc_hd__nor2_1 _15420_ (.A(net1865),
    .B(net1864),
    .Y(_07494_));
 sky130_fd_sc_hd__nor2_1 _15421_ (.A(_07493_),
    .B(_07494_),
    .Y(_07495_));
 sky130_fd_sc_hd__xor2_2 _15422_ (.A(_07478_),
    .B(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__o21a_1 _15423_ (.A1(net2229),
    .A2(net1866),
    .B1(net1868),
    .X(_07497_));
 sky130_fd_sc_hd__a21o_1 _15424_ (.A1(net2229),
    .A2(net1866),
    .B1(_07497_),
    .X(_07498_));
 sky130_fd_sc_hd__o21a_1 _15425_ (.A1(net1543),
    .A2(net2703),
    .B1(net1877),
    .X(_07499_));
 sky130_fd_sc_hd__a21oi_1 _15426_ (.A1(net1543),
    .A2(net2703),
    .B1(_07499_),
    .Y(_07500_));
 sky130_fd_sc_hd__xnor2_1 _15427_ (.A(net1273),
    .B(_07500_),
    .Y(_07501_));
 sky130_fd_sc_hd__xnor2_2 _15428_ (.A(_07496_),
    .B(_07501_),
    .Y(_07502_));
 sky130_fd_sc_hd__o21a_1 _15429_ (.A1(_07398_),
    .A2(_07400_),
    .B1(_07387_),
    .X(_07503_));
 sky130_fd_sc_hd__a21o_1 _15430_ (.A1(_07398_),
    .A2(_07400_),
    .B1(_07503_),
    .X(_07504_));
 sky130_fd_sc_hd__buf_1 _15431_ (.A(net3534),
    .X(_07505_));
 sky130_fd_sc_hd__nor2_1 _15432_ (.A(net3450),
    .B(net2690),
    .Y(_07506_));
 sky130_fd_sc_hd__o22a_1 _15433_ (.A1(net4172),
    .A2(net4166),
    .B1(net4199),
    .B2(_06977_),
    .X(_07507_));
 sky130_fd_sc_hd__o22a_1 _15434_ (.A1(net3510),
    .A2(net3505),
    .B1(net4210),
    .B2(net4208),
    .X(_07508_));
 sky130_fd_sc_hd__xnor2_1 _15435_ (.A(net3423),
    .B(net2689),
    .Y(_07509_));
 sky130_fd_sc_hd__xnor2_1 _15436_ (.A(_07506_),
    .B(_07509_),
    .Y(_07510_));
 sky130_fd_sc_hd__or2_1 _15437_ (.A(net4092),
    .B(net4089),
    .X(_07511_));
 sky130_fd_sc_hd__a31o_1 _15438_ (.A1(_07377_),
    .A2(_07511_),
    .A3(_07373_),
    .B1(_07374_),
    .X(_07512_));
 sky130_fd_sc_hd__o21a_1 _15439_ (.A1(_07372_),
    .A2(_07373_),
    .B1(_07512_),
    .X(_07513_));
 sky130_fd_sc_hd__a22o_1 _15440_ (.A1(net6631),
    .A2(\matmul0.matmul_stage_inst.d[13] ),
    .B1(\matmul0.matmul_stage_inst.c[13] ),
    .B2(net6533),
    .X(_07514_));
 sky130_fd_sc_hd__a22o_1 _15441_ (.A1(net6616),
    .A2(\matmul0.matmul_stage_inst.b[13] ),
    .B1(\matmul0.matmul_stage_inst.a[13] ),
    .B2(net6581),
    .X(_07515_));
 sky130_fd_sc_hd__nor2_1 _15442_ (.A(net4083),
    .B(net4081),
    .Y(_07516_));
 sky130_fd_sc_hd__nor2_1 _15443_ (.A(net3602),
    .B(net3419),
    .Y(_07517_));
 sky130_fd_sc_hd__o22a_1 _15444_ (.A1(net3597),
    .A2(net3591),
    .B1(net4216),
    .B2(net4214),
    .X(_07518_));
 sky130_fd_sc_hd__o22a_1 _15445_ (.A1(_06974_),
    .A2(net4201),
    .B1(net4092),
    .B2(net4089),
    .X(_07519_));
 sky130_fd_sc_hd__xnor2_1 _15446_ (.A(_07518_),
    .B(_07519_),
    .Y(_07520_));
 sky130_fd_sc_hd__xnor2_2 _15447_ (.A(_07517_),
    .B(_07520_),
    .Y(_07521_));
 sky130_fd_sc_hd__xnor2_1 _15448_ (.A(_07513_),
    .B(_07521_),
    .Y(_07522_));
 sky130_fd_sc_hd__xnor2_1 _15449_ (.A(_07510_),
    .B(_07522_),
    .Y(_07523_));
 sky130_fd_sc_hd__a21o_1 _15450_ (.A1(net1539),
    .A2(net1869),
    .B1(net1872),
    .X(_07524_));
 sky130_fd_sc_hd__o21a_1 _15451_ (.A1(net1539),
    .A2(net1869),
    .B1(_07524_),
    .X(_07525_));
 sky130_fd_sc_hd__o22a_1 _15452_ (.A1(net4161),
    .A2(net4157),
    .B1(net4143),
    .B2(net4140),
    .X(_07526_));
 sky130_fd_sc_hd__nor2_1 _15453_ (.A(net2807),
    .B(net3555),
    .Y(_07527_));
 sky130_fd_sc_hd__or2_1 _15454_ (.A(net4175),
    .B(net4173),
    .X(_07528_));
 sky130_fd_sc_hd__nand2_1 _15455_ (.A(net3412),
    .B(_07016_),
    .Y(_07529_));
 sky130_fd_sc_hd__xnor2_1 _15456_ (.A(_07527_),
    .B(_07529_),
    .Y(_07530_));
 sky130_fd_sc_hd__xnor2_1 _15457_ (.A(_07526_),
    .B(_07530_),
    .Y(_07531_));
 sky130_fd_sc_hd__a31o_1 _15458_ (.A1(net2814),
    .A2(_07063_),
    .A3(_07382_),
    .B1(_07383_),
    .X(_07532_));
 sky130_fd_sc_hd__o21a_1 _15459_ (.A1(_07381_),
    .A2(_07382_),
    .B1(_07532_),
    .X(_07533_));
 sky130_fd_sc_hd__clkbuf_1 _15460_ (.A(_07179_),
    .X(_07534_));
 sky130_fd_sc_hd__a22o_1 _15461_ (.A1(net2848),
    .A2(net2820),
    .B1(net2686),
    .B2(net2827),
    .X(_07535_));
 sky130_fd_sc_hd__and4_1 _15462_ (.A(net2827),
    .B(_07012_),
    .C(net2820),
    .D(net2686),
    .X(_07536_));
 sky130_fd_sc_hd__a21o_1 _15463_ (.A1(_07390_),
    .A2(_07535_),
    .B1(_07536_),
    .X(_07537_));
 sky130_fd_sc_hd__xor2_1 _15464_ (.A(net1861),
    .B(net1860),
    .X(_07538_));
 sky130_fd_sc_hd__xnor2_2 _15465_ (.A(net1538),
    .B(_07538_),
    .Y(_07539_));
 sky130_fd_sc_hd__xor2_1 _15466_ (.A(_07525_),
    .B(_07539_),
    .X(_07540_));
 sky130_fd_sc_hd__xnor2_2 _15467_ (.A(net1113),
    .B(_07540_),
    .Y(_07541_));
 sky130_fd_sc_hd__xor2_1 _15468_ (.A(_07504_),
    .B(_07541_),
    .X(_07542_));
 sky130_fd_sc_hd__xnor2_2 _15469_ (.A(_07502_),
    .B(_07542_),
    .Y(_07543_));
 sky130_fd_sc_hd__and3_1 _15470_ (.A(_07343_),
    .B(_07344_),
    .C(net1542),
    .X(_07544_));
 sky130_fd_sc_hd__and2_1 _15471_ (.A(net1875),
    .B(_07544_),
    .X(_07545_));
 sky130_fd_sc_hd__a21o_1 _15472_ (.A1(_07343_),
    .A2(_07344_),
    .B1(net1542),
    .X(_07546_));
 sky130_fd_sc_hd__o211a_1 _15473_ (.A1(net1875),
    .A2(_07544_),
    .B1(_07546_),
    .C1(net1274),
    .X(_07547_));
 sky130_fd_sc_hd__o21ai_1 _15474_ (.A1(_07545_),
    .A2(_07547_),
    .B1(_07402_),
    .Y(_07548_));
 sky130_fd_sc_hd__nand2_1 _15475_ (.A(net1274),
    .B(_07545_),
    .Y(_07549_));
 sky130_fd_sc_hd__o21a_1 _15476_ (.A1(net1875),
    .A2(_07544_),
    .B1(_07546_),
    .X(_07550_));
 sky130_fd_sc_hd__a211o_1 _15477_ (.A1(_07402_),
    .A2(net1274),
    .B1(net1875),
    .C1(_07546_),
    .X(_07551_));
 sky130_fd_sc_hd__o31a_1 _15478_ (.A1(_07402_),
    .A2(net1274),
    .A3(_07550_),
    .B1(_07551_),
    .X(_07552_));
 sky130_fd_sc_hd__nand3_1 _15479_ (.A(_07548_),
    .B(_07549_),
    .C(_07552_),
    .Y(_07553_));
 sky130_fd_sc_hd__xor2_1 _15480_ (.A(_07543_),
    .B(_07553_),
    .X(_07554_));
 sky130_fd_sc_hd__xor2_1 _15481_ (.A(_07475_),
    .B(_07554_),
    .X(_07555_));
 sky130_fd_sc_hd__a211o_1 _15482_ (.A1(_07341_),
    .A2(_07471_),
    .B1(_07472_),
    .C1(net675),
    .X(_07556_));
 sky130_fd_sc_hd__a21o_1 _15483_ (.A1(_07341_),
    .A2(_07471_),
    .B1(_07472_),
    .X(_07557_));
 sky130_fd_sc_hd__nand2_1 _15484_ (.A(_07557_),
    .B(net675),
    .Y(_07558_));
 sky130_fd_sc_hd__and2_1 _15485_ (.A(_07556_),
    .B(_07558_),
    .X(_07559_));
 sky130_fd_sc_hd__buf_1 _15486_ (.A(net3478),
    .X(_07560_));
 sky130_fd_sc_hd__mux2_1 _15487_ (.A0(\matmul0.matmul_stage_inst.mult1[0] ),
    .A1(net494),
    .S(net2678),
    .X(_07561_));
 sky130_fd_sc_hd__clkbuf_1 _15488_ (.A(_07561_),
    .X(_00215_));
 sky130_fd_sc_hd__and2b_1 _15489_ (.A_N(_07475_),
    .B(_07554_),
    .X(_07562_));
 sky130_fd_sc_hd__or2_1 _15490_ (.A(net1274),
    .B(net1875),
    .X(_07563_));
 sky130_fd_sc_hd__or2_1 _15491_ (.A(_07402_),
    .B(_07544_),
    .X(_07564_));
 sky130_fd_sc_hd__a22o_1 _15492_ (.A1(_07543_),
    .A2(_07563_),
    .B1(_07564_),
    .B2(_07546_),
    .X(_07565_));
 sky130_fd_sc_hd__a21o_1 _15493_ (.A1(_07543_),
    .A2(_07546_),
    .B1(_07402_),
    .X(_07566_));
 sky130_fd_sc_hd__or2_1 _15494_ (.A(_07543_),
    .B(_07544_),
    .X(_07567_));
 sky130_fd_sc_hd__a22o_1 _15495_ (.A1(net1274),
    .A2(net1875),
    .B1(_07566_),
    .B2(_07567_),
    .X(_07568_));
 sky130_fd_sc_hd__o211ai_2 _15496_ (.A1(_07543_),
    .A2(_07563_),
    .B1(_07565_),
    .C1(_07568_),
    .Y(_07569_));
 sky130_fd_sc_hd__nor2_1 _15497_ (.A(net2800),
    .B(net3440),
    .Y(_07570_));
 sky130_fd_sc_hd__o22a_1 _15498_ (.A1(net4119),
    .A2(net4114),
    .B1(net4087),
    .B2(net4086),
    .X(_07571_));
 sky130_fd_sc_hd__o21a_1 _15499_ (.A1(net6622),
    .A2(net6643),
    .B1(net7380),
    .X(_07572_));
 sky130_fd_sc_hd__o21a_1 _15500_ (.A1(net6540),
    .A2(net6594),
    .B1(\matmul0.matmul_stage_inst.e[14] ),
    .X(_07573_));
 sky130_fd_sc_hd__o22a_1 _15501_ (.A1(net4111),
    .A2(net4108),
    .B1(net4079),
    .B2(net4077),
    .X(_07574_));
 sky130_fd_sc_hd__xnor2_1 _15502_ (.A(net3407),
    .B(net3404),
    .Y(_07575_));
 sky130_fd_sc_hd__xnor2_2 _15503_ (.A(net2228),
    .B(_07575_),
    .Y(_07576_));
 sky130_fd_sc_hd__or2_1 _15504_ (.A(_07479_),
    .B(_07480_),
    .X(_07577_));
 sky130_fd_sc_hd__a32o_1 _15505_ (.A1(_07133_),
    .A2(_07146_),
    .A3(net3566),
    .B1(_07360_),
    .B2(_07577_),
    .X(_07578_));
 sky130_fd_sc_hd__o22a_1 _15506_ (.A1(net3573),
    .A2(net3569),
    .B1(net4098),
    .B2(net4096),
    .X(_07579_));
 sky130_fd_sc_hd__o22a_1 _15507_ (.A1(net4160),
    .A2(net4156),
    .B1(net4105),
    .B2(net4101),
    .X(_07580_));
 sky130_fd_sc_hd__xnor2_1 _15508_ (.A(net2677),
    .B(_07580_),
    .Y(_07581_));
 sky130_fd_sc_hd__xnor2_2 _15509_ (.A(_07476_),
    .B(_07581_),
    .Y(_07582_));
 sky130_fd_sc_hd__xor2_1 _15510_ (.A(net1859),
    .B(_07582_),
    .X(_07583_));
 sky130_fd_sc_hd__xnor2_2 _15511_ (.A(_07576_),
    .B(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__nand2_1 _15512_ (.A(net1861),
    .B(net1860),
    .Y(_07585_));
 sky130_fd_sc_hd__nor2_1 _15513_ (.A(net1861),
    .B(net1860),
    .Y(_07586_));
 sky130_fd_sc_hd__a21oi_1 _15514_ (.A1(net1538),
    .A2(_07585_),
    .B1(_07586_),
    .Y(_07587_));
 sky130_fd_sc_hd__o21ai_2 _15515_ (.A1(_07478_),
    .A2(_07494_),
    .B1(_07492_),
    .Y(_07588_));
 sky130_fd_sc_hd__xnor2_1 _15516_ (.A(net1272),
    .B(_07588_),
    .Y(_07589_));
 sky130_fd_sc_hd__xnor2_2 _15517_ (.A(_07584_),
    .B(_07589_),
    .Y(_07590_));
 sky130_fd_sc_hd__a21o_1 _15518_ (.A1(_07525_),
    .A2(_07539_),
    .B1(net1113),
    .X(_07591_));
 sky130_fd_sc_hd__o21a_1 _15519_ (.A1(_07525_),
    .A2(_07539_),
    .B1(_07591_),
    .X(_07592_));
 sky130_fd_sc_hd__nor2_1 _15520_ (.A(net3497),
    .B(net3600),
    .Y(_07593_));
 sky130_fd_sc_hd__nor2_1 _15521_ (.A(net3447),
    .B(net3518),
    .Y(_07594_));
 sky130_fd_sc_hd__nor2_1 _15522_ (.A(net2717),
    .B(net3537),
    .Y(_07595_));
 sky130_fd_sc_hd__xnor2_1 _15523_ (.A(_07594_),
    .B(_07595_),
    .Y(_07596_));
 sky130_fd_sc_hd__xnor2_1 _15524_ (.A(_07593_),
    .B(_07596_),
    .Y(_07597_));
 sky130_fd_sc_hd__or2_1 _15525_ (.A(net4083),
    .B(net4081),
    .X(_07598_));
 sky130_fd_sc_hd__a31o_1 _15526_ (.A1(net2852),
    .A2(_07598_),
    .A3(_07518_),
    .B1(_07519_),
    .X(_07599_));
 sky130_fd_sc_hd__o21a_1 _15527_ (.A1(_07517_),
    .A2(_07518_),
    .B1(_07599_),
    .X(_07600_));
 sky130_fd_sc_hd__o21a_1 _15528_ (.A1(net6642),
    .A2(net6593),
    .B1(net7401),
    .X(_07601_));
 sky130_fd_sc_hd__a22o_1 _15529_ (.A1(net6542),
    .A2(\matmul0.matmul_stage_inst.c[14] ),
    .B1(\matmul0.matmul_stage_inst.b[14] ),
    .B2(net6614),
    .X(_07602_));
 sky130_fd_sc_hd__nor2_1 _15530_ (.A(net4075),
    .B(net4074),
    .Y(_07603_));
 sky130_fd_sc_hd__nor2_1 _15531_ (.A(net2701),
    .B(net3399),
    .Y(_07604_));
 sky130_fd_sc_hd__o22a_1 _15532_ (.A1(net3597),
    .A2(net3591),
    .B1(net4092),
    .B2(net4089),
    .X(_07605_));
 sky130_fd_sc_hd__o22a_1 _15533_ (.A1(net4207),
    .A2(net4201),
    .B1(net4083),
    .B2(net4081),
    .X(_07606_));
 sky130_fd_sc_hd__xnor2_1 _15534_ (.A(_07605_),
    .B(_07606_),
    .Y(_07607_));
 sky130_fd_sc_hd__xnor2_1 _15535_ (.A(_07604_),
    .B(net2227),
    .Y(_07608_));
 sky130_fd_sc_hd__xnor2_1 _15536_ (.A(net1857),
    .B(_07608_),
    .Y(_07609_));
 sky130_fd_sc_hd__xnor2_1 _15537_ (.A(_07597_),
    .B(_07609_),
    .Y(_07610_));
 sky130_fd_sc_hd__a21o_1 _15538_ (.A1(_07513_),
    .A2(_07521_),
    .B1(_07510_),
    .X(_07611_));
 sky130_fd_sc_hd__o21a_1 _15539_ (.A1(_07513_),
    .A2(_07521_),
    .B1(_07611_),
    .X(_07612_));
 sky130_fd_sc_hd__nor2_2 _15540_ (.A(net2806),
    .B(net3557),
    .Y(_07613_));
 sky130_fd_sc_hd__nor2_1 _15541_ (.A(net3532),
    .B(net3552),
    .Y(_07614_));
 sky130_fd_sc_hd__nor2_1 _15542_ (.A(net3456),
    .B(net3554),
    .Y(_07615_));
 sky130_fd_sc_hd__xor2_1 _15543_ (.A(_07614_),
    .B(_07615_),
    .X(_07616_));
 sky130_fd_sc_hd__xnor2_2 _15544_ (.A(_07613_),
    .B(_07616_),
    .Y(_07617_));
 sky130_fd_sc_hd__a22o_1 _15545_ (.A1(net2713),
    .A2(net3494),
    .B1(net3423),
    .B2(net2689),
    .X(_07618_));
 sky130_fd_sc_hd__o21a_1 _15546_ (.A1(net3423),
    .A2(net2689),
    .B1(_07618_),
    .X(_07619_));
 sky130_fd_sc_hd__a32o_1 _15547_ (.A1(net3502),
    .A2(net2820),
    .A3(_07526_),
    .B1(_07016_),
    .B2(net3412),
    .X(_07620_));
 sky130_fd_sc_hd__o21a_1 _15548_ (.A1(_07526_),
    .A2(_07527_),
    .B1(_07620_),
    .X(_07621_));
 sky130_fd_sc_hd__xor2_1 _15549_ (.A(net1854),
    .B(net1853),
    .X(_07622_));
 sky130_fd_sc_hd__xnor2_2 _15550_ (.A(_07617_),
    .B(_07622_),
    .Y(_07623_));
 sky130_fd_sc_hd__xnor2_1 _15551_ (.A(net1109),
    .B(_07623_),
    .Y(_07624_));
 sky130_fd_sc_hd__xnor2_2 _15552_ (.A(net1270),
    .B(_07624_),
    .Y(_07625_));
 sky130_fd_sc_hd__xnor2_1 _15553_ (.A(net889),
    .B(_07625_),
    .Y(_07626_));
 sky130_fd_sc_hd__xnor2_2 _15554_ (.A(_07590_),
    .B(_07626_),
    .Y(_07627_));
 sky130_fd_sc_hd__o21ba_1 _15555_ (.A1(net1273),
    .A2(_07496_),
    .B1_N(_07500_),
    .X(_07628_));
 sky130_fd_sc_hd__a21oi_1 _15556_ (.A1(net1273),
    .A2(_07496_),
    .B1(_07628_),
    .Y(_07629_));
 sky130_fd_sc_hd__nand2_1 _15557_ (.A(net2703),
    .B(net3407),
    .Y(_07630_));
 sky130_fd_sc_hd__xor2_1 _15558_ (.A(_07629_),
    .B(_07630_),
    .X(_07631_));
 sky130_fd_sc_hd__o21ba_1 _15559_ (.A1(_07541_),
    .A2(_07502_),
    .B1_N(_07504_),
    .X(_07632_));
 sky130_fd_sc_hd__a21o_1 _15560_ (.A1(_07541_),
    .A2(_07502_),
    .B1(_07632_),
    .X(_07633_));
 sky130_fd_sc_hd__xor2_1 _15561_ (.A(_07631_),
    .B(_07633_),
    .X(_07634_));
 sky130_fd_sc_hd__xnor2_1 _15562_ (.A(_07627_),
    .B(_07634_),
    .Y(_07635_));
 sky130_fd_sc_hd__and2_1 _15563_ (.A(_07569_),
    .B(_07635_),
    .X(_07636_));
 sky130_fd_sc_hd__nor2_1 _15564_ (.A(_07569_),
    .B(_07635_),
    .Y(_07637_));
 sky130_fd_sc_hd__or2_1 _15565_ (.A(_07636_),
    .B(_07637_),
    .X(_07638_));
 sky130_fd_sc_hd__xnor2_1 _15566_ (.A(net674),
    .B(_07638_),
    .Y(_07639_));
 sky130_fd_sc_hd__xnor2_1 _15567_ (.A(net574),
    .B(_07639_),
    .Y(_07640_));
 sky130_fd_sc_hd__mux2_1 _15568_ (.A0(\matmul0.matmul_stage_inst.mult1[1] ),
    .A1(net440),
    .S(net2678),
    .X(_07641_));
 sky130_fd_sc_hd__clkbuf_1 _15569_ (.A(_07641_),
    .X(_00216_));
 sky130_fd_sc_hd__a21oi_1 _15570_ (.A1(_07569_),
    .A2(_07635_),
    .B1(net674),
    .Y(_07642_));
 sky130_fd_sc_hd__and2b_1 _15571_ (.A_N(_07633_),
    .B(_07631_),
    .X(_07643_));
 sky130_fd_sc_hd__or2b_1 _15572_ (.A(_07631_),
    .B_N(_07633_),
    .X(_07644_));
 sky130_fd_sc_hd__o21ai_2 _15573_ (.A1(_07627_),
    .A2(_07643_),
    .B1(_07644_),
    .Y(_07645_));
 sky130_fd_sc_hd__nor2_1 _15574_ (.A(_07629_),
    .B(_07630_),
    .Y(_07646_));
 sky130_fd_sc_hd__nor2_1 _15575_ (.A(net2799),
    .B(net3427),
    .Y(_07647_));
 sky130_fd_sc_hd__nand2_1 _15576_ (.A(net2830),
    .B(net3488),
    .Y(_07648_));
 sky130_fd_sc_hd__nor2_1 _15577_ (.A(net2837),
    .B(net3440),
    .Y(_07649_));
 sky130_fd_sc_hd__xor2_1 _15578_ (.A(_07648_),
    .B(_07649_),
    .X(_07650_));
 sky130_fd_sc_hd__xnor2_1 _15579_ (.A(_07647_),
    .B(_07650_),
    .Y(_07651_));
 sky130_fd_sc_hd__a31o_1 _15580_ (.A1(net2833),
    .A2(net3489),
    .A3(net2677),
    .B1(_07580_),
    .X(_07652_));
 sky130_fd_sc_hd__o21a_1 _15581_ (.A1(_07476_),
    .A2(net2677),
    .B1(_07652_),
    .X(_07653_));
 sky130_fd_sc_hd__o22a_1 _15582_ (.A1(net4160),
    .A2(net4156),
    .B1(net4098),
    .B2(net4096),
    .X(_07654_));
 sky130_fd_sc_hd__nor2_1 _15583_ (.A(net3455),
    .B(net3556),
    .Y(_07655_));
 sky130_fd_sc_hd__nor2_1 _15584_ (.A(net2805),
    .B(net3466),
    .Y(_07656_));
 sky130_fd_sc_hd__xnor2_1 _15585_ (.A(_07655_),
    .B(_07656_),
    .Y(_07657_));
 sky130_fd_sc_hd__xnor2_2 _15586_ (.A(net3398),
    .B(_07657_),
    .Y(_07658_));
 sky130_fd_sc_hd__xor2_1 _15587_ (.A(net1852),
    .B(_07658_),
    .X(_07659_));
 sky130_fd_sc_hd__xnor2_1 _15588_ (.A(_07651_),
    .B(_07659_),
    .Y(_07660_));
 sky130_fd_sc_hd__a21o_1 _15589_ (.A1(net1859),
    .A2(_07582_),
    .B1(_07576_),
    .X(_07661_));
 sky130_fd_sc_hd__o21a_1 _15590_ (.A1(net1859),
    .A2(_07582_),
    .B1(_07661_),
    .X(_07662_));
 sky130_fd_sc_hd__nor2_1 _15591_ (.A(net1854),
    .B(net1853),
    .Y(_07663_));
 sky130_fd_sc_hd__nand2_1 _15592_ (.A(net1854),
    .B(net1853),
    .Y(_07664_));
 sky130_fd_sc_hd__o21ai_1 _15593_ (.A1(_07617_),
    .A2(_07663_),
    .B1(_07664_),
    .Y(_07665_));
 sky130_fd_sc_hd__xor2_1 _15594_ (.A(net1269),
    .B(net1268),
    .X(_07666_));
 sky130_fd_sc_hd__xnor2_2 _15595_ (.A(net1108),
    .B(_07666_),
    .Y(_07667_));
 sky130_fd_sc_hd__a21o_1 _15596_ (.A1(net1109),
    .A2(_07623_),
    .B1(net1270),
    .X(_07668_));
 sky130_fd_sc_hd__o21a_1 _15597_ (.A1(net1109),
    .A2(_07623_),
    .B1(_07668_),
    .X(_07669_));
 sky130_fd_sc_hd__nor2_1 _15598_ (.A(net3447),
    .B(net3537),
    .Y(_07670_));
 sky130_fd_sc_hd__nor2_1 _15599_ (.A(net3531),
    .B(net2725),
    .Y(_07671_));
 sky130_fd_sc_hd__nor2_1 _15600_ (.A(net3551),
    .B(net3514),
    .Y(_07672_));
 sky130_fd_sc_hd__xnor2_1 _15601_ (.A(_07671_),
    .B(_07672_),
    .Y(_07673_));
 sky130_fd_sc_hd__xnor2_1 _15602_ (.A(net2676),
    .B(_07673_),
    .Y(_07674_));
 sky130_fd_sc_hd__a21o_1 _15603_ (.A1(net2687),
    .A2(_07670_),
    .B1(_07593_),
    .X(_07675_));
 sky130_fd_sc_hd__o21a_1 _15604_ (.A1(_07594_),
    .A2(_07595_),
    .B1(_07675_),
    .X(_07676_));
 sky130_fd_sc_hd__a21o_1 _15605_ (.A1(_07613_),
    .A2(_07615_),
    .B1(_07614_),
    .X(_07677_));
 sky130_fd_sc_hd__o21a_1 _15606_ (.A1(_07613_),
    .A2(_07615_),
    .B1(_07677_),
    .X(_07678_));
 sky130_fd_sc_hd__xnor2_1 _15607_ (.A(net1851),
    .B(net1537),
    .Y(_07679_));
 sky130_fd_sc_hd__xnor2_1 _15608_ (.A(_07674_),
    .B(_07679_),
    .Y(_07680_));
 sky130_fd_sc_hd__a22oi_1 _15609_ (.A1(\matmul0.matmul_stage_inst.e[15] ),
    .A2(_07151_),
    .B1(_07152_),
    .B2(net7378),
    .Y(_07681_));
 sky130_fd_sc_hd__a22oi_1 _15610_ (.A1(net6542),
    .A2(\matmul0.matmul_stage_inst.c[14] ),
    .B1(\matmul0.matmul_stage_inst.b[14] ),
    .B2(net6614),
    .Y(_07682_));
 sky130_fd_sc_hd__a22o_1 _15611_ (.A1(net6542),
    .A2(\matmul0.matmul_stage_inst.c[15] ),
    .B1(\matmul0.matmul_stage_inst.b[15] ),
    .B2(net6615),
    .X(_07683_));
 sky130_fd_sc_hd__inv_2 _15612_ (.A(net4069),
    .Y(_07684_));
 sky130_fd_sc_hd__a2bb2o_1 _15613_ (.A1_N(net2851),
    .A2_N(net4076),
    .B1(net3397),
    .B2(net3444),
    .X(_07685_));
 sky130_fd_sc_hd__or2_1 _15614_ (.A(net4076),
    .B(net4069),
    .X(_07686_));
 sky130_fd_sc_hd__nand2_1 _15615_ (.A(net2851),
    .B(_07686_),
    .Y(_07687_));
 sky130_fd_sc_hd__a21o_1 _15616_ (.A1(net4074),
    .A2(net4069),
    .B1(net4075),
    .X(_07688_));
 sky130_fd_sc_hd__and2_1 _15617_ (.A(net3444),
    .B(_07688_),
    .X(_07689_));
 sky130_fd_sc_hd__a221o_1 _15618_ (.A1(net4072),
    .A2(_07685_),
    .B1(_07687_),
    .B2(net3527),
    .C1(_07689_),
    .X(_07690_));
 sky130_fd_sc_hd__xnor2_1 _15619_ (.A(net2675),
    .B(_07690_),
    .Y(_07691_));
 sky130_fd_sc_hd__or2_1 _15620_ (.A(net4075),
    .B(net4074),
    .X(_07692_));
 sky130_fd_sc_hd__a21o_1 _15621_ (.A1(net2851),
    .A2(_07692_),
    .B1(_07605_),
    .X(_07693_));
 sky130_fd_sc_hd__buf_1 _15622_ (.A(_07692_),
    .X(_07694_));
 sky130_fd_sc_hd__and3_1 _15623_ (.A(_07377_),
    .B(_07694_),
    .C(_07605_),
    .X(_07695_));
 sky130_fd_sc_hd__a21o_1 _15624_ (.A1(_07606_),
    .A2(_07693_),
    .B1(_07695_),
    .X(_07696_));
 sky130_fd_sc_hd__nand2_1 _15625_ (.A(net2813),
    .B(_07511_),
    .Y(_07697_));
 sky130_fd_sc_hd__o22a_1 _15626_ (.A1(net3597),
    .A2(net3591),
    .B1(net4083),
    .B2(net4081),
    .X(_07698_));
 sky130_fd_sc_hd__o22a_1 _15627_ (.A1(net3513),
    .A2(net3508),
    .B1(net4216),
    .B2(net4214),
    .X(_07699_));
 sky130_fd_sc_hd__xor2_1 _15628_ (.A(_07698_),
    .B(_07699_),
    .X(_07700_));
 sky130_fd_sc_hd__xnor2_1 _15629_ (.A(_07697_),
    .B(_07700_),
    .Y(_07701_));
 sky130_fd_sc_hd__xnor2_1 _15630_ (.A(_07696_),
    .B(_07701_),
    .Y(_07702_));
 sky130_fd_sc_hd__xnor2_1 _15631_ (.A(_07691_),
    .B(_07702_),
    .Y(_07703_));
 sky130_fd_sc_hd__or2_1 _15632_ (.A(net1857),
    .B(_07608_),
    .X(_07704_));
 sky130_fd_sc_hd__and2_1 _15633_ (.A(net1857),
    .B(_07608_),
    .X(_07705_));
 sky130_fd_sc_hd__a21o_1 _15634_ (.A1(_07597_),
    .A2(_07704_),
    .B1(_07705_),
    .X(_07706_));
 sky130_fd_sc_hd__xor2_1 _15635_ (.A(net1104),
    .B(net1266),
    .X(_07707_));
 sky130_fd_sc_hd__xnor2_1 _15636_ (.A(_07680_),
    .B(_07707_),
    .Y(_07708_));
 sky130_fd_sc_hd__xor2_1 _15637_ (.A(net888),
    .B(_07708_),
    .X(_07709_));
 sky130_fd_sc_hd__xnor2_1 _15638_ (.A(_07667_),
    .B(_07709_),
    .Y(_07710_));
 sky130_fd_sc_hd__a21o_1 _15639_ (.A1(_07590_),
    .A2(_07625_),
    .B1(net889),
    .X(_07711_));
 sky130_fd_sc_hd__o21ai_2 _15640_ (.A1(_07590_),
    .A2(_07625_),
    .B1(_07711_),
    .Y(_07712_));
 sky130_fd_sc_hd__a22o_1 _15641_ (.A1(\matmul0.matmul_stage_inst.e[15] ),
    .A2(_07151_),
    .B1(_07152_),
    .B2(net7378),
    .X(_07713_));
 sky130_fd_sc_hd__or2_1 _15642_ (.A(_07572_),
    .B(_07573_),
    .X(_07714_));
 sky130_fd_sc_hd__clkbuf_1 _15643_ (.A(_07714_),
    .X(_07715_));
 sky130_fd_sc_hd__and3_1 _15644_ (.A(net2821),
    .B(net3426),
    .C(net2696),
    .X(_07716_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _15645_ (.A(_07716_),
    .X(_07717_));
 sky130_fd_sc_hd__xnor2_1 _15646_ (.A(net2661),
    .B(_07717_),
    .Y(_07718_));
 sky130_fd_sc_hd__a221o_1 _15647_ (.A1(_07570_),
    .A2(net3405),
    .B1(net2666),
    .B2(net2776),
    .C1(net2781),
    .X(_07719_));
 sky130_fd_sc_hd__or2_1 _15648_ (.A(net2696),
    .B(_07570_),
    .X(_07720_));
 sky130_fd_sc_hd__or3_1 _15649_ (.A(net2250),
    .B(net2666),
    .C(_07717_),
    .X(_07721_));
 sky130_fd_sc_hd__o21ai_1 _15650_ (.A1(net2776),
    .A2(_07720_),
    .B1(_07721_),
    .Y(_07722_));
 sky130_fd_sc_hd__nor2_1 _15651_ (.A(net4079),
    .B(net4077),
    .Y(_07723_));
 sky130_fd_sc_hd__buf_1 _15652_ (.A(net3393),
    .X(_07724_));
 sky130_fd_sc_hd__o211a_1 _15653_ (.A1(net2250),
    .A2(net2672),
    .B1(_07717_),
    .C1(_07724_),
    .X(_07725_));
 sky130_fd_sc_hd__a211o_1 _15654_ (.A1(net2661),
    .A2(_07722_),
    .B1(_07725_),
    .C1(net2755),
    .X(_07726_));
 sky130_fd_sc_hd__a32o_1 _15655_ (.A1(net2776),
    .A2(net2666),
    .A3(_07718_),
    .B1(_07719_),
    .B2(_07726_),
    .X(_07727_));
 sky130_fd_sc_hd__o21ba_1 _15656_ (.A1(_07584_),
    .A2(_07588_),
    .B1_N(net1272),
    .X(_07728_));
 sky130_fd_sc_hd__a21oi_1 _15657_ (.A1(_07584_),
    .A2(_07588_),
    .B1(_07728_),
    .Y(_07729_));
 sky130_fd_sc_hd__nand2_1 _15658_ (.A(net988),
    .B(_07729_),
    .Y(_07730_));
 sky130_fd_sc_hd__or2_1 _15659_ (.A(net988),
    .B(_07729_),
    .X(_07731_));
 sky130_fd_sc_hd__nand2_1 _15660_ (.A(_07730_),
    .B(_07731_),
    .Y(_07732_));
 sky130_fd_sc_hd__xnor2_1 _15661_ (.A(_07712_),
    .B(_07732_),
    .Y(_07733_));
 sky130_fd_sc_hd__xnor2_1 _15662_ (.A(_07710_),
    .B(_07733_),
    .Y(_07734_));
 sky130_fd_sc_hd__xor2_1 _15663_ (.A(net778),
    .B(_07734_),
    .X(_07735_));
 sky130_fd_sc_hd__xnor2_1 _15664_ (.A(_07645_),
    .B(_07735_),
    .Y(_07736_));
 sky130_fd_sc_hd__a211o_1 _15665_ (.A1(net574),
    .A2(_07642_),
    .B1(_07736_),
    .C1(_07637_),
    .X(_07737_));
 sky130_fd_sc_hd__a21o_1 _15666_ (.A1(net574),
    .A2(_07642_),
    .B1(_07637_),
    .X(_07738_));
 sky130_fd_sc_hd__nand2_1 _15667_ (.A(_07736_),
    .B(_07738_),
    .Y(_07739_));
 sky130_fd_sc_hd__and2_1 _15668_ (.A(_07737_),
    .B(_07739_),
    .X(_07740_));
 sky130_fd_sc_hd__mux2_1 _15669_ (.A0(\matmul0.matmul_stage_inst.mult1[2] ),
    .A1(net433),
    .S(net2678),
    .X(_07741_));
 sky130_fd_sc_hd__clkbuf_1 _15670_ (.A(_07741_),
    .X(_00217_));
 sky130_fd_sc_hd__nor2_1 _15671_ (.A(_07696_),
    .B(_07701_),
    .Y(_07742_));
 sky130_fd_sc_hd__nand2_1 _15672_ (.A(_07696_),
    .B(_07701_),
    .Y(_07743_));
 sky130_fd_sc_hd__o21ai_1 _15673_ (.A1(_07691_),
    .A2(_07742_),
    .B1(_07743_),
    .Y(_07744_));
 sky130_fd_sc_hd__xnor2_1 _15674_ (.A(net2701),
    .B(net3526),
    .Y(_07745_));
 sky130_fd_sc_hd__nor2_1 _15675_ (.A(net2761),
    .B(_07745_),
    .Y(_07746_));
 sky130_fd_sc_hd__a2bb2o_1 _15676_ (.A1_N(net2699),
    .A2_N(_07601_),
    .B1(net4071),
    .B2(_07746_),
    .X(_07747_));
 sky130_fd_sc_hd__o21a_1 _15677_ (.A1(net2761),
    .A2(net3399),
    .B1(_07745_),
    .X(_07748_));
 sky130_fd_sc_hd__a221o_1 _15678_ (.A1(net3395),
    .A2(_07746_),
    .B1(_07747_),
    .B2(net3397),
    .C1(_07748_),
    .X(_07749_));
 sky130_fd_sc_hd__a22o_1 _15679_ (.A1(net2671),
    .A2(net2668),
    .B1(net3395),
    .B2(net2235),
    .X(_07750_));
 sky130_fd_sc_hd__a2bb2o_1 _15680_ (.A1_N(net2674),
    .A2_N(_07687_),
    .B1(_07750_),
    .B2(net2728),
    .X(_07751_));
 sky130_fd_sc_hd__nor2_2 _15681_ (.A(net3498),
    .B(net3413),
    .Y(_07752_));
 sky130_fd_sc_hd__nor2_1 _15682_ (.A(net3447),
    .B(net3600),
    .Y(_07753_));
 sky130_fd_sc_hd__nor2_1 _15683_ (.A(net2717),
    .B(net3434),
    .Y(_07754_));
 sky130_fd_sc_hd__xnor2_1 _15684_ (.A(_07753_),
    .B(_07754_),
    .Y(_07755_));
 sky130_fd_sc_hd__xnor2_2 _15685_ (.A(_07752_),
    .B(_07755_),
    .Y(_07756_));
 sky130_fd_sc_hd__xor2_1 _15686_ (.A(net1536),
    .B(_07756_),
    .X(_07757_));
 sky130_fd_sc_hd__xnor2_1 _15687_ (.A(_07749_),
    .B(_07757_),
    .Y(_07758_));
 sky130_fd_sc_hd__buf_1 _15688_ (.A(net3537),
    .X(_07759_));
 sky130_fd_sc_hd__nor2_1 _15689_ (.A(net3550),
    .B(_07759_),
    .Y(_07760_));
 sky130_fd_sc_hd__buf_1 _15690_ (.A(net3517),
    .X(_07761_));
 sky130_fd_sc_hd__nor2_1 _15691_ (.A(net2724),
    .B(_07761_),
    .Y(_07762_));
 sky130_fd_sc_hd__buf_1 _15692_ (.A(net3556),
    .X(_07763_));
 sky130_fd_sc_hd__nor2_1 _15693_ (.A(net2694),
    .B(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__xnor2_1 _15694_ (.A(_07762_),
    .B(_07764_),
    .Y(_07765_));
 sky130_fd_sc_hd__xnor2_1 _15695_ (.A(_07760_),
    .B(_07765_),
    .Y(_07766_));
 sky130_fd_sc_hd__a21o_1 _15696_ (.A1(net2676),
    .A2(_07672_),
    .B1(_07671_),
    .X(_07767_));
 sky130_fd_sc_hd__o21a_1 _15697_ (.A1(net2676),
    .A2(_07672_),
    .B1(_07767_),
    .X(_07768_));
 sky130_fd_sc_hd__nor2_1 _15698_ (.A(net2720),
    .B(net3414),
    .Y(_07769_));
 sky130_fd_sc_hd__a21bo_1 _15699_ (.A1(_07518_),
    .A2(_07769_),
    .B1_N(_07697_),
    .X(_07770_));
 sky130_fd_sc_hd__o21a_1 _15700_ (.A1(_07698_),
    .A2(_07699_),
    .B1(_07770_),
    .X(_07771_));
 sky130_fd_sc_hd__xnor2_1 _15701_ (.A(_07768_),
    .B(net1530),
    .Y(_07772_));
 sky130_fd_sc_hd__xnor2_1 _15702_ (.A(net1535),
    .B(_07772_),
    .Y(_07773_));
 sky130_fd_sc_hd__xor2_1 _15703_ (.A(net1097),
    .B(_07773_),
    .X(_07774_));
 sky130_fd_sc_hd__xnor2_2 _15704_ (.A(net1099),
    .B(_07774_),
    .Y(_07775_));
 sky130_fd_sc_hd__a21bo_1 _15705_ (.A1(_07680_),
    .A2(net1266),
    .B1_N(net1104),
    .X(_07776_));
 sky130_fd_sc_hd__o21ai_1 _15706_ (.A1(_07680_),
    .A2(net1266),
    .B1(_07776_),
    .Y(_07777_));
 sky130_fd_sc_hd__nor2_1 _15707_ (.A(net3458),
    .B(net2766),
    .Y(_07778_));
 sky130_fd_sc_hd__nor2_1 _15708_ (.A(net2804),
    .B(net3481),
    .Y(_07779_));
 sky130_fd_sc_hd__clkbuf_1 _15709_ (.A(net3454),
    .X(_07780_));
 sky130_fd_sc_hd__nor2_1 _15710_ (.A(net2647),
    .B(net3465),
    .Y(_07781_));
 sky130_fd_sc_hd__xor2_1 _15711_ (.A(_07779_),
    .B(_07781_),
    .X(_07782_));
 sky130_fd_sc_hd__xnor2_2 _15712_ (.A(_07778_),
    .B(_07782_),
    .Y(_07783_));
 sky130_fd_sc_hd__a32o_1 _15713_ (.A1(net2735),
    .A2(_07133_),
    .A3(net3398),
    .B1(net3411),
    .B2(net2685),
    .X(_07784_));
 sky130_fd_sc_hd__o21a_1 _15714_ (.A1(net3398),
    .A2(_07656_),
    .B1(_07784_),
    .X(_07785_));
 sky130_fd_sc_hd__o22a_1 _15715_ (.A1(net3585),
    .A2(net3578),
    .B1(net4087),
    .B2(net4086),
    .X(_07786_));
 sky130_fd_sc_hd__o22a_1 _15716_ (.A1(net3574),
    .A2(net3570),
    .B1(net4095),
    .B2(net4094),
    .X(_07787_));
 sky130_fd_sc_hd__xnor2_1 _15717_ (.A(_07786_),
    .B(_07787_),
    .Y(_07788_));
 sky130_fd_sc_hd__nor2_1 _15718_ (.A(net2799),
    .B(net3392),
    .Y(_07789_));
 sky130_fd_sc_hd__xnor2_2 _15719_ (.A(net2225),
    .B(_07789_),
    .Y(_07790_));
 sky130_fd_sc_hd__xnor2_1 _15720_ (.A(_07785_),
    .B(_07790_),
    .Y(_07791_));
 sky130_fd_sc_hd__xnor2_2 _15721_ (.A(_07783_),
    .B(_07791_),
    .Y(_07792_));
 sky130_fd_sc_hd__o21a_1 _15722_ (.A1(net1852),
    .A2(_07658_),
    .B1(_07651_),
    .X(_07793_));
 sky130_fd_sc_hd__a21o_1 _15723_ (.A1(net1852),
    .A2(_07658_),
    .B1(_07793_),
    .X(_07794_));
 sky130_fd_sc_hd__o21a_1 _15724_ (.A1(net1851),
    .A2(net1537),
    .B1(_07674_),
    .X(_07795_));
 sky130_fd_sc_hd__a21o_1 _15725_ (.A1(net1851),
    .A2(net1537),
    .B1(_07795_),
    .X(_07796_));
 sky130_fd_sc_hd__xnor2_1 _15726_ (.A(_07794_),
    .B(_07796_),
    .Y(_07797_));
 sky130_fd_sc_hd__xnor2_2 _15727_ (.A(_07792_),
    .B(_07797_),
    .Y(_07798_));
 sky130_fd_sc_hd__xnor2_1 _15728_ (.A(net887),
    .B(_07798_),
    .Y(_07799_));
 sky130_fd_sc_hd__xnor2_2 _15729_ (.A(_07775_),
    .B(_07799_),
    .Y(_07800_));
 sky130_fd_sc_hd__o21a_1 _15730_ (.A1(net888),
    .A2(_07667_),
    .B1(_07708_),
    .X(_07801_));
 sky130_fd_sc_hd__a21oi_2 _15731_ (.A1(net888),
    .A2(_07667_),
    .B1(_07801_),
    .Y(_07802_));
 sky130_fd_sc_hd__a21bo_1 _15732_ (.A1(net1269),
    .A2(net1268),
    .B1_N(net1108),
    .X(_07803_));
 sky130_fd_sc_hd__o21a_1 _15733_ (.A1(net1269),
    .A2(net1268),
    .B1(_07803_),
    .X(_07804_));
 sky130_fd_sc_hd__nor2_1 _15734_ (.A(net2661),
    .B(_07717_),
    .Y(_07805_));
 sky130_fd_sc_hd__a21oi_1 _15735_ (.A1(net2250),
    .A2(_07720_),
    .B1(_07717_),
    .Y(_07806_));
 sky130_fd_sc_hd__o32a_1 _15736_ (.A1(net2250),
    .A2(net2672),
    .A3(_07805_),
    .B1(_07806_),
    .B2(_07724_),
    .X(_07807_));
 sky130_fd_sc_hd__a21bo_1 _15737_ (.A1(_07647_),
    .A2(_07649_),
    .B1_N(_07648_),
    .X(_07808_));
 sky130_fd_sc_hd__o21a_1 _15738_ (.A1(_07647_),
    .A2(_07649_),
    .B1(_07808_),
    .X(_07809_));
 sky130_fd_sc_hd__clkbuf_1 _15739_ (.A(net2672),
    .X(_07810_));
 sky130_fd_sc_hd__nor2_1 _15740_ (.A(net2780),
    .B(net2221),
    .Y(_07811_));
 sky130_fd_sc_hd__xnor2_1 _15741_ (.A(net1529),
    .B(net1850),
    .Y(_07812_));
 sky130_fd_sc_hd__o21ai_1 _15742_ (.A1(net2758),
    .A2(net1265),
    .B1(_07812_),
    .Y(_07813_));
 sky130_fd_sc_hd__inv_2 _15743_ (.A(_07813_),
    .Y(_07814_));
 sky130_fd_sc_hd__nor3_1 _15744_ (.A(net2758),
    .B(_07812_),
    .C(net1265),
    .Y(_07815_));
 sky130_fd_sc_hd__nor2_1 _15745_ (.A(_07814_),
    .B(_07815_),
    .Y(_07816_));
 sky130_fd_sc_hd__xnor2_2 _15746_ (.A(_07804_),
    .B(_07816_),
    .Y(_07817_));
 sky130_fd_sc_hd__xor2_1 _15747_ (.A(_07802_),
    .B(_07817_),
    .X(_07818_));
 sky130_fd_sc_hd__xnor2_2 _15748_ (.A(_07800_),
    .B(_07818_),
    .Y(_07819_));
 sky130_fd_sc_hd__o21a_1 _15749_ (.A1(_07712_),
    .A2(_07732_),
    .B1(_07710_),
    .X(_07820_));
 sky130_fd_sc_hd__a21o_1 _15750_ (.A1(_07712_),
    .A2(_07732_),
    .B1(_07820_),
    .X(_07821_));
 sky130_fd_sc_hd__xnor2_1 _15751_ (.A(_07819_),
    .B(_07821_),
    .Y(_07822_));
 sky130_fd_sc_hd__xnor2_1 _15752_ (.A(_07730_),
    .B(_07822_),
    .Y(_07823_));
 sky130_fd_sc_hd__nor2_1 _15753_ (.A(_07645_),
    .B(_07734_),
    .Y(_07824_));
 sky130_fd_sc_hd__a21boi_1 _15754_ (.A1(_07645_),
    .A2(_07734_),
    .B1_N(net778),
    .Y(_07825_));
 sky130_fd_sc_hd__or3_1 _15755_ (.A(_07823_),
    .B(_07824_),
    .C(_07825_),
    .X(_07826_));
 sky130_fd_sc_hd__o21ai_1 _15756_ (.A1(_07824_),
    .A2(_07825_),
    .B1(_07823_),
    .Y(_07827_));
 sky130_fd_sc_hd__nand2_1 _15757_ (.A(_07826_),
    .B(_07827_),
    .Y(_07828_));
 sky130_fd_sc_hd__xor2_1 _15758_ (.A(_07737_),
    .B(_07828_),
    .X(_07829_));
 sky130_fd_sc_hd__mux2_1 _15759_ (.A0(\matmul0.matmul_stage_inst.mult1[3] ),
    .A1(net426),
    .S(net2680),
    .X(_07830_));
 sky130_fd_sc_hd__clkbuf_1 _15760_ (.A(_07830_),
    .X(_00218_));
 sky130_fd_sc_hd__a21boi_1 _15761_ (.A1(_07737_),
    .A2(_07827_),
    .B1_N(_07826_),
    .Y(_07831_));
 sky130_fd_sc_hd__a21bo_1 _15762_ (.A1(net1536),
    .A2(_07756_),
    .B1_N(_07749_),
    .X(_07832_));
 sky130_fd_sc_hd__o21ai_1 _15763_ (.A1(net1536),
    .A2(_07756_),
    .B1(_07832_),
    .Y(_07833_));
 sky130_fd_sc_hd__nor2_1 _15764_ (.A(net3499),
    .B(net3399),
    .Y(_07834_));
 sky130_fd_sc_hd__nor2_1 _15765_ (.A(net3449),
    .B(net3438),
    .Y(_07835_));
 sky130_fd_sc_hd__xnor2_1 _15766_ (.A(_07769_),
    .B(_07835_),
    .Y(_07836_));
 sky130_fd_sc_hd__xnor2_2 _15767_ (.A(_07834_),
    .B(_07836_),
    .Y(_07837_));
 sky130_fd_sc_hd__buf_1 _15768_ (.A(net3400),
    .X(_07838_));
 sky130_fd_sc_hd__a21oi_1 _15769_ (.A1(net2700),
    .A2(net2671),
    .B1(net3526),
    .Y(_07839_));
 sky130_fd_sc_hd__a21oi_1 _15770_ (.A1(net2234),
    .A2(_07838_),
    .B1(_07839_),
    .Y(_07840_));
 sky130_fd_sc_hd__nor2_1 _15771_ (.A(net2699),
    .B(net2727),
    .Y(_07841_));
 sky130_fd_sc_hd__nand2_1 _15772_ (.A(net2700),
    .B(_07841_),
    .Y(_07842_));
 sky130_fd_sc_hd__clkbuf_1 _15773_ (.A(net3396),
    .X(_07843_));
 sky130_fd_sc_hd__o211a_1 _15774_ (.A1(net2761),
    .A2(_07840_),
    .B1(_07842_),
    .C1(net2640),
    .X(_07844_));
 sky130_fd_sc_hd__xor2_1 _15775_ (.A(_07837_),
    .B(_07844_),
    .X(_07845_));
 sky130_fd_sc_hd__nor2_1 _15776_ (.A(net3550),
    .B(net3600),
    .Y(_07846_));
 sky130_fd_sc_hd__o22a_1 _15777_ (.A1(net4138),
    .A2(net4131),
    .B1(net4198),
    .B2(net4197),
    .X(_07847_));
 sky130_fd_sc_hd__nor2_1 _15778_ (.A(net2650),
    .B(_07761_),
    .Y(_07848_));
 sky130_fd_sc_hd__xnor2_1 _15779_ (.A(net3390),
    .B(_07848_),
    .Y(_07849_));
 sky130_fd_sc_hd__xnor2_1 _15780_ (.A(_07846_),
    .B(_07849_),
    .Y(_07850_));
 sky130_fd_sc_hd__o21a_1 _15781_ (.A1(_07762_),
    .A2(_07764_),
    .B1(_07760_),
    .X(_07851_));
 sky130_fd_sc_hd__a21o_1 _15782_ (.A1(_07762_),
    .A2(_07764_),
    .B1(_07851_),
    .X(_07852_));
 sky130_fd_sc_hd__a21o_1 _15783_ (.A1(_07752_),
    .A2(_07753_),
    .B1(_07754_),
    .X(_07853_));
 sky130_fd_sc_hd__o21a_1 _15784_ (.A1(_07752_),
    .A2(_07753_),
    .B1(_07853_),
    .X(_07854_));
 sky130_fd_sc_hd__xnor2_1 _15785_ (.A(_07852_),
    .B(_07854_),
    .Y(_07855_));
 sky130_fd_sc_hd__xnor2_1 _15786_ (.A(_07850_),
    .B(_07855_),
    .Y(_07856_));
 sky130_fd_sc_hd__nor2_1 _15787_ (.A(net1264),
    .B(_07856_),
    .Y(_07857_));
 sky130_fd_sc_hd__nand2_1 _15788_ (.A(net1264),
    .B(_07856_),
    .Y(_07858_));
 sky130_fd_sc_hd__or2b_1 _15789_ (.A(_07857_),
    .B_N(_07858_),
    .X(_07859_));
 sky130_fd_sc_hd__xnor2_1 _15790_ (.A(net987),
    .B(_07859_),
    .Y(_07860_));
 sky130_fd_sc_hd__o21a_1 _15791_ (.A1(net1097),
    .A2(_07773_),
    .B1(net1099),
    .X(_07861_));
 sky130_fd_sc_hd__a21o_1 _15792_ (.A1(net1097),
    .A2(_07773_),
    .B1(_07861_),
    .X(_07862_));
 sky130_fd_sc_hd__nor2_1 _15793_ (.A(net2836),
    .B(net2658),
    .Y(_07863_));
 sky130_fd_sc_hd__buf_1 _15794_ (.A(net3439),
    .X(_07864_));
 sky130_fd_sc_hd__nor2_1 _15795_ (.A(net3458),
    .B(_07864_),
    .Y(_07865_));
 sky130_fd_sc_hd__buf_1 _15796_ (.A(net3427),
    .X(_07866_));
 sky130_fd_sc_hd__nor2_1 _15797_ (.A(net3546),
    .B(_07866_),
    .Y(_07867_));
 sky130_fd_sc_hd__xnor2_1 _15798_ (.A(_07865_),
    .B(_07867_),
    .Y(_07868_));
 sky130_fd_sc_hd__xnor2_2 _15799_ (.A(_07863_),
    .B(_07868_),
    .Y(_07869_));
 sky130_fd_sc_hd__a21o_1 _15800_ (.A1(_07778_),
    .A2(_07779_),
    .B1(_07781_),
    .X(_07870_));
 sky130_fd_sc_hd__o21a_1 _15801_ (.A1(_07778_),
    .A2(_07779_),
    .B1(_07870_),
    .X(_07871_));
 sky130_fd_sc_hd__nand2_1 _15802_ (.A(net2732),
    .B(net2788),
    .Y(_07872_));
 sky130_fd_sc_hd__nor2_1 _15803_ (.A(net2647),
    .B(net3481),
    .Y(_07873_));
 sky130_fd_sc_hd__nor2_1 _15804_ (.A(net2693),
    .B(net3465),
    .Y(_07874_));
 sky130_fd_sc_hd__xor2_1 _15805_ (.A(_07873_),
    .B(_07874_),
    .X(_07875_));
 sky130_fd_sc_hd__xnor2_2 _15806_ (.A(_07872_),
    .B(_07875_),
    .Y(_07876_));
 sky130_fd_sc_hd__xor2_1 _15807_ (.A(_07871_),
    .B(_07876_),
    .X(_07877_));
 sky130_fd_sc_hd__xnor2_2 _15808_ (.A(_07869_),
    .B(_07877_),
    .Y(_07878_));
 sky130_fd_sc_hd__nand2_1 _15809_ (.A(_07768_),
    .B(net1530),
    .Y(_07879_));
 sky130_fd_sc_hd__o21ai_1 _15810_ (.A1(_07768_),
    .A2(net1530),
    .B1(net1535),
    .Y(_07880_));
 sky130_fd_sc_hd__nand2_1 _15811_ (.A(_07785_),
    .B(_07790_),
    .Y(_07881_));
 sky130_fd_sc_hd__nor2_1 _15812_ (.A(_07785_),
    .B(_07790_),
    .Y(_07882_));
 sky130_fd_sc_hd__a21o_1 _15813_ (.A1(_07783_),
    .A2(_07881_),
    .B1(_07882_),
    .X(_07883_));
 sky130_fd_sc_hd__a21o_1 _15814_ (.A1(_07879_),
    .A2(_07880_),
    .B1(_07883_),
    .X(_07884_));
 sky130_fd_sc_hd__inv_2 _15815_ (.A(_07884_),
    .Y(_07885_));
 sky130_fd_sc_hd__and3_1 _15816_ (.A(_07883_),
    .B(_07879_),
    .C(_07880_),
    .X(_07886_));
 sky130_fd_sc_hd__or2_1 _15817_ (.A(_07885_),
    .B(_07886_),
    .X(_07887_));
 sky130_fd_sc_hd__xnor2_2 _15818_ (.A(_07878_),
    .B(_07887_),
    .Y(_07888_));
 sky130_fd_sc_hd__xnor2_1 _15819_ (.A(_07862_),
    .B(_07888_),
    .Y(_07889_));
 sky130_fd_sc_hd__xnor2_2 _15820_ (.A(net827),
    .B(_07889_),
    .Y(_07890_));
 sky130_fd_sc_hd__o21a_1 _15821_ (.A1(_07775_),
    .A2(_07798_),
    .B1(net887),
    .X(_07891_));
 sky130_fd_sc_hd__a21o_1 _15822_ (.A1(_07775_),
    .A2(_07798_),
    .B1(_07891_),
    .X(_07892_));
 sky130_fd_sc_hd__o21ba_1 _15823_ (.A1(_07794_),
    .A2(_07796_),
    .B1_N(_07792_),
    .X(_07893_));
 sky130_fd_sc_hd__a21oi_2 _15824_ (.A1(_07794_),
    .A2(_07796_),
    .B1(_07893_),
    .Y(_07894_));
 sky130_fd_sc_hd__nand2_1 _15825_ (.A(net1529),
    .B(net1850),
    .Y(_07895_));
 sky130_fd_sc_hd__buf_1 _15826_ (.A(net2660),
    .X(_07896_));
 sky130_fd_sc_hd__or3_1 _15827_ (.A(net2799),
    .B(net2216),
    .C(net2225),
    .X(_07897_));
 sky130_fd_sc_hd__nor2_1 _15828_ (.A(_07864_),
    .B(_07866_),
    .Y(_07898_));
 sky130_fd_sc_hd__o2bb2a_1 _15829_ (.A1_N(net3565),
    .A2_N(_07898_),
    .B1(net2221),
    .B2(net2821),
    .X(_07899_));
 sky130_fd_sc_hd__nand2_1 _15830_ (.A(net3425),
    .B(net2695),
    .Y(_07900_));
 sky130_fd_sc_hd__nor2_1 _15831_ (.A(net2223),
    .B(_07900_),
    .Y(_07901_));
 sky130_fd_sc_hd__and3_1 _15832_ (.A(net2799),
    .B(net3565),
    .C(net1846),
    .X(_07902_));
 sky130_fd_sc_hd__a21o_1 _15833_ (.A1(_07897_),
    .A2(_07899_),
    .B1(_07902_),
    .X(_07903_));
 sky130_fd_sc_hd__xnor2_1 _15834_ (.A(_07895_),
    .B(net1263),
    .Y(_07904_));
 sky130_fd_sc_hd__xnor2_1 _15835_ (.A(_07894_),
    .B(_07904_),
    .Y(_07905_));
 sky130_fd_sc_hd__and2_1 _15836_ (.A(_07892_),
    .B(_07905_),
    .X(_07906_));
 sky130_fd_sc_hd__nor2_1 _15837_ (.A(_07892_),
    .B(_07905_),
    .Y(_07907_));
 sky130_fd_sc_hd__nor2_1 _15838_ (.A(_07906_),
    .B(_07907_),
    .Y(_07908_));
 sky130_fd_sc_hd__xnor2_1 _15839_ (.A(_07890_),
    .B(_07908_),
    .Y(_07909_));
 sky130_fd_sc_hd__a21o_1 _15840_ (.A1(_07802_),
    .A2(_07817_),
    .B1(_07800_),
    .X(_07910_));
 sky130_fd_sc_hd__o21ai_2 _15841_ (.A1(_07802_),
    .A2(_07817_),
    .B1(_07910_),
    .Y(_07911_));
 sky130_fd_sc_hd__o21a_1 _15842_ (.A1(_07804_),
    .A2(_07815_),
    .B1(_07813_),
    .X(_07912_));
 sky130_fd_sc_hd__xnor2_1 _15843_ (.A(_07911_),
    .B(_07912_),
    .Y(_07913_));
 sky130_fd_sc_hd__xnor2_1 _15844_ (.A(_07909_),
    .B(_07913_),
    .Y(_07914_));
 sky130_fd_sc_hd__inv_2 _15845_ (.A(_07821_),
    .Y(_07915_));
 sky130_fd_sc_hd__nand2_1 _15846_ (.A(_07819_),
    .B(_07915_),
    .Y(_07916_));
 sky130_fd_sc_hd__nor2_1 _15847_ (.A(_07819_),
    .B(_07915_),
    .Y(_07917_));
 sky130_fd_sc_hd__a21o_1 _15848_ (.A1(_07730_),
    .A2(_07916_),
    .B1(_07917_),
    .X(_07918_));
 sky130_fd_sc_hd__nor2_1 _15849_ (.A(_07914_),
    .B(_07918_),
    .Y(_07919_));
 sky130_fd_sc_hd__nand2_1 _15850_ (.A(_07914_),
    .B(_07918_),
    .Y(_07920_));
 sky130_fd_sc_hd__or2b_1 _15851_ (.A(_07919_),
    .B_N(_07920_),
    .X(_07921_));
 sky130_fd_sc_hd__xnor2_1 _15852_ (.A(_07831_),
    .B(_07921_),
    .Y(_07922_));
 sky130_fd_sc_hd__mux2_1 _15853_ (.A0(\matmul0.matmul_stage_inst.mult1[4] ),
    .A1(net396),
    .S(net2680),
    .X(_07923_));
 sky130_fd_sc_hd__clkbuf_1 _15854_ (.A(_07923_),
    .X(_00219_));
 sky130_fd_sc_hd__o21a_1 _15855_ (.A1(_07831_),
    .A2(_07919_),
    .B1(_07920_),
    .X(_07924_));
 sky130_fd_sc_hd__o21ba_1 _15856_ (.A1(net827),
    .A2(_07888_),
    .B1_N(_07862_),
    .X(_07925_));
 sky130_fd_sc_hd__a21oi_1 _15857_ (.A1(net827),
    .A2(_07888_),
    .B1(_07925_),
    .Y(_07926_));
 sky130_fd_sc_hd__o21ai_1 _15858_ (.A1(net2234),
    .A2(net2727),
    .B1(_07837_),
    .Y(_07927_));
 sky130_fd_sc_hd__o31a_1 _15859_ (.A1(net2700),
    .A2(net2761),
    .A3(net2671),
    .B1(_07837_),
    .X(_07928_));
 sky130_fd_sc_hd__nand2_1 _15860_ (.A(net2699),
    .B(net2727),
    .Y(_07929_));
 sky130_fd_sc_hd__o21a_1 _15861_ (.A1(_07929_),
    .A2(net2671),
    .B1(_07837_),
    .X(_07930_));
 sky130_fd_sc_hd__o22ai_1 _15862_ (.A1(net2727),
    .A2(_07928_),
    .B1(_07930_),
    .B2(net2234),
    .Y(_07931_));
 sky130_fd_sc_hd__nor2_2 _15863_ (.A(net4075),
    .B(net4068),
    .Y(_07932_));
 sky130_fd_sc_hd__clkbuf_1 _15864_ (.A(_07932_),
    .X(_07933_));
 sky130_fd_sc_hd__a211o_1 _15865_ (.A1(net2761),
    .A2(_07927_),
    .B1(_07931_),
    .C1(net2630),
    .X(_07934_));
 sky130_fd_sc_hd__nor2_1 _15866_ (.A(net3550),
    .B(net3434),
    .Y(_07935_));
 sky130_fd_sc_hd__buf_1 _15867_ (.A(net3599),
    .X(_07936_));
 sky130_fd_sc_hd__nor2_1 _15868_ (.A(net2723),
    .B(net2627),
    .Y(_07937_));
 sky130_fd_sc_hd__nor2_1 _15869_ (.A(net2650),
    .B(net2657),
    .Y(_07938_));
 sky130_fd_sc_hd__xnor2_1 _15870_ (.A(_07937_),
    .B(_07938_),
    .Y(_07939_));
 sky130_fd_sc_hd__xnor2_1 _15871_ (.A(_07935_),
    .B(_07939_),
    .Y(_07940_));
 sky130_fd_sc_hd__a32o_1 _15872_ (.A1(net2842),
    .A2(net3432),
    .A3(net3390),
    .B1(net2683),
    .B2(net3523),
    .X(_07941_));
 sky130_fd_sc_hd__o21a_1 _15873_ (.A1(_07846_),
    .A2(net3390),
    .B1(_07941_),
    .X(_07942_));
 sky130_fd_sc_hd__and4_1 _15874_ (.A(net2714),
    .B(net2812),
    .C(net3422),
    .D(_07694_),
    .X(_07943_));
 sky130_fd_sc_hd__a22o_1 _15875_ (.A1(net2714),
    .A2(net3422),
    .B1(_07694_),
    .B2(net2813),
    .X(_07944_));
 sky130_fd_sc_hd__o21a_1 _15876_ (.A1(_07769_),
    .A2(_07943_),
    .B1(_07944_),
    .X(_07945_));
 sky130_fd_sc_hd__nor2_1 _15877_ (.A(net1845),
    .B(net1842),
    .Y(_07946_));
 sky130_fd_sc_hd__and2_1 _15878_ (.A(net1845),
    .B(net1842),
    .X(_07947_));
 sky130_fd_sc_hd__or2_1 _15879_ (.A(_07946_),
    .B(_07947_),
    .X(_07948_));
 sky130_fd_sc_hd__xnor2_1 _15880_ (.A(_07940_),
    .B(_07948_),
    .Y(_07949_));
 sky130_fd_sc_hd__o211a_1 _15881_ (.A1(net2700),
    .A2(_07929_),
    .B1(net3396),
    .C1(_07842_),
    .X(_07950_));
 sky130_fd_sc_hd__nor2_1 _15882_ (.A(net3448),
    .B(net3413),
    .Y(_07951_));
 sky130_fd_sc_hd__a2bb2o_1 _15883_ (.A1_N(net2810),
    .A2_N(_07601_),
    .B1(net3397),
    .B2(net2737),
    .X(_07952_));
 sky130_fd_sc_hd__nand2_1 _15884_ (.A(net2810),
    .B(_07686_),
    .Y(_07953_));
 sky130_fd_sc_hd__and2_1 _15885_ (.A(net2737),
    .B(net3395),
    .X(_07954_));
 sky130_fd_sc_hd__a221o_1 _15886_ (.A1(net4071),
    .A2(_07952_),
    .B1(_07953_),
    .B2(net2718),
    .C1(_07954_),
    .X(_07955_));
 sky130_fd_sc_hd__xor2_1 _15887_ (.A(_07951_),
    .B(_07955_),
    .X(_07956_));
 sky130_fd_sc_hd__xnor2_1 _15888_ (.A(net1525),
    .B(net1523),
    .Y(_07957_));
 sky130_fd_sc_hd__or2_1 _15889_ (.A(_07949_),
    .B(_07957_),
    .X(_07958_));
 sky130_fd_sc_hd__nand2_1 _15890_ (.A(_07949_),
    .B(_07957_),
    .Y(_07959_));
 sky130_fd_sc_hd__nand2_1 _15891_ (.A(_07958_),
    .B(_07959_),
    .Y(_07960_));
 sky130_fd_sc_hd__xor2_1 _15892_ (.A(net984),
    .B(_07960_),
    .X(_07961_));
 sky130_fd_sc_hd__o21ai_1 _15893_ (.A1(net987),
    .A2(_07857_),
    .B1(_07858_),
    .Y(_07962_));
 sky130_fd_sc_hd__nor2_1 _15894_ (.A(net2647),
    .B(net2765),
    .Y(_07963_));
 sky130_fd_sc_hd__nor2_1 _15895_ (.A(net3530),
    .B(net3481),
    .Y(_07964_));
 sky130_fd_sc_hd__nor2_1 _15896_ (.A(net3515),
    .B(net3465),
    .Y(_07965_));
 sky130_fd_sc_hd__xor2_1 _15897_ (.A(_07964_),
    .B(_07965_),
    .X(_07966_));
 sky130_fd_sc_hd__xnor2_1 _15898_ (.A(_07963_),
    .B(_07966_),
    .Y(_07967_));
 sky130_fd_sc_hd__o21ai_1 _15899_ (.A1(net2647),
    .A2(net2748),
    .B1(_07872_),
    .Y(_07968_));
 sky130_fd_sc_hd__and3_1 _15900_ (.A(net2732),
    .B(net2788),
    .C(_07873_),
    .X(_07969_));
 sky130_fd_sc_hd__a21o_1 _15901_ (.A1(_07874_),
    .A2(_07968_),
    .B1(_07969_),
    .X(_07970_));
 sky130_fd_sc_hd__a211o_1 _15902_ (.A1(net2846),
    .A2(net2695),
    .B1(net3439),
    .C1(net2803),
    .X(_07971_));
 sky130_fd_sc_hd__a211o_1 _15903_ (.A1(net2734),
    .A2(net3425),
    .B1(net3427),
    .C1(net3460),
    .X(_07972_));
 sky130_fd_sc_hd__a211o_1 _15904_ (.A1(_07971_),
    .A2(_07972_),
    .B1(net3546),
    .C1(net3392),
    .X(_07973_));
 sky130_fd_sc_hd__o211ai_1 _15905_ (.A1(net3546),
    .A2(net3392),
    .B1(_07971_),
    .C1(_07972_),
    .Y(_07974_));
 sky130_fd_sc_hd__and2_1 _15906_ (.A(_07973_),
    .B(_07974_),
    .X(_07975_));
 sky130_fd_sc_hd__xor2_1 _15907_ (.A(_07970_),
    .B(net1522),
    .X(_07976_));
 sky130_fd_sc_hd__xnor2_1 _15908_ (.A(_07967_),
    .B(_07976_),
    .Y(_07977_));
 sky130_fd_sc_hd__a21o_1 _15909_ (.A1(_07871_),
    .A2(_07876_),
    .B1(_07869_),
    .X(_07978_));
 sky130_fd_sc_hd__o21a_1 _15910_ (.A1(_07871_),
    .A2(_07876_),
    .B1(_07978_),
    .X(_07979_));
 sky130_fd_sc_hd__o21a_1 _15911_ (.A1(_07852_),
    .A2(_07854_),
    .B1(_07850_),
    .X(_07980_));
 sky130_fd_sc_hd__a21o_1 _15912_ (.A1(_07852_),
    .A2(_07854_),
    .B1(_07980_),
    .X(_07981_));
 sky130_fd_sc_hd__xnor2_1 _15913_ (.A(_07979_),
    .B(net1094),
    .Y(_07982_));
 sky130_fd_sc_hd__xnor2_1 _15914_ (.A(_07977_),
    .B(_07982_),
    .Y(_07983_));
 sky130_fd_sc_hd__or2_1 _15915_ (.A(net884),
    .B(_07983_),
    .X(_07984_));
 sky130_fd_sc_hd__nand2_1 _15916_ (.A(net884),
    .B(_07983_),
    .Y(_07985_));
 sky130_fd_sc_hd__nand2_1 _15917_ (.A(_07984_),
    .B(_07985_),
    .Y(_07986_));
 sky130_fd_sc_hd__xnor2_1 _15918_ (.A(net826),
    .B(_07986_),
    .Y(_07987_));
 sky130_fd_sc_hd__o21a_1 _15919_ (.A1(_07878_),
    .A2(_07886_),
    .B1(_07884_),
    .X(_07988_));
 sky130_fd_sc_hd__o21a_1 _15920_ (.A1(_07865_),
    .A2(_07867_),
    .B1(_07863_),
    .X(_07989_));
 sky130_fd_sc_hd__clkbuf_1 _15921_ (.A(net2666),
    .X(_07990_));
 sky130_fd_sc_hd__a32o_1 _15922_ (.A1(net2829),
    .A2(net2846),
    .A3(_07898_),
    .B1(net2212),
    .B2(net2836),
    .X(_07991_));
 sky130_fd_sc_hd__and4_1 _15923_ (.A(net2836),
    .B(net2829),
    .C(net2846),
    .D(net1846),
    .X(_07992_));
 sky130_fd_sc_hd__o21ba_1 _15924_ (.A1(_07989_),
    .A2(_07991_),
    .B1_N(_07992_),
    .X(_07993_));
 sky130_fd_sc_hd__xnor2_1 _15925_ (.A(net1527),
    .B(net1262),
    .Y(_07994_));
 sky130_fd_sc_hd__xnor2_1 _15926_ (.A(_07988_),
    .B(_07994_),
    .Y(_07995_));
 sky130_fd_sc_hd__xor2_1 _15927_ (.A(_07987_),
    .B(_07995_),
    .X(_07996_));
 sky130_fd_sc_hd__xnor2_1 _15928_ (.A(_07926_),
    .B(_07996_),
    .Y(_07997_));
 sky130_fd_sc_hd__nand2_1 _15929_ (.A(_07892_),
    .B(_07905_),
    .Y(_07998_));
 sky130_fd_sc_hd__o21ai_2 _15930_ (.A1(_07890_),
    .A2(_07907_),
    .B1(_07998_),
    .Y(_07999_));
 sky130_fd_sc_hd__o21a_1 _15931_ (.A1(_07894_),
    .A2(net1263),
    .B1(_07895_),
    .X(_08000_));
 sky130_fd_sc_hd__a21oi_1 _15932_ (.A1(_07894_),
    .A2(net1263),
    .B1(_08000_),
    .Y(_08001_));
 sky130_fd_sc_hd__xnor2_1 _15933_ (.A(_07999_),
    .B(_08001_),
    .Y(_08002_));
 sky130_fd_sc_hd__xnor2_1 _15934_ (.A(_07997_),
    .B(_08002_),
    .Y(_08003_));
 sky130_fd_sc_hd__nor2_1 _15935_ (.A(_07911_),
    .B(_07912_),
    .Y(_08004_));
 sky130_fd_sc_hd__nand2_1 _15936_ (.A(_07911_),
    .B(_07912_),
    .Y(_08005_));
 sky130_fd_sc_hd__o21a_1 _15937_ (.A1(_07909_),
    .A2(_08004_),
    .B1(_08005_),
    .X(_08006_));
 sky130_fd_sc_hd__and2_1 _15938_ (.A(_08003_),
    .B(_08006_),
    .X(_08007_));
 sky130_fd_sc_hd__nor2_1 _15939_ (.A(_08003_),
    .B(_08006_),
    .Y(_08008_));
 sky130_fd_sc_hd__or2_1 _15940_ (.A(_08007_),
    .B(_08008_),
    .X(_08009_));
 sky130_fd_sc_hd__xnor2_1 _15941_ (.A(net425),
    .B(_08009_),
    .Y(_08010_));
 sky130_fd_sc_hd__mux2_1 _15942_ (.A0(\matmul0.matmul_stage_inst.mult1[5] ),
    .A1(net389),
    .S(_07560_),
    .X(_08011_));
 sky130_fd_sc_hd__clkbuf_1 _15943_ (.A(_08011_),
    .X(_00220_));
 sky130_fd_sc_hd__or2b_1 _15944_ (.A(_07987_),
    .B_N(_07995_),
    .X(_08012_));
 sky130_fd_sc_hd__and2b_1 _15945_ (.A_N(_07995_),
    .B(_07987_),
    .X(_08013_));
 sky130_fd_sc_hd__a21oi_1 _15946_ (.A1(_07926_),
    .A2(_08012_),
    .B1(_08013_),
    .Y(_08014_));
 sky130_fd_sc_hd__a21bo_1 _15947_ (.A1(net1527),
    .A2(net1262),
    .B1_N(_07988_),
    .X(_08015_));
 sky130_fd_sc_hd__o21ai_2 _15948_ (.A1(net1527),
    .A2(net1262),
    .B1(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__inv_2 _15949_ (.A(_07958_),
    .Y(_08017_));
 sky130_fd_sc_hd__o21ai_2 _15950_ (.A1(net984),
    .A2(_08017_),
    .B1(_07959_),
    .Y(_08018_));
 sky130_fd_sc_hd__nor2_1 _15951_ (.A(net2693),
    .B(_07156_),
    .Y(_08019_));
 sky130_fd_sc_hd__nor2_1 _15952_ (.A(net2652),
    .B(net2748),
    .Y(_08020_));
 sky130_fd_sc_hd__nor2_1 _15953_ (.A(net2753),
    .B(net2653),
    .Y(_08021_));
 sky130_fd_sc_hd__xnor2_1 _15954_ (.A(_08020_),
    .B(_08021_),
    .Y(_08022_));
 sky130_fd_sc_hd__xnor2_1 _15955_ (.A(_08019_),
    .B(_08022_),
    .Y(_08023_));
 sky130_fd_sc_hd__o21a_1 _15956_ (.A1(_07963_),
    .A2(_07964_),
    .B1(_07965_),
    .X(_08024_));
 sky130_fd_sc_hd__a21o_1 _15957_ (.A1(_07963_),
    .A2(_07964_),
    .B1(_08024_),
    .X(_08025_));
 sky130_fd_sc_hd__nor2_1 _15958_ (.A(net2803),
    .B(net2633),
    .Y(_08026_));
 sky130_fd_sc_hd__nor2_1 _15959_ (.A(net3460),
    .B(net2660),
    .Y(_08027_));
 sky130_fd_sc_hd__nor2_2 _15960_ (.A(net2646),
    .B(net2637),
    .Y(_08028_));
 sky130_fd_sc_hd__xnor2_1 _15961_ (.A(_08027_),
    .B(_08028_),
    .Y(_08029_));
 sky130_fd_sc_hd__xnor2_1 _15962_ (.A(_08026_),
    .B(_08029_),
    .Y(_08030_));
 sky130_fd_sc_hd__xor2_1 _15963_ (.A(_08025_),
    .B(_08030_),
    .X(_08031_));
 sky130_fd_sc_hd__xnor2_1 _15964_ (.A(_08023_),
    .B(_08031_),
    .Y(_08032_));
 sky130_fd_sc_hd__o21ba_1 _15965_ (.A1(_07970_),
    .A2(net1522),
    .B1_N(_07967_),
    .X(_08033_));
 sky130_fd_sc_hd__a21o_1 _15966_ (.A1(_07970_),
    .A2(net1522),
    .B1(_08033_),
    .X(_08034_));
 sky130_fd_sc_hd__o21ba_1 _15967_ (.A1(_07940_),
    .A2(_07947_),
    .B1_N(_07946_),
    .X(_08035_));
 sky130_fd_sc_hd__xor2_1 _15968_ (.A(_08034_),
    .B(net1261),
    .X(_08036_));
 sky130_fd_sc_hd__xnor2_1 _15969_ (.A(_08032_),
    .B(_08036_),
    .Y(_08037_));
 sky130_fd_sc_hd__nor2_1 _15970_ (.A(net2708),
    .B(net3416),
    .Y(_08038_));
 sky130_fd_sc_hd__nor2_1 _15971_ (.A(net2649),
    .B(net2626),
    .Y(_08039_));
 sky130_fd_sc_hd__buf_1 _15972_ (.A(net3436),
    .X(_08040_));
 sky130_fd_sc_hd__nor2_1 _15973_ (.A(net2722),
    .B(net2624),
    .Y(_08041_));
 sky130_fd_sc_hd__xor2_1 _15974_ (.A(_08039_),
    .B(_08041_),
    .X(_08042_));
 sky130_fd_sc_hd__xnor2_1 _15975_ (.A(_08038_),
    .B(_08042_),
    .Y(_08043_));
 sky130_fd_sc_hd__o21ai_1 _15976_ (.A1(net2718),
    .A2(net3399),
    .B1(_07953_),
    .Y(_08044_));
 sky130_fd_sc_hd__o21a_1 _15977_ (.A1(_07951_),
    .A2(_07954_),
    .B1(_08044_),
    .X(_08045_));
 sky130_fd_sc_hd__a21o_1 _15978_ (.A1(_07935_),
    .A2(_07938_),
    .B1(_07937_),
    .X(_08046_));
 sky130_fd_sc_hd__o21a_1 _15979_ (.A1(_07935_),
    .A2(_07938_),
    .B1(_08046_),
    .X(_08047_));
 sky130_fd_sc_hd__xnor2_1 _15980_ (.A(net1518),
    .B(_08047_),
    .Y(_08048_));
 sky130_fd_sc_hd__xnor2_2 _15981_ (.A(net1520),
    .B(_08048_),
    .Y(_08049_));
 sky130_fd_sc_hd__and2_1 _15982_ (.A(net1525),
    .B(net1523),
    .X(_08050_));
 sky130_fd_sc_hd__or3b_1 _15983_ (.A(net2762),
    .B(_07932_),
    .C_N(net3444),
    .X(_08051_));
 sky130_fd_sc_hd__or2b_1 _15984_ (.A(_08050_),
    .B_N(net2205),
    .X(_08052_));
 sky130_fd_sc_hd__xnor2_2 _15985_ (.A(net2239),
    .B(net3499),
    .Y(_08053_));
 sky130_fd_sc_hd__nor2_1 _15986_ (.A(net2712),
    .B(net4076),
    .Y(_08054_));
 sky130_fd_sc_hd__a31oi_1 _15987_ (.A1(net2712),
    .A2(net4071),
    .A3(_08053_),
    .B1(_08054_),
    .Y(_08055_));
 sky130_fd_sc_hd__nor2_1 _15988_ (.A(net3449),
    .B(_07838_),
    .Y(_08056_));
 sky130_fd_sc_hd__nand3_1 _15989_ (.A(net2712),
    .B(net3394),
    .C(_08053_),
    .Y(_08057_));
 sky130_fd_sc_hd__o221a_1 _15990_ (.A1(net4068),
    .A2(_08055_),
    .B1(_08056_),
    .B2(_08053_),
    .C1(_08057_),
    .X(_08058_));
 sky130_fd_sc_hd__xnor2_1 _15991_ (.A(_08052_),
    .B(net1258),
    .Y(_08059_));
 sky130_fd_sc_hd__xor2_1 _15992_ (.A(_08049_),
    .B(_08059_),
    .X(_08060_));
 sky130_fd_sc_hd__and2_1 _15993_ (.A(_08037_),
    .B(net883),
    .X(_08061_));
 sky130_fd_sc_hd__or2_1 _15994_ (.A(_08037_),
    .B(net883),
    .X(_08062_));
 sky130_fd_sc_hd__and2b_1 _15995_ (.A_N(_08061_),
    .B(_08062_),
    .X(_08063_));
 sky130_fd_sc_hd__xnor2_1 _15996_ (.A(_08018_),
    .B(_08063_),
    .Y(_08064_));
 sky130_fd_sc_hd__and2_1 _15997_ (.A(net884),
    .B(_07983_),
    .X(_08065_));
 sky130_fd_sc_hd__o21a_1 _15998_ (.A1(net826),
    .A2(_08065_),
    .B1(_07984_),
    .X(_08066_));
 sky130_fd_sc_hd__o21a_1 _15999_ (.A1(_07979_),
    .A2(net1094),
    .B1(_07977_),
    .X(_08067_));
 sky130_fd_sc_hd__a21o_1 _16000_ (.A1(_07979_),
    .A2(net1094),
    .B1(_08067_),
    .X(_08068_));
 sky130_fd_sc_hd__o32a_1 _16001_ (.A1(net3459),
    .A2(net2803),
    .A3(_07900_),
    .B1(net2224),
    .B2(net2829),
    .X(_08069_));
 sky130_fd_sc_hd__and4_1 _16002_ (.A(net3546),
    .B(net2846),
    .C(net2732),
    .D(net1846),
    .X(_08070_));
 sky130_fd_sc_hd__a21oi_1 _16003_ (.A1(_07973_),
    .A2(_08069_),
    .B1(_08070_),
    .Y(_08071_));
 sky130_fd_sc_hd__xnor2_1 _16004_ (.A(net1521),
    .B(net1257),
    .Y(_08072_));
 sky130_fd_sc_hd__xnor2_2 _16005_ (.A(_08068_),
    .B(_08072_),
    .Y(_08073_));
 sky130_fd_sc_hd__xnor2_1 _16006_ (.A(_08066_),
    .B(_08073_),
    .Y(_08074_));
 sky130_fd_sc_hd__xnor2_1 _16007_ (.A(_08064_),
    .B(_08074_),
    .Y(_08075_));
 sky130_fd_sc_hd__xnor2_1 _16008_ (.A(_08016_),
    .B(net673),
    .Y(_08076_));
 sky130_fd_sc_hd__xnor2_1 _16009_ (.A(_08014_),
    .B(_08076_),
    .Y(_08077_));
 sky130_fd_sc_hd__or2b_1 _16010_ (.A(_08001_),
    .B_N(_07999_),
    .X(_08078_));
 sky130_fd_sc_hd__and2b_1 _16011_ (.A_N(_07999_),
    .B(_08001_),
    .X(_08079_));
 sky130_fd_sc_hd__a21oi_1 _16012_ (.A1(_07997_),
    .A2(_08078_),
    .B1(_08079_),
    .Y(_08080_));
 sky130_fd_sc_hd__nand2_1 _16013_ (.A(_08077_),
    .B(_08080_),
    .Y(_08081_));
 sky130_fd_sc_hd__or2_1 _16014_ (.A(_08077_),
    .B(_08080_),
    .X(_08082_));
 sky130_fd_sc_hd__nand2_1 _16015_ (.A(_08081_),
    .B(_08082_),
    .Y(_08083_));
 sky130_fd_sc_hd__inv_2 _16016_ (.A(_08007_),
    .Y(_08084_));
 sky130_fd_sc_hd__a21o_1 _16017_ (.A1(net425),
    .A2(_08084_),
    .B1(_08008_),
    .X(_08085_));
 sky130_fd_sc_hd__xnor2_1 _16018_ (.A(_08083_),
    .B(_08085_),
    .Y(_08086_));
 sky130_fd_sc_hd__mux2_1 _16019_ (.A0(\matmul0.matmul_stage_inst.mult1[6] ),
    .A1(net359),
    .S(net2679),
    .X(_08087_));
 sky130_fd_sc_hd__clkbuf_1 _16020_ (.A(_08087_),
    .X(_00221_));
 sky130_fd_sc_hd__or2b_1 _16021_ (.A(_08008_),
    .B_N(_08082_),
    .X(_08088_));
 sky130_fd_sc_hd__nand2_1 _16022_ (.A(_08007_),
    .B(_08082_),
    .Y(_08089_));
 sky130_fd_sc_hd__o211ai_1 _16023_ (.A1(net425),
    .A2(_08088_),
    .B1(_08089_),
    .C1(_08081_),
    .Y(_08090_));
 sky130_fd_sc_hd__or2_1 _16024_ (.A(_08016_),
    .B(net673),
    .X(_08091_));
 sky130_fd_sc_hd__and2_1 _16025_ (.A(_08016_),
    .B(net673),
    .X(_08092_));
 sky130_fd_sc_hd__a21oi_1 _16026_ (.A1(_08014_),
    .A2(_08091_),
    .B1(_08092_),
    .Y(_08093_));
 sky130_fd_sc_hd__nor2_1 _16027_ (.A(net2708),
    .B(net3400),
    .Y(_08094_));
 sky130_fd_sc_hd__nor2_1 _16028_ (.A(net2649),
    .B(net2624),
    .Y(_08095_));
 sky130_fd_sc_hd__nor2_1 _16029_ (.A(net2722),
    .B(net3417),
    .Y(_08096_));
 sky130_fd_sc_hd__xnor2_1 _16030_ (.A(_08095_),
    .B(_08096_),
    .Y(_08097_));
 sky130_fd_sc_hd__xnor2_2 _16031_ (.A(_08094_),
    .B(_08097_),
    .Y(_08098_));
 sky130_fd_sc_hd__o21ai_1 _16032_ (.A1(net2239),
    .A2(_08056_),
    .B1(net2812),
    .Y(_08099_));
 sky130_fd_sc_hd__nand2_1 _16033_ (.A(net2239),
    .B(_08056_),
    .Y(_08100_));
 sky130_fd_sc_hd__a21oi_1 _16034_ (.A1(_08099_),
    .A2(_08100_),
    .B1(_07932_),
    .Y(_08101_));
 sky130_fd_sc_hd__a21o_1 _16035_ (.A1(_08038_),
    .A2(_08039_),
    .B1(_08041_),
    .X(_08102_));
 sky130_fd_sc_hd__o21a_1 _16036_ (.A1(_08038_),
    .A2(_08039_),
    .B1(_08102_),
    .X(_08103_));
 sky130_fd_sc_hd__xor2_1 _16037_ (.A(net1516),
    .B(_08103_),
    .X(_08104_));
 sky130_fd_sc_hd__xnor2_2 _16038_ (.A(_08098_),
    .B(_08104_),
    .Y(_08105_));
 sky130_fd_sc_hd__xnor2_1 _16039_ (.A(net2712),
    .B(_08053_),
    .Y(_08106_));
 sky130_fd_sc_hd__a21o_1 _16040_ (.A1(_07929_),
    .A2(net1260),
    .B1(net2700),
    .X(_08107_));
 sky130_fd_sc_hd__o21a_1 _16041_ (.A1(_07841_),
    .A2(net1260),
    .B1(_08107_),
    .X(_08108_));
 sky130_fd_sc_hd__xor2_1 _16042_ (.A(net1515),
    .B(_08108_),
    .X(_08109_));
 sky130_fd_sc_hd__nand2_1 _16043_ (.A(net2640),
    .B(_08109_),
    .Y(_08110_));
 sky130_fd_sc_hd__xnor2_1 _16044_ (.A(_08105_),
    .B(_08110_),
    .Y(_08111_));
 sky130_fd_sc_hd__a21bo_1 _16045_ (.A1(net1518),
    .A2(_08047_),
    .B1_N(net1520),
    .X(_08112_));
 sky130_fd_sc_hd__o21a_1 _16046_ (.A1(net1518),
    .A2(_08047_),
    .B1(_08112_),
    .X(_08113_));
 sky130_fd_sc_hd__nor2_2 _16047_ (.A(net2646),
    .B(net2633),
    .Y(_08114_));
 sky130_fd_sc_hd__nor2_1 _16048_ (.A(net2802),
    .B(net2660),
    .Y(_08115_));
 sky130_fd_sc_hd__nor2_1 _16049_ (.A(net2692),
    .B(net2637),
    .Y(_08116_));
 sky130_fd_sc_hd__xnor2_1 _16050_ (.A(_08115_),
    .B(_08116_),
    .Y(_08117_));
 sky130_fd_sc_hd__xnor2_1 _16051_ (.A(_08114_),
    .B(_08117_),
    .Y(_08118_));
 sky130_fd_sc_hd__a21o_1 _16052_ (.A1(_08019_),
    .A2(_08020_),
    .B1(_08021_),
    .X(_08119_));
 sky130_fd_sc_hd__o21a_1 _16053_ (.A1(_08019_),
    .A2(_08020_),
    .B1(_08119_),
    .X(_08120_));
 sky130_fd_sc_hd__nor2_2 _16054_ (.A(net2652),
    .B(net2764),
    .Y(_08121_));
 sky130_fd_sc_hd__nor2_1 _16055_ (.A(net2747),
    .B(net2656),
    .Y(_08122_));
 sky130_fd_sc_hd__nor2_1 _16056_ (.A(net2753),
    .B(net2627),
    .Y(_08123_));
 sky130_fd_sc_hd__xnor2_1 _16057_ (.A(_08122_),
    .B(_08123_),
    .Y(_08124_));
 sky130_fd_sc_hd__xnor2_2 _16058_ (.A(_08121_),
    .B(_08124_),
    .Y(_08125_));
 sky130_fd_sc_hd__xnor2_1 _16059_ (.A(_08120_),
    .B(_08125_),
    .Y(_08126_));
 sky130_fd_sc_hd__xnor2_1 _16060_ (.A(_08118_),
    .B(_08126_),
    .Y(_08127_));
 sky130_fd_sc_hd__a21o_1 _16061_ (.A1(_08025_),
    .A2(_08030_),
    .B1(_08023_),
    .X(_08128_));
 sky130_fd_sc_hd__o21a_1 _16062_ (.A1(_08025_),
    .A2(_08030_),
    .B1(_08128_),
    .X(_08129_));
 sky130_fd_sc_hd__xor2_1 _16063_ (.A(_08127_),
    .B(net1092),
    .X(_08130_));
 sky130_fd_sc_hd__xnor2_1 _16064_ (.A(net1093),
    .B(_08130_),
    .Y(_08131_));
 sky130_fd_sc_hd__or2_1 _16065_ (.A(net2205),
    .B(_08049_),
    .X(_08132_));
 sky130_fd_sc_hd__nor2_1 _16066_ (.A(net1525),
    .B(net1258),
    .Y(_08133_));
 sky130_fd_sc_hd__and2_1 _16067_ (.A(net2205),
    .B(net1258),
    .X(_08134_));
 sky130_fd_sc_hd__o21a_1 _16068_ (.A1(_08050_),
    .A2(_08134_),
    .B1(_08049_),
    .X(_08135_));
 sky130_fd_sc_hd__a221o_1 _16069_ (.A1(_08050_),
    .A2(net1258),
    .B1(_08132_),
    .B2(_08133_),
    .C1(_08135_),
    .X(_08136_));
 sky130_fd_sc_hd__xor2_1 _16070_ (.A(_08131_),
    .B(_08136_),
    .X(_08137_));
 sky130_fd_sc_hd__xnor2_2 _16071_ (.A(net776),
    .B(_08137_),
    .Y(_08138_));
 sky130_fd_sc_hd__a21bo_1 _16072_ (.A1(_08034_),
    .A2(net1261),
    .B1_N(_08032_),
    .X(_08139_));
 sky130_fd_sc_hd__o21a_1 _16073_ (.A1(_08034_),
    .A2(net1261),
    .B1(_08139_),
    .X(_08140_));
 sky130_fd_sc_hd__o21ai_1 _16074_ (.A1(net2662),
    .A2(_08028_),
    .B1(_08026_),
    .Y(_08141_));
 sky130_fd_sc_hd__nand2_1 _16075_ (.A(net2662),
    .B(_08028_),
    .Y(_08142_));
 sky130_fd_sc_hd__a21oi_1 _16076_ (.A1(_08141_),
    .A2(_08142_),
    .B1(net3460),
    .Y(_08143_));
 sky130_fd_sc_hd__a211oi_1 _16077_ (.A1(_08026_),
    .A2(_08028_),
    .B1(net2846),
    .C1(net2224),
    .Y(_08144_));
 sky130_fd_sc_hd__a311o_1 _16078_ (.A1(net2224),
    .A2(_08026_),
    .A3(_08028_),
    .B1(_08143_),
    .C1(_08144_),
    .X(_08145_));
 sky130_fd_sc_hd__xor2_1 _16079_ (.A(net1517),
    .B(net1256),
    .X(_08146_));
 sky130_fd_sc_hd__xnor2_2 _16080_ (.A(_08140_),
    .B(_08146_),
    .Y(_08147_));
 sky130_fd_sc_hd__a21o_1 _16081_ (.A1(_08018_),
    .A2(_08062_),
    .B1(_08061_),
    .X(_08148_));
 sky130_fd_sc_hd__xnor2_1 _16082_ (.A(_08147_),
    .B(_08148_),
    .Y(_08149_));
 sky130_fd_sc_hd__xor2_2 _16083_ (.A(_08138_),
    .B(_08149_),
    .X(_08150_));
 sky130_fd_sc_hd__nand2_1 _16084_ (.A(_08066_),
    .B(_08073_),
    .Y(_08151_));
 sky130_fd_sc_hd__nor2_1 _16085_ (.A(_08066_),
    .B(_08073_),
    .Y(_08152_));
 sky130_fd_sc_hd__a21o_1 _16086_ (.A1(_08064_),
    .A2(_08151_),
    .B1(_08152_),
    .X(_08153_));
 sky130_fd_sc_hd__a21o_1 _16087_ (.A1(_08068_),
    .A2(net1257),
    .B1(net1521),
    .X(_08154_));
 sky130_fd_sc_hd__o21a_1 _16088_ (.A1(_08068_),
    .A2(net1257),
    .B1(_08154_),
    .X(_08155_));
 sky130_fd_sc_hd__xor2_1 _16089_ (.A(_08153_),
    .B(_08155_),
    .X(_08156_));
 sky130_fd_sc_hd__xnor2_1 _16090_ (.A(_08150_),
    .B(_08156_),
    .Y(_08157_));
 sky130_fd_sc_hd__and2_1 _16091_ (.A(net572),
    .B(_08157_),
    .X(_08158_));
 sky130_fd_sc_hd__nor2_1 _16092_ (.A(net572),
    .B(_08157_),
    .Y(_08159_));
 sky130_fd_sc_hd__nor2_1 _16093_ (.A(_08158_),
    .B(_08159_),
    .Y(_08160_));
 sky130_fd_sc_hd__xnor2_1 _16094_ (.A(net385),
    .B(net493),
    .Y(_08161_));
 sky130_fd_sc_hd__mux2_1 _16095_ (.A0(\matmul0.matmul_stage_inst.mult1[7] ),
    .A1(net354),
    .S(net2679),
    .X(_08162_));
 sky130_fd_sc_hd__clkbuf_1 _16096_ (.A(_08162_),
    .X(_00222_));
 sky130_fd_sc_hd__a21o_1 _16097_ (.A1(net2699),
    .A2(net2727),
    .B1(net1260),
    .X(_08163_));
 sky130_fd_sc_hd__and2b_1 _16098_ (.A_N(_07841_),
    .B(net1260),
    .X(_08164_));
 sky130_fd_sc_hd__a21oi_2 _16099_ (.A1(net2234),
    .A2(_08163_),
    .B1(_08164_),
    .Y(_08165_));
 sky130_fd_sc_hd__o21ai_1 _16100_ (.A1(net2630),
    .A2(_08165_),
    .B1(_08105_),
    .Y(_08166_));
 sky130_fd_sc_hd__a211o_1 _16101_ (.A1(_08105_),
    .A2(_08165_),
    .B1(net1515),
    .C1(net1526),
    .X(_08167_));
 sky130_fd_sc_hd__o21ai_1 _16102_ (.A1(_08105_),
    .A2(_08165_),
    .B1(_08167_),
    .Y(_08168_));
 sky130_fd_sc_hd__a32o_1 _16103_ (.A1(net1526),
    .A2(net1515),
    .A3(_08166_),
    .B1(_08168_),
    .B2(net2640),
    .X(_08169_));
 sky130_fd_sc_hd__nor2_2 _16104_ (.A(net2648),
    .B(net3418),
    .Y(_08170_));
 sky130_fd_sc_hd__o2bb2a_1 _16105_ (.A1_N(net3561),
    .A2_N(_07684_),
    .B1(net4075),
    .B2(net2840),
    .X(_08171_));
 sky130_fd_sc_hd__nor2_1 _16106_ (.A(net2707),
    .B(_07932_),
    .Y(_08172_));
 sky130_fd_sc_hd__nand2_1 _16107_ (.A(net3561),
    .B(net3394),
    .Y(_08173_));
 sky130_fd_sc_hd__o221a_1 _16108_ (.A1(net4074),
    .A2(_08171_),
    .B1(_08172_),
    .B2(net2816),
    .C1(_08173_),
    .X(_08174_));
 sky130_fd_sc_hd__xnor2_1 _16109_ (.A(_08170_),
    .B(_08174_),
    .Y(_08175_));
 sky130_fd_sc_hd__a21o_1 _16110_ (.A1(_08094_),
    .A2(_08095_),
    .B1(_08096_),
    .X(_08176_));
 sky130_fd_sc_hd__o21a_1 _16111_ (.A1(_08094_),
    .A2(_08095_),
    .B1(_08176_),
    .X(_08177_));
 sky130_fd_sc_hd__a21o_1 _16112_ (.A1(net3449),
    .A2(net2719),
    .B1(net3499),
    .X(_08178_));
 sky130_fd_sc_hd__nand2_1 _16113_ (.A(net2712),
    .B(net2239),
    .Y(_08179_));
 sky130_fd_sc_hd__a21oi_1 _16114_ (.A1(_08178_),
    .A2(_08179_),
    .B1(_07932_),
    .Y(_08180_));
 sky130_fd_sc_hd__xnor2_1 _16115_ (.A(_08177_),
    .B(_08180_),
    .Y(_08181_));
 sky130_fd_sc_hd__xnor2_1 _16116_ (.A(net1512),
    .B(_08181_),
    .Y(_08182_));
 sky130_fd_sc_hd__a31o_1 _16117_ (.A1(net2700),
    .A2(_07841_),
    .A3(net1515),
    .B1(net2630),
    .X(_08183_));
 sky130_fd_sc_hd__nor2_1 _16118_ (.A(net2206),
    .B(net1513),
    .Y(_08184_));
 sky130_fd_sc_hd__nor2_2 _16119_ (.A(net1254),
    .B(net1253),
    .Y(_08185_));
 sky130_fd_sc_hd__xnor2_1 _16120_ (.A(net1091),
    .B(_08185_),
    .Y(_08186_));
 sky130_fd_sc_hd__nor2_1 _16121_ (.A(net2752),
    .B(net3435),
    .Y(_08187_));
 sky130_fd_sc_hd__nor2_1 _16122_ (.A(net3484),
    .B(net3599),
    .Y(_08188_));
 sky130_fd_sc_hd__nor2_1 _16123_ (.A(net2656),
    .B(net2764),
    .Y(_08189_));
 sky130_fd_sc_hd__xnor2_1 _16124_ (.A(_08188_),
    .B(_08189_),
    .Y(_08190_));
 sky130_fd_sc_hd__xnor2_1 _16125_ (.A(_08187_),
    .B(_08190_),
    .Y(_08191_));
 sky130_fd_sc_hd__a21o_1 _16126_ (.A1(_08121_),
    .A2(_08122_),
    .B1(_08123_),
    .X(_08192_));
 sky130_fd_sc_hd__o21a_1 _16127_ (.A1(_08121_),
    .A2(_08122_),
    .B1(_08192_),
    .X(_08193_));
 sky130_fd_sc_hd__a211o_1 _16128_ (.A1(net3492),
    .A2(net2697),
    .B1(net3442),
    .C1(net3516),
    .X(_08194_));
 sky130_fd_sc_hd__a211o_1 _16129_ (.A1(net3522),
    .A2(net3424),
    .B1(net3429),
    .C1(net3533),
    .X(_08195_));
 sky130_fd_sc_hd__a211o_1 _16130_ (.A1(_08194_),
    .A2(_08195_),
    .B1(net2645),
    .C1(net2659),
    .X(_08196_));
 sky130_fd_sc_hd__o211ai_1 _16131_ (.A1(net2645),
    .A2(net2659),
    .B1(_08194_),
    .C1(_08195_),
    .Y(_08197_));
 sky130_fd_sc_hd__and2_1 _16132_ (.A(_08196_),
    .B(_08197_),
    .X(_08198_));
 sky130_fd_sc_hd__xnor2_1 _16133_ (.A(_08193_),
    .B(_08198_),
    .Y(_08199_));
 sky130_fd_sc_hd__xnor2_1 _16134_ (.A(_08191_),
    .B(_08199_),
    .Y(_08200_));
 sky130_fd_sc_hd__a21o_1 _16135_ (.A1(net1516),
    .A2(_08103_),
    .B1(_08098_),
    .X(_08201_));
 sky130_fd_sc_hd__o21a_1 _16136_ (.A1(net1516),
    .A2(_08103_),
    .B1(_08201_),
    .X(_08202_));
 sky130_fd_sc_hd__a21o_1 _16137_ (.A1(_08120_),
    .A2(_08125_),
    .B1(_08118_),
    .X(_08203_));
 sky130_fd_sc_hd__o21a_1 _16138_ (.A1(_08120_),
    .A2(_08125_),
    .B1(_08203_),
    .X(_08204_));
 sky130_fd_sc_hd__xnor2_1 _16139_ (.A(net1089),
    .B(net983),
    .Y(_08205_));
 sky130_fd_sc_hd__xnor2_1 _16140_ (.A(_08200_),
    .B(_08205_),
    .Y(_08206_));
 sky130_fd_sc_hd__or2_1 _16141_ (.A(_08186_),
    .B(_08206_),
    .X(_08207_));
 sky130_fd_sc_hd__nand2_1 _16142_ (.A(_08186_),
    .B(_08206_),
    .Y(_08208_));
 sky130_fd_sc_hd__nand2_1 _16143_ (.A(_08207_),
    .B(_08208_),
    .Y(_08209_));
 sky130_fd_sc_hd__xnor2_1 _16144_ (.A(net774),
    .B(_08209_),
    .Y(_08210_));
 sky130_fd_sc_hd__o21a_1 _16145_ (.A1(_08131_),
    .A2(_08136_),
    .B1(net776),
    .X(_08211_));
 sky130_fd_sc_hd__a21oi_1 _16146_ (.A1(_08131_),
    .A2(_08136_),
    .B1(_08211_),
    .Y(_08212_));
 sky130_fd_sc_hd__o21a_1 _16147_ (.A1(net1093),
    .A2(net1092),
    .B1(_08127_),
    .X(_08213_));
 sky130_fd_sc_hd__a21oi_2 _16148_ (.A1(net1093),
    .A2(net1092),
    .B1(_08213_),
    .Y(_08214_));
 sky130_fd_sc_hd__o21a_1 _16149_ (.A1(net2662),
    .A2(_08114_),
    .B1(_08116_),
    .X(_08215_));
 sky130_fd_sc_hd__a21oi_1 _16150_ (.A1(net2662),
    .A2(_08114_),
    .B1(_08215_),
    .Y(_08216_));
 sky130_fd_sc_hd__nor2_1 _16151_ (.A(net2802),
    .B(_08216_),
    .Y(_08217_));
 sky130_fd_sc_hd__a211oi_1 _16152_ (.A1(_08114_),
    .A2(_08116_),
    .B1(net2733),
    .C1(net2223),
    .Y(_08218_));
 sky130_fd_sc_hd__a311o_1 _16153_ (.A1(net2223),
    .A2(_08114_),
    .A3(_08116_),
    .B1(_08217_),
    .C1(_08218_),
    .X(_08219_));
 sky130_fd_sc_hd__and4_1 _16154_ (.A(net3459),
    .B(net2733),
    .C(net3409),
    .D(net1849),
    .X(_08220_));
 sky130_fd_sc_hd__xor2_1 _16155_ (.A(net1088),
    .B(net1511),
    .X(_08221_));
 sky130_fd_sc_hd__xnor2_2 _16156_ (.A(_08214_),
    .B(_08221_),
    .Y(_08222_));
 sky130_fd_sc_hd__xor2_1 _16157_ (.A(_08212_),
    .B(_08222_),
    .X(_08223_));
 sky130_fd_sc_hd__xor2_1 _16158_ (.A(net672),
    .B(_08223_),
    .X(_08224_));
 sky130_fd_sc_hd__a21o_1 _16159_ (.A1(_08140_),
    .A2(net1256),
    .B1(net1517),
    .X(_08225_));
 sky130_fd_sc_hd__o21a_1 _16160_ (.A1(_08140_),
    .A2(net1256),
    .B1(_08225_),
    .X(_08226_));
 sky130_fd_sc_hd__nor2_1 _16161_ (.A(_08138_),
    .B(_08148_),
    .Y(_08227_));
 sky130_fd_sc_hd__nand2_1 _16162_ (.A(_08138_),
    .B(_08148_),
    .Y(_08228_));
 sky130_fd_sc_hd__o21ai_2 _16163_ (.A1(_08147_),
    .A2(_08227_),
    .B1(_08228_),
    .Y(_08229_));
 sky130_fd_sc_hd__xor2_1 _16164_ (.A(_08226_),
    .B(_08229_),
    .X(_08230_));
 sky130_fd_sc_hd__xnor2_1 _16165_ (.A(_08224_),
    .B(_08230_),
    .Y(_08231_));
 sky130_fd_sc_hd__a21bo_1 _16166_ (.A1(_08150_),
    .A2(_08155_),
    .B1_N(_08153_),
    .X(_08232_));
 sky130_fd_sc_hd__o21ai_2 _16167_ (.A1(_08150_),
    .A2(_08155_),
    .B1(_08232_),
    .Y(_08233_));
 sky130_fd_sc_hd__xor2_1 _16168_ (.A(_08231_),
    .B(_08233_),
    .X(_08234_));
 sky130_fd_sc_hd__o21ba_1 _16169_ (.A1(net386),
    .A2(_08159_),
    .B1_N(_08158_),
    .X(_08235_));
 sky130_fd_sc_hd__xnor2_1 _16170_ (.A(_08234_),
    .B(_08235_),
    .Y(_08236_));
 sky130_fd_sc_hd__mux2_1 _16171_ (.A0(\matmul0.matmul_stage_inst.mult1[8] ),
    .A1(net311),
    .S(net2681),
    .X(_08237_));
 sky130_fd_sc_hd__clkbuf_1 _16172_ (.A(_08237_),
    .X(_00223_));
 sky130_fd_sc_hd__nand2_1 _16173_ (.A(net493),
    .B(net492),
    .Y(_08238_));
 sky130_fd_sc_hd__o2bb2a_1 _16174_ (.A1_N(net572),
    .A2_N(_08157_),
    .B1(_08231_),
    .B2(_08233_),
    .X(_08239_));
 sky130_fd_sc_hd__a21o_1 _16175_ (.A1(_08231_),
    .A2(_08233_),
    .B1(_08239_),
    .X(_08240_));
 sky130_fd_sc_hd__o21a_1 _16176_ (.A1(net385),
    .A2(_08238_),
    .B1(net424),
    .X(_08241_));
 sky130_fd_sc_hd__a21o_1 _16177_ (.A1(_08226_),
    .A2(_08229_),
    .B1(_08224_),
    .X(_08242_));
 sky130_fd_sc_hd__o21a_1 _16178_ (.A1(_08226_),
    .A2(_08229_),
    .B1(_08242_),
    .X(_08243_));
 sky130_fd_sc_hd__a21o_1 _16179_ (.A1(net672),
    .A2(_08222_),
    .B1(_08212_),
    .X(_08244_));
 sky130_fd_sc_hd__o21ai_2 _16180_ (.A1(net672),
    .A2(_08222_),
    .B1(_08244_),
    .Y(_08245_));
 sky130_fd_sc_hd__and2_1 _16181_ (.A(_08186_),
    .B(_08206_),
    .X(_08246_));
 sky130_fd_sc_hd__o21ai_4 _16182_ (.A1(net774),
    .A2(_08246_),
    .B1(_08207_),
    .Y(_08247_));
 sky130_fd_sc_hd__a21o_1 _16183_ (.A1(net1089),
    .A2(net983),
    .B1(_08200_),
    .X(_08248_));
 sky130_fd_sc_hd__o21a_1 _16184_ (.A1(net1089),
    .A2(net983),
    .B1(_08248_),
    .X(_08249_));
 sky130_fd_sc_hd__o32a_1 _16185_ (.A1(net2692),
    .A2(net2651),
    .A3(net2214),
    .B1(net2222),
    .B2(net3409),
    .X(_08250_));
 sky130_fd_sc_hd__and4_1 _16186_ (.A(net3492),
    .B(net2645),
    .C(net3522),
    .D(net1849),
    .X(_08251_));
 sky130_fd_sc_hd__a21oi_1 _16187_ (.A1(_08196_),
    .A2(_08250_),
    .B1(_08251_),
    .Y(_08252_));
 sky130_fd_sc_hd__nand2_1 _16188_ (.A(net2211),
    .B(net2215),
    .Y(_08253_));
 sky130_fd_sc_hd__or4_1 _16189_ (.A(net2691),
    .B(net2731),
    .C(net2645),
    .D(_08253_),
    .X(_08254_));
 sky130_fd_sc_hd__xnor2_1 _16190_ (.A(net1251),
    .B(net1508),
    .Y(_08255_));
 sky130_fd_sc_hd__xnor2_2 _16191_ (.A(_08249_),
    .B(_08255_),
    .Y(_08256_));
 sky130_fd_sc_hd__xnor2_1 _16192_ (.A(net2721),
    .B(net2707),
    .Y(_08257_));
 sky130_fd_sc_hd__buf_1 _16193_ (.A(net2670),
    .X(_08258_));
 sky130_fd_sc_hd__o211a_1 _16194_ (.A1(_07932_),
    .A2(_08257_),
    .B1(net2682),
    .C1(_08258_),
    .X(_08259_));
 sky130_fd_sc_hd__a211o_1 _16195_ (.A1(net2682),
    .A2(net2670),
    .B1(_07932_),
    .C1(_08257_),
    .X(_08260_));
 sky130_fd_sc_hd__and2b_1 _16196_ (.A_N(_08259_),
    .B(_08260_),
    .X(_08261_));
 sky130_fd_sc_hd__buf_1 _16197_ (.A(_08180_),
    .X(_08262_));
 sky130_fd_sc_hd__a22o_1 _16198_ (.A1(net2840),
    .A2(net3394),
    .B1(_08170_),
    .B2(net2670),
    .X(_08263_));
 sky130_fd_sc_hd__a22oi_4 _16199_ (.A1(_08170_),
    .A2(_08172_),
    .B1(_08263_),
    .B2(net2815),
    .Y(_08264_));
 sky130_fd_sc_hd__xnor2_1 _16200_ (.A(net1250),
    .B(_08264_),
    .Y(_08265_));
 sky130_fd_sc_hd__xnor2_1 _16201_ (.A(_08261_),
    .B(_08265_),
    .Y(_08266_));
 sky130_fd_sc_hd__xor2_2 _16202_ (.A(_08185_),
    .B(net981),
    .X(_08267_));
 sky130_fd_sc_hd__a21bo_1 _16203_ (.A1(_08177_),
    .A2(_08262_),
    .B1_N(net1512),
    .X(_08268_));
 sky130_fd_sc_hd__o21ai_1 _16204_ (.A1(_08177_),
    .A2(_08262_),
    .B1(_08268_),
    .Y(_08269_));
 sky130_fd_sc_hd__nor2_1 _16205_ (.A(net2752),
    .B(net3416),
    .Y(_08270_));
 sky130_fd_sc_hd__nand2_1 _16206_ (.A(net3431),
    .B(net2786),
    .Y(_08271_));
 sky130_fd_sc_hd__nor2_1 _16207_ (.A(net2746),
    .B(net3435),
    .Y(_08272_));
 sky130_fd_sc_hd__xnor2_1 _16208_ (.A(_08271_),
    .B(_08272_),
    .Y(_08273_));
 sky130_fd_sc_hd__xnor2_1 _16209_ (.A(_08270_),
    .B(_08273_),
    .Y(_08274_));
 sky130_fd_sc_hd__a21o_1 _16210_ (.A1(_08187_),
    .A2(_08188_),
    .B1(_08189_),
    .X(_08275_));
 sky130_fd_sc_hd__o21a_1 _16211_ (.A1(_08187_),
    .A2(_08188_),
    .B1(_08275_),
    .X(_08276_));
 sky130_fd_sc_hd__o211a_1 _16212_ (.A1(net3516),
    .A2(net3429),
    .B1(net3424),
    .C1(net3587),
    .X(_08277_));
 sky130_fd_sc_hd__o211a_1 _16213_ (.A1(net2655),
    .A2(net3442),
    .B1(net2697),
    .C1(net3522),
    .X(_08278_));
 sky130_fd_sc_hd__nor2_1 _16214_ (.A(_08277_),
    .B(_08278_),
    .Y(_08279_));
 sky130_fd_sc_hd__nor2_1 _16215_ (.A(net2691),
    .B(net2659),
    .Y(_08280_));
 sky130_fd_sc_hd__xnor2_2 _16216_ (.A(_08279_),
    .B(_08280_),
    .Y(_08281_));
 sky130_fd_sc_hd__xor2_1 _16217_ (.A(_08276_),
    .B(_08281_),
    .X(_08282_));
 sky130_fd_sc_hd__xnor2_1 _16218_ (.A(_08274_),
    .B(_08282_),
    .Y(_08283_));
 sky130_fd_sc_hd__a21o_1 _16219_ (.A1(_08193_),
    .A2(_08198_),
    .B1(_08191_),
    .X(_08284_));
 sky130_fd_sc_hd__o21a_1 _16220_ (.A1(_08193_),
    .A2(_08198_),
    .B1(_08284_),
    .X(_08285_));
 sky130_fd_sc_hd__nor2_1 _16221_ (.A(_08283_),
    .B(_08285_),
    .Y(_08286_));
 sky130_fd_sc_hd__nand2_1 _16222_ (.A(_08283_),
    .B(_08285_),
    .Y(_08287_));
 sky130_fd_sc_hd__or2b_1 _16223_ (.A(_08286_),
    .B_N(_08287_),
    .X(_08288_));
 sky130_fd_sc_hd__xnor2_1 _16224_ (.A(net979),
    .B(_08288_),
    .Y(_08289_));
 sky130_fd_sc_hd__buf_1 _16225_ (.A(net1254),
    .X(_08290_));
 sky130_fd_sc_hd__or2_1 _16226_ (.A(net2206),
    .B(net1513),
    .X(_08291_));
 sky130_fd_sc_hd__clkbuf_1 _16227_ (.A(_08291_),
    .X(_08292_));
 sky130_fd_sc_hd__o21ai_2 _16228_ (.A1(net1091),
    .A2(_08290_),
    .B1(net1085),
    .Y(_08293_));
 sky130_fd_sc_hd__xnor2_1 _16229_ (.A(_08289_),
    .B(_08293_),
    .Y(_08294_));
 sky130_fd_sc_hd__xnor2_2 _16230_ (.A(_08267_),
    .B(_08294_),
    .Y(_08295_));
 sky130_fd_sc_hd__xor2_2 _16231_ (.A(_08256_),
    .B(_08295_),
    .X(_08296_));
 sky130_fd_sc_hd__xnor2_4 _16232_ (.A(_08247_),
    .B(_08296_),
    .Y(_08297_));
 sky130_fd_sc_hd__a21bo_1 _16233_ (.A1(net1088),
    .A2(net1511),
    .B1_N(_08214_),
    .X(_08298_));
 sky130_fd_sc_hd__o21a_2 _16234_ (.A1(net1088),
    .A2(net1511),
    .B1(_08298_),
    .X(_08299_));
 sky130_fd_sc_hd__xor2_1 _16235_ (.A(_08297_),
    .B(_08299_),
    .X(_08300_));
 sky130_fd_sc_hd__xnor2_1 _16236_ (.A(_08245_),
    .B(_08300_),
    .Y(_08301_));
 sky130_fd_sc_hd__nand2_1 _16237_ (.A(net491),
    .B(_08301_),
    .Y(_08302_));
 sky130_fd_sc_hd__or2_1 _16238_ (.A(net491),
    .B(_08301_),
    .X(_08303_));
 sky130_fd_sc_hd__and2_1 _16239_ (.A(_08302_),
    .B(_08303_),
    .X(_08304_));
 sky130_fd_sc_hd__xnor2_1 _16240_ (.A(_08241_),
    .B(_08304_),
    .Y(_08305_));
 sky130_fd_sc_hd__mux2_1 _16241_ (.A0(\matmul0.matmul_stage_inst.mult1[9] ),
    .A1(net305),
    .S(net2681),
    .X(_08306_));
 sky130_fd_sc_hd__clkbuf_1 _16242_ (.A(_08306_),
    .X(_00224_));
 sky130_fd_sc_hd__o21a_1 _16243_ (.A1(_08256_),
    .A2(_08295_),
    .B1(_08247_),
    .X(_08307_));
 sky130_fd_sc_hd__a21o_1 _16244_ (.A1(_08256_),
    .A2(_08295_),
    .B1(_08307_),
    .X(_08308_));
 sky130_fd_sc_hd__o21ba_1 _16245_ (.A1(_08267_),
    .A2(_08293_),
    .B1_N(_08289_),
    .X(_08309_));
 sky130_fd_sc_hd__a21oi_1 _16246_ (.A1(_08267_),
    .A2(_08293_),
    .B1(_08309_),
    .Y(_08310_));
 sky130_fd_sc_hd__a21oi_2 _16247_ (.A1(net979),
    .A2(_08287_),
    .B1(_08286_),
    .Y(_08311_));
 sky130_fd_sc_hd__nand2_1 _16248_ (.A(net3587),
    .B(net2215),
    .Y(_08312_));
 sky130_fd_sc_hd__nor2_1 _16249_ (.A(net2651),
    .B(_08312_),
    .Y(_08313_));
 sky130_fd_sc_hd__xnor2_1 _16250_ (.A(net2210),
    .B(_08313_),
    .Y(_08314_));
 sky130_fd_sc_hd__o221a_1 _16251_ (.A1(net2220),
    .A2(_08279_),
    .B1(_08312_),
    .B2(net2651),
    .C1(net3492),
    .X(_08315_));
 sky130_fd_sc_hd__a21oi_1 _16252_ (.A1(net2691),
    .A2(_08314_),
    .B1(_08315_),
    .Y(_08316_));
 sky130_fd_sc_hd__xnor2_1 _16253_ (.A(net1509),
    .B(net1083),
    .Y(_08317_));
 sky130_fd_sc_hd__xnor2_2 _16254_ (.A(_08311_),
    .B(_08317_),
    .Y(_08318_));
 sky130_fd_sc_hd__nor2_2 _16255_ (.A(net2751),
    .B(net2643),
    .Y(_08319_));
 sky130_fd_sc_hd__nor2_1 _16256_ (.A(net2746),
    .B(net3415),
    .Y(_08320_));
 sky130_fd_sc_hd__nor2_1 _16257_ (.A(net2246),
    .B(_08040_),
    .Y(_08321_));
 sky130_fd_sc_hd__xnor2_1 _16258_ (.A(_08320_),
    .B(_08321_),
    .Y(_08322_));
 sky130_fd_sc_hd__xor2_2 _16259_ (.A(_08319_),
    .B(_08322_),
    .X(_08323_));
 sky130_fd_sc_hd__o21ba_1 _16260_ (.A1(_08270_),
    .A2(_08272_),
    .B1_N(_08271_),
    .X(_08324_));
 sky130_fd_sc_hd__a21o_1 _16261_ (.A1(_08270_),
    .A2(_08272_),
    .B1(_08324_),
    .X(_08325_));
 sky130_fd_sc_hd__o211a_1 _16262_ (.A1(net2655),
    .A2(net2632),
    .B1(net3424),
    .C1(net3431),
    .X(_08326_));
 sky130_fd_sc_hd__o211a_1 _16263_ (.A1(net2626),
    .A2(net2636),
    .B1(net2697),
    .C1(net3587),
    .X(_08327_));
 sky130_fd_sc_hd__nor2_1 _16264_ (.A(_08326_),
    .B(_08327_),
    .Y(_08328_));
 sky130_fd_sc_hd__or3_1 _16265_ (.A(net2651),
    .B(net2659),
    .C(_08328_),
    .X(_08329_));
 sky130_fd_sc_hd__o21ai_1 _16266_ (.A1(net2651),
    .A2(net2220),
    .B1(_08328_),
    .Y(_08330_));
 sky130_fd_sc_hd__and2_1 _16267_ (.A(_08329_),
    .B(_08330_),
    .X(_08331_));
 sky130_fd_sc_hd__xnor2_1 _16268_ (.A(_08325_),
    .B(net1249),
    .Y(_08332_));
 sky130_fd_sc_hd__xnor2_2 _16269_ (.A(_08323_),
    .B(_08332_),
    .Y(_08333_));
 sky130_fd_sc_hd__o21ba_1 _16270_ (.A1(_08264_),
    .A2(_08261_),
    .B1_N(net1250),
    .X(_08334_));
 sky130_fd_sc_hd__a21o_1 _16271_ (.A1(_08264_),
    .A2(_08261_),
    .B1(_08334_),
    .X(_08335_));
 sky130_fd_sc_hd__a21bo_1 _16272_ (.A1(_08276_),
    .A2(_08281_),
    .B1_N(_08274_),
    .X(_08336_));
 sky130_fd_sc_hd__o21ai_2 _16273_ (.A1(_08276_),
    .A2(_08281_),
    .B1(_08336_),
    .Y(_08337_));
 sky130_fd_sc_hd__xnor2_1 _16274_ (.A(net978),
    .B(_08337_),
    .Y(_08338_));
 sky130_fd_sc_hd__xnor2_2 _16275_ (.A(_08333_),
    .B(_08338_),
    .Y(_08339_));
 sky130_fd_sc_hd__and2b_1 _16276_ (.A_N(net1087),
    .B(net981),
    .X(_08340_));
 sky130_fd_sc_hd__a21oi_1 _16277_ (.A1(net2707),
    .A2(_08258_),
    .B1(net2721),
    .Y(_08341_));
 sky130_fd_sc_hd__a21o_1 _16278_ (.A1(net2840),
    .A2(net2644),
    .B1(_08341_),
    .X(_08342_));
 sky130_fd_sc_hd__a31o_1 _16279_ (.A1(net2721),
    .A2(net2707),
    .A3(net2648),
    .B1(_07932_),
    .X(_08343_));
 sky130_fd_sc_hd__a21o_1 _16280_ (.A1(net2682),
    .A2(_08342_),
    .B1(_08343_),
    .X(_08344_));
 sky130_fd_sc_hd__xnor2_1 _16281_ (.A(net1250),
    .B(_08344_),
    .Y(_08345_));
 sky130_fd_sc_hd__xor2_1 _16282_ (.A(_08185_),
    .B(net1081),
    .X(_08346_));
 sky130_fd_sc_hd__o21ai_1 _16283_ (.A1(net1253),
    .A2(_08340_),
    .B1(_08346_),
    .Y(_08347_));
 sky130_fd_sc_hd__inv_2 _16284_ (.A(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__nor3_1 _16285_ (.A(net1253),
    .B(_08346_),
    .C(_08340_),
    .Y(_08349_));
 sky130_fd_sc_hd__nor2_1 _16286_ (.A(_08348_),
    .B(_08349_),
    .Y(_08350_));
 sky130_fd_sc_hd__xnor2_2 _16287_ (.A(_08339_),
    .B(_08350_),
    .Y(_08351_));
 sky130_fd_sc_hd__xor2_1 _16288_ (.A(_08318_),
    .B(_08351_),
    .X(_08352_));
 sky130_fd_sc_hd__xnor2_1 _16289_ (.A(_08310_),
    .B(_08352_),
    .Y(_08353_));
 sky130_fd_sc_hd__a21bo_1 _16290_ (.A1(_08249_),
    .A2(net1251),
    .B1_N(net1508),
    .X(_08354_));
 sky130_fd_sc_hd__o21a_1 _16291_ (.A1(_08249_),
    .A2(net1251),
    .B1(_08354_),
    .X(_08355_));
 sky130_fd_sc_hd__nor2_1 _16292_ (.A(_08353_),
    .B(net724),
    .Y(_08356_));
 sky130_fd_sc_hd__nand2_1 _16293_ (.A(_08353_),
    .B(net724),
    .Y(_08357_));
 sky130_fd_sc_hd__and2b_1 _16294_ (.A_N(_08356_),
    .B(_08357_),
    .X(_08358_));
 sky130_fd_sc_hd__xnor2_2 _16295_ (.A(_08308_),
    .B(_08358_),
    .Y(_08359_));
 sky130_fd_sc_hd__and3_1 _16296_ (.A(net491),
    .B(_08297_),
    .C(_08299_),
    .X(_08360_));
 sky130_fd_sc_hd__nor2_1 _16297_ (.A(net491),
    .B(_08299_),
    .Y(_08361_));
 sky130_fd_sc_hd__and2b_1 _16298_ (.A_N(_08297_),
    .B(_08361_),
    .X(_08362_));
 sky130_fd_sc_hd__mux2_1 _16299_ (.A0(_08360_),
    .A1(_08362_),
    .S(_08245_),
    .X(_08363_));
 sky130_fd_sc_hd__a21oi_1 _16300_ (.A1(net491),
    .A2(_08299_),
    .B1(_08297_),
    .Y(_08364_));
 sky130_fd_sc_hd__or2_1 _16301_ (.A(_08361_),
    .B(_08364_),
    .X(_08365_));
 sky130_fd_sc_hd__o21bai_1 _16302_ (.A1(_08245_),
    .A2(_08365_),
    .B1_N(_08360_),
    .Y(_08366_));
 sky130_fd_sc_hd__a21o_1 _16303_ (.A1(_08245_),
    .A2(_08365_),
    .B1(_08362_),
    .X(_08367_));
 sky130_fd_sc_hd__mux2_1 _16304_ (.A0(_08366_),
    .A1(_08367_),
    .S(_08241_),
    .X(_08368_));
 sky130_fd_sc_hd__or2_1 _16305_ (.A(_08363_),
    .B(_08368_),
    .X(_08369_));
 sky130_fd_sc_hd__xnor2_1 _16306_ (.A(_08359_),
    .B(_08369_),
    .Y(_08370_));
 sky130_fd_sc_hd__mux2_1 _16307_ (.A0(\matmul0.matmul_stage_inst.mult1[10] ),
    .A1(net247),
    .S(net3478),
    .X(_08371_));
 sky130_fd_sc_hd__clkbuf_1 _16308_ (.A(_08371_),
    .X(_00225_));
 sky130_fd_sc_hd__a21bo_1 _16309_ (.A1(_08297_),
    .A2(_08299_),
    .B1_N(_08245_),
    .X(_08372_));
 sky130_fd_sc_hd__o21a_1 _16310_ (.A1(_08297_),
    .A2(_08299_),
    .B1(_08372_),
    .X(_08373_));
 sky130_fd_sc_hd__nand2_1 _16311_ (.A(net424),
    .B(_08302_),
    .Y(_08374_));
 sky130_fd_sc_hd__a22o_1 _16312_ (.A1(_08359_),
    .A2(_08373_),
    .B1(_08374_),
    .B2(_08303_),
    .X(_08375_));
 sky130_fd_sc_hd__and4b_1 _16313_ (.A_N(net385),
    .B(net493),
    .C(net492),
    .D(_08304_),
    .X(_08376_));
 sky130_fd_sc_hd__o22ai_1 _16314_ (.A1(_08359_),
    .A2(_08373_),
    .B1(_08375_),
    .B2(_08376_),
    .Y(_08377_));
 sky130_fd_sc_hd__a21o_1 _16315_ (.A1(_08308_),
    .A2(_08357_),
    .B1(_08356_),
    .X(_08378_));
 sky130_fd_sc_hd__a21bo_1 _16316_ (.A1(_08318_),
    .A2(_08351_),
    .B1_N(_08310_),
    .X(_08379_));
 sky130_fd_sc_hd__o21ai_1 _16317_ (.A1(_08318_),
    .A2(_08351_),
    .B1(_08379_),
    .Y(_08380_));
 sky130_fd_sc_hd__inv_2 _16318_ (.A(net571),
    .Y(_08381_));
 sky130_fd_sc_hd__mux2_1 _16319_ (.A0(net2815),
    .A1(net1250),
    .S(net2648),
    .X(_08382_));
 sky130_fd_sc_hd__a211o_1 _16320_ (.A1(net2721),
    .A2(net2707),
    .B1(net2648),
    .C1(_08258_),
    .X(_08383_));
 sky130_fd_sc_hd__o211a_1 _16321_ (.A1(net2815),
    .A2(net2682),
    .B1(net1250),
    .C1(_08383_),
    .X(_08384_));
 sky130_fd_sc_hd__a21oi_1 _16322_ (.A1(net2841),
    .A2(_08382_),
    .B1(_08384_),
    .Y(_08385_));
 sky130_fd_sc_hd__nor2_1 _16323_ (.A(net2629),
    .B(_08385_),
    .Y(_08386_));
 sky130_fd_sc_hd__nand2_1 _16324_ (.A(net2791),
    .B(net2639),
    .Y(_08387_));
 sky130_fd_sc_hd__nand2_1 _16325_ (.A(net2783),
    .B(net3402),
    .Y(_08388_));
 sky130_fd_sc_hd__nand2_1 _16326_ (.A(net2772),
    .B(net2204),
    .Y(_08389_));
 sky130_fd_sc_hd__xnor2_1 _16327_ (.A(_08388_),
    .B(_08389_),
    .Y(_08390_));
 sky130_fd_sc_hd__xor2_1 _16328_ (.A(_08387_),
    .B(_08390_),
    .X(_08391_));
 sky130_fd_sc_hd__o21a_1 _16329_ (.A1(_08319_),
    .A2(_08320_),
    .B1(_08321_),
    .X(_08392_));
 sky130_fd_sc_hd__a21o_1 _16330_ (.A1(_08319_),
    .A2(_08320_),
    .B1(_08392_),
    .X(_08393_));
 sky130_fd_sc_hd__o211a_1 _16331_ (.A1(net2626),
    .A2(net2632),
    .B1(net3424),
    .C1(net3421),
    .X(_08394_));
 sky130_fd_sc_hd__o211a_1 _16332_ (.A1(_08040_),
    .A2(net2636),
    .B1(net2697),
    .C1(net3431),
    .X(_08395_));
 sky130_fd_sc_hd__nor2_1 _16333_ (.A(_08394_),
    .B(_08395_),
    .Y(_08396_));
 sky130_fd_sc_hd__nor2_1 _16334_ (.A(net2654),
    .B(net2218),
    .Y(_08397_));
 sky130_fd_sc_hd__xnor2_1 _16335_ (.A(net1840),
    .B(_08397_),
    .Y(_08398_));
 sky130_fd_sc_hd__nand2_1 _16336_ (.A(_08393_),
    .B(_08398_),
    .Y(_08399_));
 sky130_fd_sc_hd__or2_1 _16337_ (.A(_08393_),
    .B(_08398_),
    .X(_08400_));
 sky130_fd_sc_hd__nand2_1 _16338_ (.A(_08399_),
    .B(_08400_),
    .Y(_08401_));
 sky130_fd_sc_hd__xnor2_1 _16339_ (.A(net1248),
    .B(_08401_),
    .Y(_08402_));
 sky130_fd_sc_hd__o21ba_1 _16340_ (.A1(_08325_),
    .A2(net1249),
    .B1_N(_08323_),
    .X(_08403_));
 sky130_fd_sc_hd__a21o_1 _16341_ (.A1(_08325_),
    .A2(net1249),
    .B1(_08403_),
    .X(_08404_));
 sky130_fd_sc_hd__and2_1 _16342_ (.A(_08402_),
    .B(_08404_),
    .X(_08405_));
 sky130_fd_sc_hd__or2_1 _16343_ (.A(_08402_),
    .B(_08404_),
    .X(_08406_));
 sky130_fd_sc_hd__and2b_1 _16344_ (.A_N(_08405_),
    .B(_08406_),
    .X(_08407_));
 sky130_fd_sc_hd__xnor2_2 _16345_ (.A(net882),
    .B(_08407_),
    .Y(_08408_));
 sky130_fd_sc_hd__a21oi_1 _16346_ (.A1(net2682),
    .A2(net3561),
    .B1(_08343_),
    .Y(_08409_));
 sky130_fd_sc_hd__xnor2_1 _16347_ (.A(net1250),
    .B(_08409_),
    .Y(_08410_));
 sky130_fd_sc_hd__o21a_1 _16348_ (.A1(net1087),
    .A2(net1081),
    .B1(net1085),
    .X(_08411_));
 sky130_fd_sc_hd__xnor2_1 _16349_ (.A(net1079),
    .B(_08411_),
    .Y(_08412_));
 sky130_fd_sc_hd__xnor2_2 _16350_ (.A(_08408_),
    .B(_08412_),
    .Y(_08413_));
 sky130_fd_sc_hd__a21o_1 _16351_ (.A1(net978),
    .A2(_08337_),
    .B1(_08333_),
    .X(_08414_));
 sky130_fd_sc_hd__o21ai_2 _16352_ (.A1(net978),
    .A2(_08337_),
    .B1(_08414_),
    .Y(_08415_));
 sky130_fd_sc_hd__o221a_1 _16353_ (.A1(net3522),
    .A2(net2222),
    .B1(_08312_),
    .B2(_07936_),
    .C1(_08329_),
    .X(_08416_));
 sky130_fd_sc_hd__and4_1 _16354_ (.A(net2651),
    .B(net3587),
    .C(net3431),
    .D(net1848),
    .X(_08417_));
 sky130_fd_sc_hd__nor2_1 _16355_ (.A(_08416_),
    .B(_08417_),
    .Y(_08418_));
 sky130_fd_sc_hd__and3_1 _16356_ (.A(net2691),
    .B(net2210),
    .C(_08313_),
    .X(_08419_));
 sky130_fd_sc_hd__xor2_1 _16357_ (.A(_08418_),
    .B(net1247),
    .X(_08420_));
 sky130_fd_sc_hd__xnor2_2 _16358_ (.A(_08415_),
    .B(_08420_),
    .Y(_08421_));
 sky130_fd_sc_hd__a21oi_1 _16359_ (.A1(_08339_),
    .A2(_08347_),
    .B1(_08349_),
    .Y(_08422_));
 sky130_fd_sc_hd__xor2_1 _16360_ (.A(_08421_),
    .B(_08422_),
    .X(_08423_));
 sky130_fd_sc_hd__xnor2_1 _16361_ (.A(_08413_),
    .B(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__a21o_1 _16362_ (.A1(_08311_),
    .A2(net1083),
    .B1(net1509),
    .X(_08425_));
 sky130_fd_sc_hd__o21ai_1 _16363_ (.A1(_08311_),
    .A2(net1083),
    .B1(_08425_),
    .Y(_08426_));
 sky130_fd_sc_hd__or2_2 _16364_ (.A(_08424_),
    .B(net773),
    .X(_08427_));
 sky130_fd_sc_hd__nand2_2 _16365_ (.A(_08424_),
    .B(net773),
    .Y(_08428_));
 sky130_fd_sc_hd__nand2_1 _16366_ (.A(_08427_),
    .B(_08428_),
    .Y(_08429_));
 sky130_fd_sc_hd__xnor2_1 _16367_ (.A(_08381_),
    .B(_08429_),
    .Y(_08430_));
 sky130_fd_sc_hd__xnor2_1 _16368_ (.A(net490),
    .B(_08430_),
    .Y(_08431_));
 sky130_fd_sc_hd__xnor2_1 _16369_ (.A(net303),
    .B(_08431_),
    .Y(_08432_));
 sky130_fd_sc_hd__mux2_1 _16370_ (.A0(\matmul0.matmul_stage_inst.mult1[11] ),
    .A1(net276),
    .S(net3478),
    .X(_08433_));
 sky130_fd_sc_hd__clkbuf_1 _16371_ (.A(_08433_),
    .X(_00226_));
 sky130_fd_sc_hd__a21o_1 _16372_ (.A1(_08418_),
    .A2(net1247),
    .B1(_08415_),
    .X(_08434_));
 sky130_fd_sc_hd__o21ai_1 _16373_ (.A1(_08418_),
    .A2(net1247),
    .B1(_08434_),
    .Y(_08435_));
 sky130_fd_sc_hd__o21ba_1 _16374_ (.A1(net1087),
    .A2(net1079),
    .B1_N(_08408_),
    .X(_08436_));
 sky130_fd_sc_hd__mux2_1 _16375_ (.A0(_08408_),
    .A1(net1087),
    .S(net1079),
    .X(_08437_));
 sky130_fd_sc_hd__o21ba_1 _16376_ (.A1(net1081),
    .A2(_08436_),
    .B1_N(_08437_),
    .X(_08438_));
 sky130_fd_sc_hd__nand2_1 _16377_ (.A(_08408_),
    .B(net1079),
    .Y(_08439_));
 sky130_fd_sc_hd__mux2_1 _16378_ (.A0(_08438_),
    .A1(_08439_),
    .S(net1252),
    .X(_08440_));
 sky130_fd_sc_hd__o21ai_1 _16379_ (.A1(net2841),
    .A2(net2682),
    .B1(net1250),
    .Y(_08441_));
 sky130_fd_sc_hd__nor2_1 _16380_ (.A(net2707),
    .B(net2648),
    .Y(_08442_));
 sky130_fd_sc_hd__o21ai_1 _16381_ (.A1(net1250),
    .A2(_08442_),
    .B1(net2815),
    .Y(_08443_));
 sky130_fd_sc_hd__a21o_1 _16382_ (.A1(_08441_),
    .A2(_08443_),
    .B1(net2629),
    .X(_08444_));
 sky130_fd_sc_hd__mux2_1 _16383_ (.A0(net1252),
    .A1(net1087),
    .S(net1079),
    .X(_08445_));
 sky130_fd_sc_hd__xor2_2 _16384_ (.A(net976),
    .B(_08445_),
    .X(_08446_));
 sky130_fd_sc_hd__a21bo_1 _16385_ (.A1(net1248),
    .A2(_08400_),
    .B1_N(_08399_),
    .X(_08447_));
 sky130_fd_sc_hd__nor2_1 _16386_ (.A(net2625),
    .B(net2218),
    .Y(_08448_));
 sky130_fd_sc_hd__nor2_1 _16387_ (.A(net2623),
    .B(net2631),
    .Y(_08449_));
 sky130_fd_sc_hd__clkbuf_1 _16388_ (.A(net3415),
    .X(_08450_));
 sky130_fd_sc_hd__nor2_1 _16389_ (.A(net2635),
    .B(net2622),
    .Y(_08451_));
 sky130_fd_sc_hd__xnor2_1 _16390_ (.A(_08449_),
    .B(_08451_),
    .Y(_08452_));
 sky130_fd_sc_hd__xnor2_2 _16391_ (.A(_08448_),
    .B(_08452_),
    .Y(_08453_));
 sky130_fd_sc_hd__nand2_1 _16392_ (.A(net2772),
    .B(net2642),
    .Y(_08454_));
 sky130_fd_sc_hd__nor2_1 _16393_ (.A(net2750),
    .B(_08454_),
    .Y(_08455_));
 sky130_fd_sc_hd__nor2_1 _16394_ (.A(net2791),
    .B(net2772),
    .Y(_08456_));
 sky130_fd_sc_hd__nor2_1 _16395_ (.A(net3402),
    .B(net2642),
    .Y(_08457_));
 sky130_fd_sc_hd__o22a_1 _16396_ (.A1(net2204),
    .A2(_08388_),
    .B1(_08457_),
    .B2(net2791),
    .X(_08458_));
 sky130_fd_sc_hd__o32a_1 _16397_ (.A1(net2783),
    .A2(_08455_),
    .A3(_08456_),
    .B1(_08458_),
    .B2(net2744),
    .X(_08459_));
 sky130_fd_sc_hd__or3_1 _16398_ (.A(net2245),
    .B(net2642),
    .C(net2639),
    .X(_08460_));
 sky130_fd_sc_hd__o31a_1 _16399_ (.A1(net2772),
    .A2(net2204),
    .A3(_08387_),
    .B1(_08460_),
    .X(_08461_));
 sky130_fd_sc_hd__a2111o_1 _16400_ (.A1(net2791),
    .A2(net2621),
    .B1(net2642),
    .C1(net2772),
    .D1(net2245),
    .X(_08462_));
 sky130_fd_sc_hd__o221a_1 _16401_ (.A1(net2628),
    .A2(_08459_),
    .B1(_08461_),
    .B2(net3402),
    .C1(_08462_),
    .X(_08463_));
 sky130_fd_sc_hd__xnor2_2 _16402_ (.A(_08453_),
    .B(net1246),
    .Y(_08464_));
 sky130_fd_sc_hd__xnor2_1 _16403_ (.A(_08447_),
    .B(_08464_),
    .Y(_08465_));
 sky130_fd_sc_hd__xnor2_1 _16404_ (.A(_08446_),
    .B(_08465_),
    .Y(_08466_));
 sky130_fd_sc_hd__o21ai_2 _16405_ (.A1(net882),
    .A2(_08405_),
    .B1(_08406_),
    .Y(_08467_));
 sky130_fd_sc_hd__or3_1 _16406_ (.A(net2625),
    .B(net2623),
    .C(net2213),
    .X(_08468_));
 sky130_fd_sc_hd__nand2_1 _16407_ (.A(net2654),
    .B(net2209),
    .Y(_08469_));
 sky130_fd_sc_hd__o31a_1 _16408_ (.A1(net2654),
    .A2(net2218),
    .A3(net1840),
    .B1(_08469_),
    .X(_08470_));
 sky130_fd_sc_hd__or2_1 _16409_ (.A(_08469_),
    .B(_08468_),
    .X(_08471_));
 sky130_fd_sc_hd__a21bo_1 _16410_ (.A1(_08468_),
    .A2(_08470_),
    .B1_N(_08471_),
    .X(_08472_));
 sky130_fd_sc_hd__xnor2_1 _16411_ (.A(net1507),
    .B(_08472_),
    .Y(_08473_));
 sky130_fd_sc_hd__xnor2_2 _16412_ (.A(_08467_),
    .B(_08473_),
    .Y(_08474_));
 sky130_fd_sc_hd__xor2_1 _16413_ (.A(_08466_),
    .B(_08474_),
    .X(_08475_));
 sky130_fd_sc_hd__xnor2_1 _16414_ (.A(_08440_),
    .B(_08475_),
    .Y(_08476_));
 sky130_fd_sc_hd__o21ba_1 _16415_ (.A1(_08421_),
    .A2(_08413_),
    .B1_N(_08422_),
    .X(_08477_));
 sky130_fd_sc_hd__a21o_1 _16416_ (.A1(_08421_),
    .A2(_08413_),
    .B1(_08477_),
    .X(_08478_));
 sky130_fd_sc_hd__xor2_1 _16417_ (.A(_08476_),
    .B(_08478_),
    .X(_08479_));
 sky130_fd_sc_hd__xnor2_2 _16418_ (.A(net723),
    .B(_08479_),
    .Y(_08480_));
 sky130_fd_sc_hd__nand2_1 _16419_ (.A(net490),
    .B(net571),
    .Y(_08481_));
 sky130_fd_sc_hd__or2_1 _16420_ (.A(net490),
    .B(net571),
    .X(_08482_));
 sky130_fd_sc_hd__inv_2 _16421_ (.A(_08427_),
    .Y(_08483_));
 sky130_fd_sc_hd__o21ai_1 _16422_ (.A1(_08381_),
    .A2(_08483_),
    .B1(_08428_),
    .Y(_08484_));
 sky130_fd_sc_hd__o22a_1 _16423_ (.A1(net571),
    .A2(_08427_),
    .B1(_08484_),
    .B2(net490),
    .X(_08485_));
 sky130_fd_sc_hd__o2bb2a_1 _16424_ (.A1_N(net490),
    .A2_N(_08484_),
    .B1(_08428_),
    .B2(_08381_),
    .X(_08486_));
 sky130_fd_sc_hd__mux2_1 _16425_ (.A0(_08485_),
    .A1(_08486_),
    .S(net303),
    .X(_08487_));
 sky130_fd_sc_hd__o221a_1 _16426_ (.A1(_08428_),
    .A2(_08481_),
    .B1(_08482_),
    .B2(_08427_),
    .C1(_08487_),
    .X(_08488_));
 sky130_fd_sc_hd__xor2_1 _16427_ (.A(_08480_),
    .B(_08488_),
    .X(_08489_));
 sky130_fd_sc_hd__mux2_1 _16428_ (.A0(\matmul0.matmul_stage_inst.mult1[12] ),
    .A1(net209),
    .S(net3475),
    .X(_08490_));
 sky130_fd_sc_hd__clkbuf_1 _16429_ (.A(_08490_),
    .X(_00227_));
 sky130_fd_sc_hd__nor2_1 _16430_ (.A(net490),
    .B(net571),
    .Y(_08491_));
 sky130_fd_sc_hd__a21bo_1 _16431_ (.A1(_08480_),
    .A2(_08481_),
    .B1_N(net303),
    .X(_08492_));
 sky130_fd_sc_hd__o21a_1 _16432_ (.A1(_08480_),
    .A2(_08491_),
    .B1(_08492_),
    .X(_08493_));
 sky130_fd_sc_hd__nand2_1 _16433_ (.A(net303),
    .B(_08482_),
    .Y(_08494_));
 sky130_fd_sc_hd__a22o_1 _16434_ (.A1(_08428_),
    .A2(_08480_),
    .B1(_08481_),
    .B2(_08494_),
    .X(_08495_));
 sky130_fd_sc_hd__o221a_1 _16435_ (.A1(_08428_),
    .A2(_08480_),
    .B1(_08493_),
    .B2(_08483_),
    .C1(_08495_),
    .X(_08496_));
 sky130_fd_sc_hd__and2_1 _16436_ (.A(net723),
    .B(_08478_),
    .X(_08497_));
 sky130_fd_sc_hd__or2_1 _16437_ (.A(net723),
    .B(_08478_),
    .X(_08498_));
 sky130_fd_sc_hd__o21a_1 _16438_ (.A1(_08476_),
    .A2(_08497_),
    .B1(_08498_),
    .X(_08499_));
 sky130_fd_sc_hd__a21o_1 _16439_ (.A1(_08466_),
    .A2(_08474_),
    .B1(_08440_),
    .X(_08500_));
 sky130_fd_sc_hd__o21ai_1 _16440_ (.A1(_08466_),
    .A2(_08474_),
    .B1(_08500_),
    .Y(_08501_));
 sky130_fd_sc_hd__xnor2_1 _16441_ (.A(net976),
    .B(_08465_),
    .Y(_08502_));
 sky130_fd_sc_hd__o21a_1 _16442_ (.A1(net1086),
    .A2(_08502_),
    .B1(net1078),
    .X(_08503_));
 sky130_fd_sc_hd__a21oi_1 _16443_ (.A1(net1084),
    .A2(_08502_),
    .B1(_08503_),
    .Y(_08504_));
 sky130_fd_sc_hd__inv_2 _16444_ (.A(_08453_),
    .Y(_08505_));
 sky130_fd_sc_hd__or3_1 _16445_ (.A(net2772),
    .B(net2621),
    .C(net2204),
    .X(_08506_));
 sky130_fd_sc_hd__a21o_1 _16446_ (.A1(_08389_),
    .A2(_08506_),
    .B1(_08387_),
    .X(_08507_));
 sky130_fd_sc_hd__or3_1 _16447_ (.A(net2621),
    .B(net2639),
    .C(_08389_),
    .X(_08508_));
 sky130_fd_sc_hd__a21o_1 _16448_ (.A1(_08507_),
    .A2(_08508_),
    .B1(net2245),
    .X(_08509_));
 sky130_fd_sc_hd__o21a_1 _16449_ (.A1(_08505_),
    .A2(net1246),
    .B1(net1245),
    .X(_08510_));
 sky130_fd_sc_hd__nor2_1 _16450_ (.A(net2634),
    .B(net2641),
    .Y(_08511_));
 sky130_fd_sc_hd__nor2_1 _16451_ (.A(net2623),
    .B(net2217),
    .Y(_08512_));
 sky130_fd_sc_hd__nor2_1 _16452_ (.A(net2622),
    .B(net2631),
    .Y(_08513_));
 sky130_fd_sc_hd__xnor2_1 _16453_ (.A(_08512_),
    .B(_08513_),
    .Y(_08514_));
 sky130_fd_sc_hd__xnor2_1 _16454_ (.A(_08511_),
    .B(_08514_),
    .Y(_08515_));
 sky130_fd_sc_hd__a21o_1 _16455_ (.A1(net2744),
    .A2(net2204),
    .B1(net2750),
    .X(_08516_));
 sky130_fd_sc_hd__a21oi_1 _16456_ (.A1(_08454_),
    .A2(_08516_),
    .B1(net2245),
    .Y(_08517_));
 sky130_fd_sc_hd__a211o_1 _16457_ (.A1(net2245),
    .A2(_08456_),
    .B1(_08517_),
    .C1(net2628),
    .X(_08518_));
 sky130_fd_sc_hd__xor2_2 _16458_ (.A(net1244),
    .B(_08518_),
    .X(_08519_));
 sky130_fd_sc_hd__xnor2_1 _16459_ (.A(_08510_),
    .B(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__xnor2_1 _16460_ (.A(_08446_),
    .B(net975),
    .Y(_08521_));
 sky130_fd_sc_hd__inv_2 _16461_ (.A(net976),
    .Y(_08522_));
 sky130_fd_sc_hd__o21a_1 _16462_ (.A1(_08447_),
    .A2(_08464_),
    .B1(_08522_),
    .X(_08523_));
 sky130_fd_sc_hd__a21o_1 _16463_ (.A1(_08447_),
    .A2(_08464_),
    .B1(_08523_),
    .X(_08524_));
 sky130_fd_sc_hd__nor2_1 _16464_ (.A(_08449_),
    .B(_08451_),
    .Y(_08525_));
 sky130_fd_sc_hd__or3_1 _16465_ (.A(net2623),
    .B(net2622),
    .C(net2213),
    .X(_08526_));
 sky130_fd_sc_hd__nand2_1 _16466_ (.A(net2625),
    .B(net2209),
    .Y(_08527_));
 sky130_fd_sc_hd__o311a_1 _16467_ (.A1(net2625),
    .A2(net2218),
    .A3(_08525_),
    .B1(_08526_),
    .C1(_08527_),
    .X(_08528_));
 sky130_fd_sc_hd__or2_1 _16468_ (.A(_08527_),
    .B(_08526_),
    .X(_08529_));
 sky130_fd_sc_hd__nor2b_1 _16469_ (.A(_08528_),
    .B_N(_08529_),
    .Y(_08530_));
 sky130_fd_sc_hd__xor2_1 _16470_ (.A(_08471_),
    .B(_08530_),
    .X(_08531_));
 sky130_fd_sc_hd__xnor2_2 _16471_ (.A(_08524_),
    .B(_08531_),
    .Y(_08532_));
 sky130_fd_sc_hd__xor2_1 _16472_ (.A(_08521_),
    .B(_08532_),
    .X(_08533_));
 sky130_fd_sc_hd__xnor2_1 _16473_ (.A(_08504_),
    .B(_08533_),
    .Y(_08534_));
 sky130_fd_sc_hd__o21ba_1 _16474_ (.A1(_08467_),
    .A2(_08472_),
    .B1_N(net1507),
    .X(_08535_));
 sky130_fd_sc_hd__a21oi_1 _16475_ (.A1(_08467_),
    .A2(_08472_),
    .B1(_08535_),
    .Y(_08536_));
 sky130_fd_sc_hd__or2b_1 _16476_ (.A(_08534_),
    .B_N(net671),
    .X(_08537_));
 sky130_fd_sc_hd__and2b_1 _16477_ (.A_N(net671),
    .B(_08534_),
    .X(_08538_));
 sky130_fd_sc_hd__inv_2 _16478_ (.A(_08538_),
    .Y(_08539_));
 sky130_fd_sc_hd__nand2_1 _16479_ (.A(_08537_),
    .B(_08539_),
    .Y(_08540_));
 sky130_fd_sc_hd__xnor2_1 _16480_ (.A(_08501_),
    .B(_08540_),
    .Y(_08541_));
 sky130_fd_sc_hd__nor2_1 _16481_ (.A(_08499_),
    .B(_08541_),
    .Y(_08542_));
 sky130_fd_sc_hd__nand2_1 _16482_ (.A(_08499_),
    .B(_08541_),
    .Y(_08543_));
 sky130_fd_sc_hd__or2b_1 _16483_ (.A(_08542_),
    .B_N(_08543_),
    .X(_08544_));
 sky130_fd_sc_hd__xnor2_1 _16484_ (.A(net208),
    .B(_08544_),
    .Y(_08545_));
 sky130_fd_sc_hd__mux2_1 _16485_ (.A0(\matmul0.matmul_stage_inst.mult1[13] ),
    .A1(net181),
    .S(net3475),
    .X(_08546_));
 sky130_fd_sc_hd__clkbuf_1 _16486_ (.A(_08546_),
    .X(_00228_));
 sky130_fd_sc_hd__o21ai_1 _16487_ (.A1(net208),
    .A2(_08542_),
    .B1(_08543_),
    .Y(_08547_));
 sky130_fd_sc_hd__a21o_1 _16488_ (.A1(_08501_),
    .A2(_08537_),
    .B1(_08538_),
    .X(_08548_));
 sky130_fd_sc_hd__a21o_1 _16489_ (.A1(_08521_),
    .A2(_08532_),
    .B1(_08504_),
    .X(_08549_));
 sky130_fd_sc_hd__o21a_1 _16490_ (.A1(_08521_),
    .A2(_08532_),
    .B1(_08549_),
    .X(_08550_));
 sky130_fd_sc_hd__nand2_1 _16491_ (.A(_08522_),
    .B(net975),
    .Y(_08551_));
 sky130_fd_sc_hd__or2_1 _16492_ (.A(_08522_),
    .B(net975),
    .X(_08552_));
 sky130_fd_sc_hd__o211a_1 _16493_ (.A1(net1084),
    .A2(net1078),
    .B1(_08551_),
    .C1(_08552_),
    .X(_08553_));
 sky130_fd_sc_hd__a21oi_2 _16494_ (.A1(net1086),
    .A2(net1078),
    .B1(_08553_),
    .Y(_08554_));
 sky130_fd_sc_hd__nor2_2 _16495_ (.A(net2634),
    .B(net2628),
    .Y(_08555_));
 sky130_fd_sc_hd__nor2_1 _16496_ (.A(net2621),
    .B(net2217),
    .Y(_08556_));
 sky130_fd_sc_hd__nor2_1 _16497_ (.A(net2631),
    .B(net2641),
    .Y(_08557_));
 sky130_fd_sc_hd__xnor2_1 _16498_ (.A(_08556_),
    .B(_08557_),
    .Y(_08558_));
 sky130_fd_sc_hd__xnor2_2 _16499_ (.A(_08555_),
    .B(_08558_),
    .Y(_08559_));
 sky130_fd_sc_hd__nand2_1 _16500_ (.A(net2772),
    .B(net2783),
    .Y(_08560_));
 sky130_fd_sc_hd__nand2_1 _16501_ (.A(net2750),
    .B(net2744),
    .Y(_08561_));
 sky130_fd_sc_hd__o221a_1 _16502_ (.A1(net2750),
    .A2(_08560_),
    .B1(_08561_),
    .B2(net2783),
    .C1(net2638),
    .X(_08562_));
 sky130_fd_sc_hd__xor2_1 _16503_ (.A(_08559_),
    .B(_08562_),
    .X(_08563_));
 sky130_fd_sc_hd__o31a_1 _16504_ (.A1(net2245),
    .A2(net2204),
    .A3(_08456_),
    .B1(net1244),
    .X(_08564_));
 sky130_fd_sc_hd__a21o_1 _16505_ (.A1(net2791),
    .A2(net2772),
    .B1(_08564_),
    .X(_08565_));
 sky130_fd_sc_hd__a21o_1 _16506_ (.A1(_08561_),
    .A2(net1244),
    .B1(net2784),
    .X(_08566_));
 sky130_fd_sc_hd__and4_1 _16507_ (.A(net2638),
    .B(_08563_),
    .C(_08565_),
    .D(_08566_),
    .X(_08567_));
 sky130_fd_sc_hd__a31oi_1 _16508_ (.A1(net2638),
    .A2(_08565_),
    .A3(_08566_),
    .B1(_08563_),
    .Y(_08568_));
 sky130_fd_sc_hd__or2_1 _16509_ (.A(net880),
    .B(net879),
    .X(_08569_));
 sky130_fd_sc_hd__xnor2_1 _16510_ (.A(net881),
    .B(_08569_),
    .Y(_08570_));
 sky130_fd_sc_hd__o21a_1 _16511_ (.A1(_08510_),
    .A2(_08519_),
    .B1(net977),
    .X(_08571_));
 sky130_fd_sc_hd__a21o_1 _16512_ (.A1(_08510_),
    .A2(_08519_),
    .B1(_08571_),
    .X(_08572_));
 sky130_fd_sc_hd__o21a_1 _16513_ (.A1(net2665),
    .A2(_08511_),
    .B1(_08513_),
    .X(_08573_));
 sky130_fd_sc_hd__a21o_1 _16514_ (.A1(net2665),
    .A2(_08511_),
    .B1(_08573_),
    .X(_08574_));
 sky130_fd_sc_hd__nand2_1 _16515_ (.A(_08511_),
    .B(_08513_),
    .Y(_08575_));
 sky130_fd_sc_hd__and3_1 _16516_ (.A(net2623),
    .B(net2208),
    .C(_08575_),
    .X(_08576_));
 sky130_fd_sc_hd__nor2_1 _16517_ (.A(net2208),
    .B(_08575_),
    .Y(_08577_));
 sky130_fd_sc_hd__a211o_1 _16518_ (.A1(net3420),
    .A2(_08574_),
    .B1(_08576_),
    .C1(_08577_),
    .X(_08578_));
 sky130_fd_sc_hd__xnor2_1 _16519_ (.A(_08529_),
    .B(net1243),
    .Y(_08579_));
 sky130_fd_sc_hd__xnor2_1 _16520_ (.A(_08572_),
    .B(_08579_),
    .Y(_08580_));
 sky130_fd_sc_hd__nor2_1 _16521_ (.A(_08570_),
    .B(_08580_),
    .Y(_08581_));
 sky130_fd_sc_hd__nand2_1 _16522_ (.A(_08570_),
    .B(_08580_),
    .Y(_08582_));
 sky130_fd_sc_hd__or2b_1 _16523_ (.A(_08581_),
    .B_N(_08582_),
    .X(_08583_));
 sky130_fd_sc_hd__a21bo_1 _16524_ (.A1(_08524_),
    .A2(_08530_),
    .B1_N(_08471_),
    .X(_08584_));
 sky130_fd_sc_hd__o21ai_2 _16525_ (.A1(_08524_),
    .A2(_08530_),
    .B1(_08584_),
    .Y(_08585_));
 sky130_fd_sc_hd__xnor2_1 _16526_ (.A(_08583_),
    .B(_08585_),
    .Y(_08586_));
 sky130_fd_sc_hd__xnor2_1 _16527_ (.A(_08554_),
    .B(_08586_),
    .Y(_08587_));
 sky130_fd_sc_hd__xnor2_1 _16528_ (.A(_08550_),
    .B(_08587_),
    .Y(_08588_));
 sky130_fd_sc_hd__and2_1 _16529_ (.A(_08548_),
    .B(_08588_),
    .X(_08589_));
 sky130_fd_sc_hd__or2_1 _16530_ (.A(_08548_),
    .B(_08588_),
    .X(_08590_));
 sky130_fd_sc_hd__or2b_1 _16531_ (.A(_08589_),
    .B_N(_08590_),
    .X(_08591_));
 sky130_fd_sc_hd__xor2_1 _16532_ (.A(_08547_),
    .B(_08591_),
    .X(_08592_));
 sky130_fd_sc_hd__mux2_1 _16533_ (.A0(\matmul0.matmul_stage_inst.mult1[14] ),
    .A1(net167),
    .S(net3474),
    .X(_08593_));
 sky130_fd_sc_hd__clkbuf_1 _16534_ (.A(_08593_),
    .X(_00229_));
 sky130_fd_sc_hd__nand2_1 _16535_ (.A(_08522_),
    .B(net880),
    .Y(_08594_));
 sky130_fd_sc_hd__nor2_1 _16536_ (.A(net1086),
    .B(_08594_),
    .Y(_08595_));
 sky130_fd_sc_hd__o21ba_1 _16537_ (.A1(net976),
    .A2(net879),
    .B1_N(net880),
    .X(_08596_));
 sky130_fd_sc_hd__o21ai_1 _16538_ (.A1(net1084),
    .A2(_08596_),
    .B1(_08594_),
    .Y(_08597_));
 sky130_fd_sc_hd__a22o_1 _16539_ (.A1(net976),
    .A2(net879),
    .B1(_08596_),
    .B2(net1086),
    .X(_08598_));
 sky130_fd_sc_hd__mux2_1 _16540_ (.A0(_08597_),
    .A1(_08598_),
    .S(net1078),
    .X(_08599_));
 sky130_fd_sc_hd__a311o_1 _16541_ (.A1(net1084),
    .A2(net976),
    .A3(net879),
    .B1(_08595_),
    .C1(_08599_),
    .X(_08600_));
 sky130_fd_sc_hd__nand2_1 _16542_ (.A(net2744),
    .B(net2245),
    .Y(_08601_));
 sky130_fd_sc_hd__or2b_1 _16543_ (.A(_08559_),
    .B_N(_08560_),
    .X(_08602_));
 sky130_fd_sc_hd__a22o_1 _16544_ (.A1(_08559_),
    .A2(_08601_),
    .B1(_08602_),
    .B2(net2791),
    .X(_08603_));
 sky130_fd_sc_hd__nand2_1 _16545_ (.A(net2638),
    .B(_08603_),
    .Y(_08604_));
 sky130_fd_sc_hd__xnor2_1 _16546_ (.A(net2634),
    .B(net2631),
    .Y(_08605_));
 sky130_fd_sc_hd__o211a_1 _16547_ (.A1(net2628),
    .A2(_08605_),
    .B1(net2621),
    .C1(net2208),
    .X(_08606_));
 sky130_fd_sc_hd__a211o_1 _16548_ (.A1(net2621),
    .A2(net2208),
    .B1(net2628),
    .C1(_08605_),
    .X(_08607_));
 sky130_fd_sc_hd__or2b_1 _16549_ (.A(_08606_),
    .B_N(_08607_),
    .X(_08608_));
 sky130_fd_sc_hd__a21o_1 _16550_ (.A1(_08555_),
    .A2(_08556_),
    .B1(_08557_),
    .X(_08609_));
 sky130_fd_sc_hd__o21a_1 _16551_ (.A1(_08555_),
    .A2(_08556_),
    .B1(_08609_),
    .X(_08610_));
 sky130_fd_sc_hd__xnor2_1 _16552_ (.A(_08562_),
    .B(_08610_),
    .Y(_08611_));
 sky130_fd_sc_hd__xnor2_1 _16553_ (.A(_08608_),
    .B(_08611_),
    .Y(_08612_));
 sky130_fd_sc_hd__a31o_1 _16554_ (.A1(net2624),
    .A2(net3401),
    .A3(net1847),
    .B1(net2664),
    .X(_08613_));
 sky130_fd_sc_hd__or4_1 _16555_ (.A(net3420),
    .B(net2622),
    .C(net2219),
    .D(net1841),
    .X(_08614_));
 sky130_fd_sc_hd__and3_1 _16556_ (.A(_08258_),
    .B(_08613_),
    .C(_08614_),
    .X(_08615_));
 sky130_fd_sc_hd__xnor2_1 _16557_ (.A(_08612_),
    .B(net1242),
    .Y(_08616_));
 sky130_fd_sc_hd__xnor2_1 _16558_ (.A(_08604_),
    .B(_08616_),
    .Y(_08617_));
 sky130_fd_sc_hd__xnor2_1 _16559_ (.A(net881),
    .B(_08617_),
    .Y(_08618_));
 sky130_fd_sc_hd__a21bo_1 _16560_ (.A1(_08529_),
    .A2(_08572_),
    .B1_N(net1243),
    .X(_08619_));
 sky130_fd_sc_hd__o21a_1 _16561_ (.A1(_08529_),
    .A2(_08572_),
    .B1(_08619_),
    .X(_08620_));
 sky130_fd_sc_hd__xnor2_1 _16562_ (.A(_08618_),
    .B(_08620_),
    .Y(_08621_));
 sky130_fd_sc_hd__xnor2_1 _16563_ (.A(_08600_),
    .B(_08621_),
    .Y(_08622_));
 sky130_fd_sc_hd__a21oi_1 _16564_ (.A1(_08582_),
    .A2(_08585_),
    .B1(_08581_),
    .Y(_08623_));
 sky130_fd_sc_hd__nand2_1 _16565_ (.A(_08581_),
    .B(_08585_),
    .Y(_08624_));
 sky130_fd_sc_hd__o21a_1 _16566_ (.A1(_08554_),
    .A2(_08623_),
    .B1(_08624_),
    .X(_08625_));
 sky130_fd_sc_hd__nor2_1 _16567_ (.A(_08550_),
    .B(_08625_),
    .Y(_08626_));
 sky130_fd_sc_hd__nor2_1 _16568_ (.A(_08554_),
    .B(_08624_),
    .Y(_08627_));
 sky130_fd_sc_hd__nor2_1 _16569_ (.A(_08582_),
    .B(_08585_),
    .Y(_08628_));
 sky130_fd_sc_hd__o21a_1 _16570_ (.A1(_08550_),
    .A2(_08554_),
    .B1(_08628_),
    .X(_08629_));
 sky130_fd_sc_hd__a31o_1 _16571_ (.A1(_08550_),
    .A2(_08554_),
    .A3(_08623_),
    .B1(_08629_),
    .X(_08630_));
 sky130_fd_sc_hd__or3_1 _16572_ (.A(_08626_),
    .B(_08627_),
    .C(_08630_),
    .X(_08631_));
 sky130_fd_sc_hd__xnor2_1 _16573_ (.A(_08622_),
    .B(_08631_),
    .Y(_08632_));
 sky130_fd_sc_hd__o21a_1 _16574_ (.A1(_08547_),
    .A2(_08589_),
    .B1(_08590_),
    .X(_08633_));
 sky130_fd_sc_hd__xnor2_1 _16575_ (.A(_08632_),
    .B(_08633_),
    .Y(_08634_));
 sky130_fd_sc_hd__mux2_1 _16576_ (.A0(\matmul0.matmul_stage_inst.mult1[15] ),
    .A1(net161),
    .S(net3474),
    .X(_08635_));
 sky130_fd_sc_hd__clkbuf_1 _16577_ (.A(_08635_),
    .X(_00230_));
 sky130_fd_sc_hd__buf_1 _16578_ (.A(net3471),
    .X(_08636_));
 sky130_fd_sc_hd__mux2_1 _16579_ (.A0(\matmul0.matmul_stage_inst.mult2[0] ),
    .A1(net494),
    .S(net2620),
    .X(_08637_));
 sky130_fd_sc_hd__clkbuf_1 _16580_ (.A(_08637_),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _16581_ (.A0(\matmul0.matmul_stage_inst.mult2[1] ),
    .A1(net440),
    .S(net2620),
    .X(_08638_));
 sky130_fd_sc_hd__clkbuf_1 _16582_ (.A(_08638_),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _16583_ (.A0(\matmul0.matmul_stage_inst.mult2[2] ),
    .A1(net433),
    .S(net2619),
    .X(_08639_));
 sky130_fd_sc_hd__clkbuf_1 _16584_ (.A(_08639_),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _16585_ (.A0(\matmul0.matmul_stage_inst.mult2[3] ),
    .A1(net426),
    .S(net2619),
    .X(_08640_));
 sky130_fd_sc_hd__clkbuf_1 _16586_ (.A(_08640_),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _16587_ (.A0(\matmul0.matmul_stage_inst.mult2[4] ),
    .A1(net396),
    .S(net2617),
    .X(_08641_));
 sky130_fd_sc_hd__clkbuf_1 _16588_ (.A(_08641_),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _16589_ (.A0(\matmul0.matmul_stage_inst.mult2[5] ),
    .A1(net389),
    .S(net2617),
    .X(_08642_));
 sky130_fd_sc_hd__clkbuf_1 _16590_ (.A(_08642_),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _16591_ (.A0(\matmul0.matmul_stage_inst.mult2[6] ),
    .A1(net359),
    .S(net2616),
    .X(_08643_));
 sky130_fd_sc_hd__clkbuf_1 _16592_ (.A(_08643_),
    .X(_00237_));
 sky130_fd_sc_hd__or2_1 _16593_ (.A(\svm0.state[1] ),
    .B(\svm0.state[0] ),
    .X(_08644_));
 sky130_fd_sc_hd__and2_1 _16594_ (.A(net5185),
    .B(net4253),
    .X(_08645_));
 sky130_fd_sc_hd__inv_2 _16595_ (.A(net6658),
    .Y(_08646_));
 sky130_fd_sc_hd__clkbuf_1 _16596_ (.A(_08646_),
    .X(_08647_));
 sky130_fd_sc_hd__mux2_1 _16597_ (.A0(_08644_),
    .A1(net3389),
    .S(net3388),
    .X(_08648_));
 sky130_fd_sc_hd__or2_1 _16598_ (.A(\svm0.delta[0] ),
    .B(net2614),
    .X(_08649_));
 sky130_fd_sc_hd__clkbuf_1 _16599_ (.A(_08649_),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _16600_ (.A0(\matmul0.matmul_stage_inst.mult2[7] ),
    .A1(net354),
    .S(net2616),
    .X(_08650_));
 sky130_fd_sc_hd__clkbuf_1 _16601_ (.A(_08650_),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _16602_ (.A0(\matmul0.matmul_stage_inst.mult2[8] ),
    .A1(net311),
    .S(net2618),
    .X(_08651_));
 sky130_fd_sc_hd__clkbuf_1 _16603_ (.A(_08651_),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _16604_ (.A0(\matmul0.matmul_stage_inst.mult2[9] ),
    .A1(net305),
    .S(net2618),
    .X(_08652_));
 sky130_fd_sc_hd__clkbuf_1 _16605_ (.A(_08652_),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _16606_ (.A0(\matmul0.matmul_stage_inst.mult2[10] ),
    .A1(net247),
    .S(net3471),
    .X(_08653_));
 sky130_fd_sc_hd__clkbuf_1 _16607_ (.A(_08653_),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _16608_ (.A0(\matmul0.matmul_stage_inst.mult2[11] ),
    .A1(net276),
    .S(net3471),
    .X(_08654_));
 sky130_fd_sc_hd__clkbuf_1 _16609_ (.A(_08654_),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _16610_ (.A0(\matmul0.matmul_stage_inst.mult2[12] ),
    .A1(net209),
    .S(net3468),
    .X(_08655_));
 sky130_fd_sc_hd__clkbuf_1 _16611_ (.A(_08655_),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _16612_ (.A0(\matmul0.matmul_stage_inst.mult2[13] ),
    .A1(net181),
    .S(net3468),
    .X(_08656_));
 sky130_fd_sc_hd__clkbuf_1 _16613_ (.A(_08656_),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _16614_ (.A0(\matmul0.matmul_stage_inst.mult2[14] ),
    .A1(net167),
    .S(net3467),
    .X(_08657_));
 sky130_fd_sc_hd__clkbuf_1 _16615_ (.A(_08657_),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _16616_ (.A0(\matmul0.matmul_stage_inst.mult2[15] ),
    .A1(net161),
    .S(net3467),
    .X(_08658_));
 sky130_fd_sc_hd__clkbuf_1 _16617_ (.A(_08658_),
    .X(_00247_));
 sky130_fd_sc_hd__xor2_1 _16618_ (.A(\matmul0.matmul_stage_inst.mult2[0] ),
    .B(\matmul0.matmul_stage_inst.mult1[0] ),
    .X(_08659_));
 sky130_fd_sc_hd__mux2_1 _16619_ (.A0(net7373),
    .A1(net4063),
    .S(net6558),
    .X(_08660_));
 sky130_fd_sc_hd__clkbuf_1 _16620_ (.A(_08660_),
    .X(_00248_));
 sky130_fd_sc_hd__nand2_1 _16621_ (.A(\matmul0.matmul_stage_inst.mult2[0] ),
    .B(\matmul0.matmul_stage_inst.mult1[0] ),
    .Y(_08661_));
 sky130_fd_sc_hd__xor2_1 _16622_ (.A(\matmul0.matmul_stage_inst.mult2[1] ),
    .B(\matmul0.matmul_stage_inst.mult1[1] ),
    .X(_08662_));
 sky130_fd_sc_hd__xnor2_1 _16623_ (.A(_08661_),
    .B(_08662_),
    .Y(_08663_));
 sky130_fd_sc_hd__mux2_1 _16624_ (.A0(\matmul0.alpha_pass[1] ),
    .A1(net3383),
    .S(net6551),
    .X(_08664_));
 sky130_fd_sc_hd__clkbuf_1 _16625_ (.A(_08664_),
    .X(_00249_));
 sky130_fd_sc_hd__nand2_1 _16626_ (.A(\matmul0.matmul_stage_inst.mult2[1] ),
    .B(\matmul0.matmul_stage_inst.mult1[1] ),
    .Y(_08665_));
 sky130_fd_sc_hd__o211ai_2 _16627_ (.A1(\matmul0.matmul_stage_inst.mult2[1] ),
    .A2(\matmul0.matmul_stage_inst.mult1[1] ),
    .B1(\matmul0.matmul_stage_inst.mult2[0] ),
    .C1(\matmul0.matmul_stage_inst.mult1[0] ),
    .Y(_08666_));
 sky130_fd_sc_hd__nand2_1 _16628_ (.A(_08665_),
    .B(_08666_),
    .Y(_08667_));
 sky130_fd_sc_hd__xnor2_1 _16629_ (.A(\matmul0.matmul_stage_inst.mult2[2] ),
    .B(\matmul0.matmul_stage_inst.mult1[2] ),
    .Y(_08668_));
 sky130_fd_sc_hd__xnor2_1 _16630_ (.A(_08667_),
    .B(_08668_),
    .Y(_08669_));
 sky130_fd_sc_hd__mux2_1 _16631_ (.A0(\matmul0.alpha_pass[2] ),
    .A1(net2613),
    .S(net6552),
    .X(_08670_));
 sky130_fd_sc_hd__clkbuf_1 _16632_ (.A(_08670_),
    .X(_00250_));
 sky130_fd_sc_hd__inv_2 _16633_ (.A(\matmul0.matmul_stage_inst.mult1[2] ),
    .Y(_08671_));
 sky130_fd_sc_hd__a21o_1 _16634_ (.A1(_08665_),
    .A2(_08666_),
    .B1(_08671_),
    .X(_08672_));
 sky130_fd_sc_hd__inv_2 _16635_ (.A(\matmul0.matmul_stage_inst.mult2[2] ),
    .Y(_08673_));
 sky130_fd_sc_hd__a31o_1 _16636_ (.A1(_08671_),
    .A2(_08665_),
    .A3(_08666_),
    .B1(_08673_),
    .X(_08674_));
 sky130_fd_sc_hd__nand2_1 _16637_ (.A(_08672_),
    .B(_08674_),
    .Y(_08675_));
 sky130_fd_sc_hd__xnor2_1 _16638_ (.A(\matmul0.matmul_stage_inst.mult2[3] ),
    .B(\matmul0.matmul_stage_inst.mult1[3] ),
    .Y(_08676_));
 sky130_fd_sc_hd__xnor2_1 _16639_ (.A(_08675_),
    .B(_08676_),
    .Y(_08677_));
 sky130_fd_sc_hd__mux2_1 _16640_ (.A0(\matmul0.alpha_pass[3] ),
    .A1(net2202),
    .S(net6552),
    .X(_08678_));
 sky130_fd_sc_hd__clkbuf_1 _16641_ (.A(_08678_),
    .X(_00251_));
 sky130_fd_sc_hd__inv_2 _16642_ (.A(\matmul0.matmul_stage_inst.mult1[3] ),
    .Y(_08679_));
 sky130_fd_sc_hd__inv_2 _16643_ (.A(\matmul0.matmul_stage_inst.mult2[3] ),
    .Y(_08680_));
 sky130_fd_sc_hd__a31o_1 _16644_ (.A1(_08679_),
    .A2(_08672_),
    .A3(_08674_),
    .B1(_08680_),
    .X(_08681_));
 sky130_fd_sc_hd__a21boi_2 _16645_ (.A1(\matmul0.matmul_stage_inst.mult1[3] ),
    .A2(_08675_),
    .B1_N(_08681_),
    .Y(_08682_));
 sky130_fd_sc_hd__xor2_1 _16646_ (.A(\matmul0.matmul_stage_inst.mult2[4] ),
    .B(\matmul0.matmul_stage_inst.mult1[4] ),
    .X(_08683_));
 sky130_fd_sc_hd__xnor2_1 _16647_ (.A(_08682_),
    .B(_08683_),
    .Y(_08684_));
 sky130_fd_sc_hd__mux2_1 _16648_ (.A0(net7328),
    .A1(net1838),
    .S(net6551),
    .X(_08685_));
 sky130_fd_sc_hd__clkbuf_1 _16649_ (.A(_08685_),
    .X(_00252_));
 sky130_fd_sc_hd__inv_2 _16650_ (.A(\matmul0.matmul_stage_inst.mult1[4] ),
    .Y(_08686_));
 sky130_fd_sc_hd__o21ba_1 _16651_ (.A1(_08686_),
    .A2(_08682_),
    .B1_N(\matmul0.matmul_stage_inst.mult2[4] ),
    .X(_08687_));
 sky130_fd_sc_hd__a21o_1 _16652_ (.A1(_08686_),
    .A2(_08682_),
    .B1(_08687_),
    .X(_08688_));
 sky130_fd_sc_hd__xor2_1 _16653_ (.A(\matmul0.matmul_stage_inst.mult2[5] ),
    .B(\matmul0.matmul_stage_inst.mult1[5] ),
    .X(_08689_));
 sky130_fd_sc_hd__xnor2_1 _16654_ (.A(_08688_),
    .B(_08689_),
    .Y(_08690_));
 sky130_fd_sc_hd__mux2_1 _16655_ (.A0(net7316),
    .A1(net1240),
    .S(net6554),
    .X(_08691_));
 sky130_fd_sc_hd__clkbuf_1 _16656_ (.A(_08691_),
    .X(_00253_));
 sky130_fd_sc_hd__inv_2 _16657_ (.A(\matmul0.matmul_stage_inst.mult1[5] ),
    .Y(_08692_));
 sky130_fd_sc_hd__o21ba_1 _16658_ (.A1(_08692_),
    .A2(_08688_),
    .B1_N(\matmul0.matmul_stage_inst.mult2[5] ),
    .X(_08693_));
 sky130_fd_sc_hd__a21o_1 _16659_ (.A1(_08692_),
    .A2(_08688_),
    .B1(_08693_),
    .X(_08694_));
 sky130_fd_sc_hd__xor2_1 _16660_ (.A(\matmul0.matmul_stage_inst.mult2[6] ),
    .B(\matmul0.matmul_stage_inst.mult1[6] ),
    .X(_08695_));
 sky130_fd_sc_hd__xnor2_1 _16661_ (.A(_08694_),
    .B(_08695_),
    .Y(_08696_));
 sky130_fd_sc_hd__mux2_1 _16662_ (.A0(\matmul0.alpha_pass[6] ),
    .A1(net972),
    .S(net6563),
    .X(_08697_));
 sky130_fd_sc_hd__clkbuf_1 _16663_ (.A(_08697_),
    .X(_00254_));
 sky130_fd_sc_hd__inv_2 _16664_ (.A(\matmul0.matmul_stage_inst.mult1[6] ),
    .Y(_08698_));
 sky130_fd_sc_hd__o21ba_1 _16665_ (.A1(_08698_),
    .A2(_08694_),
    .B1_N(\matmul0.matmul_stage_inst.mult2[6] ),
    .X(_08699_));
 sky130_fd_sc_hd__a21o_1 _16666_ (.A1(_08698_),
    .A2(_08694_),
    .B1(_08699_),
    .X(_08700_));
 sky130_fd_sc_hd__xor2_1 _16667_ (.A(\matmul0.matmul_stage_inst.mult2[7] ),
    .B(\matmul0.matmul_stage_inst.mult1[7] ),
    .X(_08701_));
 sky130_fd_sc_hd__xnor2_1 _16668_ (.A(_08700_),
    .B(_08701_),
    .Y(_08702_));
 sky130_fd_sc_hd__mux2_1 _16669_ (.A0(\matmul0.alpha_pass[7] ),
    .A1(net823),
    .S(net6563),
    .X(_08703_));
 sky130_fd_sc_hd__clkbuf_1 _16670_ (.A(_08703_),
    .X(_00255_));
 sky130_fd_sc_hd__inv_2 _16671_ (.A(\matmul0.matmul_stage_inst.mult1[7] ),
    .Y(_08704_));
 sky130_fd_sc_hd__a21bo_1 _16672_ (.A1(_08704_),
    .A2(_08700_),
    .B1_N(\matmul0.matmul_stage_inst.mult2[7] ),
    .X(_08705_));
 sky130_fd_sc_hd__o21a_1 _16673_ (.A1(_08704_),
    .A2(_08700_),
    .B1(_08705_),
    .X(_08706_));
 sky130_fd_sc_hd__xor2_1 _16674_ (.A(\matmul0.matmul_stage_inst.mult2[8] ),
    .B(\matmul0.matmul_stage_inst.mult1[8] ),
    .X(_08707_));
 sky130_fd_sc_hd__xnor2_1 _16675_ (.A(_08706_),
    .B(_08707_),
    .Y(_08708_));
 sky130_fd_sc_hd__mux2_1 _16676_ (.A0(net7281),
    .A1(net720),
    .S(net6549),
    .X(_08709_));
 sky130_fd_sc_hd__clkbuf_1 _16677_ (.A(_08709_),
    .X(_00256_));
 sky130_fd_sc_hd__inv_2 _16678_ (.A(\matmul0.matmul_stage_inst.mult1[8] ),
    .Y(_08710_));
 sky130_fd_sc_hd__o21ba_1 _16679_ (.A1(_08710_),
    .A2(_08706_),
    .B1_N(\matmul0.matmul_stage_inst.mult2[8] ),
    .X(_08711_));
 sky130_fd_sc_hd__a21o_1 _16680_ (.A1(_08710_),
    .A2(_08706_),
    .B1(_08711_),
    .X(_08712_));
 sky130_fd_sc_hd__xor2_1 _16681_ (.A(\matmul0.matmul_stage_inst.mult2[9] ),
    .B(\matmul0.matmul_stage_inst.mult1[9] ),
    .X(_08713_));
 sky130_fd_sc_hd__xnor2_1 _16682_ (.A(_08712_),
    .B(_08713_),
    .Y(_08714_));
 sky130_fd_sc_hd__mux2_1 _16683_ (.A0(\matmul0.alpha_pass[9] ),
    .A1(net619),
    .S(net6550),
    .X(_08715_));
 sky130_fd_sc_hd__clkbuf_1 _16684_ (.A(_08715_),
    .X(_00257_));
 sky130_fd_sc_hd__inv_2 _16685_ (.A(\matmul0.matmul_stage_inst.mult1[9] ),
    .Y(_08716_));
 sky130_fd_sc_hd__o21ba_1 _16686_ (.A1(_08716_),
    .A2(_08712_),
    .B1_N(\matmul0.matmul_stage_inst.mult2[9] ),
    .X(_08717_));
 sky130_fd_sc_hd__a21o_1 _16687_ (.A1(_08716_),
    .A2(_08712_),
    .B1(_08717_),
    .X(_08718_));
 sky130_fd_sc_hd__xor2_1 _16688_ (.A(\matmul0.matmul_stage_inst.mult2[10] ),
    .B(\matmul0.matmul_stage_inst.mult1[10] ),
    .X(_08719_));
 sky130_fd_sc_hd__xnor2_1 _16689_ (.A(_08718_),
    .B(_08719_),
    .Y(_08720_));
 sky130_fd_sc_hd__mux2_1 _16690_ (.A0(\matmul0.alpha_pass[10] ),
    .A1(net528),
    .S(net6550),
    .X(_08721_));
 sky130_fd_sc_hd__clkbuf_1 _16691_ (.A(_08721_),
    .X(_00258_));
 sky130_fd_sc_hd__inv_2 _16692_ (.A(\matmul0.matmul_stage_inst.mult1[10] ),
    .Y(_08722_));
 sky130_fd_sc_hd__o21ba_1 _16693_ (.A1(_08722_),
    .A2(_08718_),
    .B1_N(\matmul0.matmul_stage_inst.mult2[10] ),
    .X(_08723_));
 sky130_fd_sc_hd__a21o_1 _16694_ (.A1(_08722_),
    .A2(_08718_),
    .B1(_08723_),
    .X(_08724_));
 sky130_fd_sc_hd__xor2_1 _16695_ (.A(\matmul0.matmul_stage_inst.mult2[11] ),
    .B(\matmul0.matmul_stage_inst.mult1[11] ),
    .X(_08725_));
 sky130_fd_sc_hd__xnor2_1 _16696_ (.A(_08724_),
    .B(_08725_),
    .Y(_08726_));
 sky130_fd_sc_hd__mux2_1 _16697_ (.A0(\matmul0.alpha_pass[11] ),
    .A1(net423),
    .S(net6550),
    .X(_08727_));
 sky130_fd_sc_hd__clkbuf_1 _16698_ (.A(_08727_),
    .X(_00259_));
 sky130_fd_sc_hd__inv_2 _16699_ (.A(\matmul0.matmul_stage_inst.mult1[11] ),
    .Y(_08728_));
 sky130_fd_sc_hd__o21ba_1 _16700_ (.A1(_08728_),
    .A2(_08724_),
    .B1_N(\matmul0.matmul_stage_inst.mult2[11] ),
    .X(_08729_));
 sky130_fd_sc_hd__a21o_1 _16701_ (.A1(_08728_),
    .A2(_08724_),
    .B1(_08729_),
    .X(_08730_));
 sky130_fd_sc_hd__xor2_1 _16702_ (.A(\matmul0.matmul_stage_inst.mult2[12] ),
    .B(\matmul0.matmul_stage_inst.mult1[12] ),
    .X(_08731_));
 sky130_fd_sc_hd__xnor2_1 _16703_ (.A(net383),
    .B(_08731_),
    .Y(_08732_));
 sky130_fd_sc_hd__mux2_1 _16704_ (.A0(\matmul0.alpha_pass[12] ),
    .A1(net353),
    .S(net6557),
    .X(_08733_));
 sky130_fd_sc_hd__clkbuf_1 _16705_ (.A(_08733_),
    .X(_00260_));
 sky130_fd_sc_hd__inv_2 _16706_ (.A(\matmul0.matmul_stage_inst.mult1[12] ),
    .Y(_08734_));
 sky130_fd_sc_hd__o21ba_1 _16707_ (.A1(_08734_),
    .A2(net383),
    .B1_N(\matmul0.matmul_stage_inst.mult2[12] ),
    .X(_08735_));
 sky130_fd_sc_hd__a21o_1 _16708_ (.A1(_08734_),
    .A2(net383),
    .B1(_08735_),
    .X(_08736_));
 sky130_fd_sc_hd__xor2_1 _16709_ (.A(net7375),
    .B(\matmul0.matmul_stage_inst.mult1[13] ),
    .X(_08737_));
 sky130_fd_sc_hd__xnor2_1 _16710_ (.A(_08736_),
    .B(_08737_),
    .Y(_08738_));
 sky130_fd_sc_hd__mux2_1 _16711_ (.A0(net7224),
    .A1(_08738_),
    .S(net6548),
    .X(_08739_));
 sky130_fd_sc_hd__clkbuf_1 _16712_ (.A(_08739_),
    .X(_00261_));
 sky130_fd_sc_hd__inv_2 _16713_ (.A(\matmul0.matmul_stage_inst.mult1[13] ),
    .Y(_08740_));
 sky130_fd_sc_hd__o21ba_1 _16714_ (.A1(_08740_),
    .A2(_08736_),
    .B1_N(net7375),
    .X(_08741_));
 sky130_fd_sc_hd__a21o_1 _16715_ (.A1(_08740_),
    .A2(_08736_),
    .B1(_08741_),
    .X(_08742_));
 sky130_fd_sc_hd__xor2_1 _16716_ (.A(\matmul0.matmul_stage_inst.mult2[14] ),
    .B(\matmul0.matmul_stage_inst.mult1[14] ),
    .X(_08743_));
 sky130_fd_sc_hd__xnor2_1 _16717_ (.A(_08742_),
    .B(_08743_),
    .Y(_08744_));
 sky130_fd_sc_hd__mux2_1 _16718_ (.A0(\matmul0.alpha_pass[14] ),
    .A1(_08744_),
    .S(net6557),
    .X(_08745_));
 sky130_fd_sc_hd__clkbuf_1 _16719_ (.A(_08745_),
    .X(_00262_));
 sky130_fd_sc_hd__xor2_1 _16720_ (.A(\matmul0.matmul_stage_inst.mult2[15] ),
    .B(\matmul0.matmul_stage_inst.mult1[15] ),
    .X(_08746_));
 sky130_fd_sc_hd__nor2_1 _16721_ (.A(\matmul0.matmul_stage_inst.mult2[14] ),
    .B(\matmul0.matmul_stage_inst.mult1[14] ),
    .Y(_08747_));
 sky130_fd_sc_hd__nand2_1 _16722_ (.A(\matmul0.matmul_stage_inst.mult2[14] ),
    .B(\matmul0.matmul_stage_inst.mult1[14] ),
    .Y(_08748_));
 sky130_fd_sc_hd__o21a_1 _16723_ (.A1(_08742_),
    .A2(_08747_),
    .B1(_08748_),
    .X(_08749_));
 sky130_fd_sc_hd__xnor2_1 _16724_ (.A(_08746_),
    .B(_08749_),
    .Y(_08750_));
 sky130_fd_sc_hd__mux2_1 _16725_ (.A0(\matmul0.alpha_pass[15] ),
    .A1(_08750_),
    .S(net6557),
    .X(_08751_));
 sky130_fd_sc_hd__clkbuf_1 _16726_ (.A(_08751_),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _16727_ (.A0(net7575),
    .A1(\matmul0.b[0] ),
    .S(net3702),
    .X(_08752_));
 sky130_fd_sc_hd__clkbuf_1 _16728_ (.A(_08752_),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _16729_ (.A0(net7574),
    .A1(\matmul0.b[1] ),
    .S(net3702),
    .X(_08753_));
 sky130_fd_sc_hd__clkbuf_1 _16730_ (.A(_08753_),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _16731_ (.A0(\matmul0.b_in[2] ),
    .A1(\matmul0.b[2] ),
    .S(net3703),
    .X(_08754_));
 sky130_fd_sc_hd__clkbuf_1 _16732_ (.A(_08754_),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _16733_ (.A0(net7573),
    .A1(\matmul0.b[3] ),
    .S(net3702),
    .X(_08755_));
 sky130_fd_sc_hd__clkbuf_1 _16734_ (.A(_08755_),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _16735_ (.A0(net9226),
    .A1(\matmul0.b[4] ),
    .S(net3703),
    .X(_08756_));
 sky130_fd_sc_hd__clkbuf_1 _16736_ (.A(_08756_),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _16737_ (.A0(net7571),
    .A1(\matmul0.b[5] ),
    .S(net3702),
    .X(_08757_));
 sky130_fd_sc_hd__clkbuf_1 _16738_ (.A(_08757_),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _16739_ (.A0(net7568),
    .A1(\matmul0.b[6] ),
    .S(net3702),
    .X(_08758_));
 sky130_fd_sc_hd__clkbuf_1 _16740_ (.A(_08758_),
    .X(_00270_));
 sky130_fd_sc_hd__clkbuf_1 _16741_ (.A(net4291),
    .X(_08759_));
 sky130_fd_sc_hd__mux2_1 _16742_ (.A0(net7567),
    .A1(\matmul0.b[7] ),
    .S(net3381),
    .X(_08760_));
 sky130_fd_sc_hd__clkbuf_1 _16743_ (.A(_08760_),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _16744_ (.A0(\matmul0.b_in[8] ),
    .A1(\matmul0.b[8] ),
    .S(net3381),
    .X(_08761_));
 sky130_fd_sc_hd__clkbuf_1 _16745_ (.A(_08761_),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _16746_ (.A0(net7566),
    .A1(\matmul0.b[9] ),
    .S(net3380),
    .X(_08762_));
 sky130_fd_sc_hd__clkbuf_1 _16747_ (.A(_08762_),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _16748_ (.A0(net7564),
    .A1(\matmul0.b[10] ),
    .S(net3380),
    .X(_08763_));
 sky130_fd_sc_hd__clkbuf_1 _16749_ (.A(_08763_),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _16750_ (.A0(net7562),
    .A1(net9242),
    .S(net3380),
    .X(_08764_));
 sky130_fd_sc_hd__clkbuf_1 _16751_ (.A(_08764_),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _16752_ (.A0(net7561),
    .A1(net9230),
    .S(net3380),
    .X(_08765_));
 sky130_fd_sc_hd__clkbuf_1 _16753_ (.A(_08765_),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _16754_ (.A0(net7559),
    .A1(\matmul0.b[13] ),
    .S(net3381),
    .X(_08766_));
 sky130_fd_sc_hd__clkbuf_1 _16755_ (.A(_08766_),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _16756_ (.A0(net7556),
    .A1(\matmul0.b[14] ),
    .S(net3381),
    .X(_08767_));
 sky130_fd_sc_hd__clkbuf_1 _16757_ (.A(_08767_),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _16758_ (.A0(net7553),
    .A1(\matmul0.b[15] ),
    .S(net3382),
    .X(_08768_));
 sky130_fd_sc_hd__clkbuf_1 _16759_ (.A(_08768_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _16760_ (.A0(\matmul0.a_in[0] ),
    .A1(\matmul0.a[0] ),
    .S(net3382),
    .X(_08769_));
 sky130_fd_sc_hd__clkbuf_1 _16761_ (.A(_08769_),
    .X(_00280_));
 sky130_fd_sc_hd__clkbuf_2 _16762_ (.A(net4291),
    .X(_08770_));
 sky130_fd_sc_hd__mux2_1 _16763_ (.A0(\matmul0.a_in[1] ),
    .A1(\matmul0.a[1] ),
    .S(net3378),
    .X(_08771_));
 sky130_fd_sc_hd__clkbuf_1 _16764_ (.A(_08771_),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _16765_ (.A0(\matmul0.a_in[2] ),
    .A1(\matmul0.a[2] ),
    .S(net3378),
    .X(_08772_));
 sky130_fd_sc_hd__clkbuf_1 _16766_ (.A(_08772_),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _16767_ (.A0(net9158),
    .A1(\matmul0.a[3] ),
    .S(net3378),
    .X(_08773_));
 sky130_fd_sc_hd__clkbuf_1 _16768_ (.A(_08773_),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _16769_ (.A0(\matmul0.a_in[4] ),
    .A1(\matmul0.a[4] ),
    .S(net3378),
    .X(_08774_));
 sky130_fd_sc_hd__clkbuf_1 _16770_ (.A(_08774_),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _16771_ (.A0(\matmul0.a_in[5] ),
    .A1(\matmul0.a[5] ),
    .S(net3378),
    .X(_08775_));
 sky130_fd_sc_hd__clkbuf_1 _16772_ (.A(_08775_),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _16773_ (.A0(\matmul0.a_in[6] ),
    .A1(\matmul0.a[6] ),
    .S(_08770_),
    .X(_08776_));
 sky130_fd_sc_hd__clkbuf_1 _16774_ (.A(_08776_),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _16775_ (.A0(\matmul0.a_in[7] ),
    .A1(\matmul0.a[7] ),
    .S(_08770_),
    .X(_08777_));
 sky130_fd_sc_hd__clkbuf_1 _16776_ (.A(_08777_),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _16777_ (.A0(net7600),
    .A1(\matmul0.a[8] ),
    .S(_08770_),
    .X(_08778_));
 sky130_fd_sc_hd__clkbuf_1 _16778_ (.A(_08778_),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _16779_ (.A0(net7598),
    .A1(\matmul0.a[9] ),
    .S(net3379),
    .X(_08779_));
 sky130_fd_sc_hd__clkbuf_1 _16780_ (.A(_08779_),
    .X(_00289_));
 sky130_fd_sc_hd__mux2_1 _16781_ (.A0(net7595),
    .A1(\matmul0.a[10] ),
    .S(net3379),
    .X(_08780_));
 sky130_fd_sc_hd__clkbuf_1 _16782_ (.A(_08780_),
    .X(_00290_));
 sky130_fd_sc_hd__clkbuf_1 _16783_ (.A(net4289),
    .X(_08781_));
 sky130_fd_sc_hd__mux2_1 _16784_ (.A0(net7592),
    .A1(\matmul0.a[11] ),
    .S(net3373),
    .X(_08782_));
 sky130_fd_sc_hd__clkbuf_1 _16785_ (.A(_08782_),
    .X(_00291_));
 sky130_fd_sc_hd__mux2_1 _16786_ (.A0(net7589),
    .A1(\matmul0.a[12] ),
    .S(net3372),
    .X(_08783_));
 sky130_fd_sc_hd__clkbuf_1 _16787_ (.A(_08783_),
    .X(_00292_));
 sky130_fd_sc_hd__mux2_1 _16788_ (.A0(net7585),
    .A1(\matmul0.a[13] ),
    .S(net3372),
    .X(_08784_));
 sky130_fd_sc_hd__clkbuf_1 _16789_ (.A(_08784_),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _16790_ (.A0(net7581),
    .A1(\matmul0.a[14] ),
    .S(net3373),
    .X(_08785_));
 sky130_fd_sc_hd__clkbuf_1 _16791_ (.A(_08785_),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _16792_ (.A0(net7577),
    .A1(\matmul0.a[15] ),
    .S(net3373),
    .X(_08786_));
 sky130_fd_sc_hd__clkbuf_1 _16793_ (.A(_08786_),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _16794_ (.A0(\cordic0.cos[0] ),
    .A1(\matmul0.cos[0] ),
    .S(net3370),
    .X(_08787_));
 sky130_fd_sc_hd__clkbuf_1 _16795_ (.A(_08787_),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_1 _16796_ (.A0(net9240),
    .A1(net7182),
    .S(net3369),
    .X(_08788_));
 sky130_fd_sc_hd__clkbuf_1 _16797_ (.A(_08788_),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_1 _16798_ (.A0(\cordic0.cos[2] ),
    .A1(\matmul0.cos[2] ),
    .S(net3370),
    .X(_08789_));
 sky130_fd_sc_hd__clkbuf_1 _16799_ (.A(_08789_),
    .X(_00298_));
 sky130_fd_sc_hd__mux2_1 _16800_ (.A0(net8968),
    .A1(\matmul0.cos[3] ),
    .S(net3370),
    .X(_08790_));
 sky130_fd_sc_hd__clkbuf_1 _16801_ (.A(_08790_),
    .X(_00299_));
 sky130_fd_sc_hd__mux2_1 _16802_ (.A0(\cordic0.cos[4] ),
    .A1(net7180),
    .S(net3369),
    .X(_08791_));
 sky130_fd_sc_hd__clkbuf_1 _16803_ (.A(_08791_),
    .X(_00300_));
 sky130_fd_sc_hd__buf_1 _16804_ (.A(net4287),
    .X(_08792_));
 sky130_fd_sc_hd__mux2_1 _16805_ (.A0(net9241),
    .A1(\matmul0.cos[5] ),
    .S(_08792_),
    .X(_08793_));
 sky130_fd_sc_hd__clkbuf_1 _16806_ (.A(_08793_),
    .X(_00301_));
 sky130_fd_sc_hd__mux2_1 _16807_ (.A0(net8975),
    .A1(\matmul0.cos[6] ),
    .S(net3368),
    .X(_08794_));
 sky130_fd_sc_hd__clkbuf_1 _16808_ (.A(_08794_),
    .X(_00302_));
 sky130_fd_sc_hd__mux2_1 _16809_ (.A0(net9038),
    .A1(\matmul0.cos[7] ),
    .S(net3367),
    .X(_08795_));
 sky130_fd_sc_hd__clkbuf_1 _16810_ (.A(_08795_),
    .X(_00303_));
 sky130_fd_sc_hd__mux2_1 _16811_ (.A0(\cordic0.cos[8] ),
    .A1(\matmul0.cos[8] ),
    .S(net3367),
    .X(_08796_));
 sky130_fd_sc_hd__clkbuf_1 _16812_ (.A(_08796_),
    .X(_00304_));
 sky130_fd_sc_hd__mux2_1 _16813_ (.A0(net8972),
    .A1(\matmul0.cos[9] ),
    .S(net3367),
    .X(_08797_));
 sky130_fd_sc_hd__clkbuf_1 _16814_ (.A(_08797_),
    .X(_00305_));
 sky130_fd_sc_hd__mux2_1 _16815_ (.A0(\cordic0.cos[10] ),
    .A1(\matmul0.cos[10] ),
    .S(net3368),
    .X(_08798_));
 sky130_fd_sc_hd__clkbuf_1 _16816_ (.A(_08798_),
    .X(_00306_));
 sky130_fd_sc_hd__mux2_1 _16817_ (.A0(net9210),
    .A1(\matmul0.cos[11] ),
    .S(net3368),
    .X(_08799_));
 sky130_fd_sc_hd__clkbuf_1 _16818_ (.A(_08799_),
    .X(_00307_));
 sky130_fd_sc_hd__mux2_1 _16819_ (.A0(\cordic0.cos[12] ),
    .A1(\matmul0.cos[12] ),
    .S(_08792_),
    .X(_08800_));
 sky130_fd_sc_hd__clkbuf_1 _16820_ (.A(_08800_),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_1 _16821_ (.A0(net9233),
    .A1(\matmul0.cos[13] ),
    .S(net3368),
    .X(_08801_));
 sky130_fd_sc_hd__clkbuf_1 _16822_ (.A(_08801_),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_1 _16823_ (.A0(net6431),
    .A1(\matmul0.sin[0] ),
    .S(net3367),
    .X(_08802_));
 sky130_fd_sc_hd__clkbuf_1 _16824_ (.A(_08802_),
    .X(_00310_));
 sky130_fd_sc_hd__buf_1 _16825_ (.A(net4287),
    .X(_08803_));
 sky130_fd_sc_hd__mux2_1 _16826_ (.A0(net6430),
    .A1(\matmul0.sin[1] ),
    .S(net3365),
    .X(_08804_));
 sky130_fd_sc_hd__clkbuf_1 _16827_ (.A(_08804_),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _16828_ (.A0(\cordic0.sin[2] ),
    .A1(\matmul0.sin[2] ),
    .S(net3365),
    .X(_08805_));
 sky130_fd_sc_hd__clkbuf_1 _16829_ (.A(_08805_),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _16830_ (.A0(net6428),
    .A1(\matmul0.sin[3] ),
    .S(net3365),
    .X(_08806_));
 sky130_fd_sc_hd__clkbuf_1 _16831_ (.A(_08806_),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _16832_ (.A0(net6427),
    .A1(\matmul0.sin[4] ),
    .S(_08803_),
    .X(_08807_));
 sky130_fd_sc_hd__clkbuf_1 _16833_ (.A(_08807_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _16834_ (.A0(net6425),
    .A1(\matmul0.sin[5] ),
    .S(net3366),
    .X(_08808_));
 sky130_fd_sc_hd__clkbuf_1 _16835_ (.A(_08808_),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _16836_ (.A0(net9245),
    .A1(\matmul0.sin[6] ),
    .S(net3366),
    .X(_08809_));
 sky130_fd_sc_hd__clkbuf_1 _16837_ (.A(_08809_),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _16838_ (.A0(net6424),
    .A1(\matmul0.sin[7] ),
    .S(net3366),
    .X(_08810_));
 sky130_fd_sc_hd__clkbuf_1 _16839_ (.A(_08810_),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _16840_ (.A0(net6423),
    .A1(\matmul0.sin[8] ),
    .S(net3366),
    .X(_08811_));
 sky130_fd_sc_hd__clkbuf_1 _16841_ (.A(_08811_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _16842_ (.A0(\cordic0.sin[9] ),
    .A1(\matmul0.sin[9] ),
    .S(net3366),
    .X(_08812_));
 sky130_fd_sc_hd__clkbuf_1 _16843_ (.A(_08812_),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _16844_ (.A0(net6422),
    .A1(\matmul0.sin[10] ),
    .S(net3365),
    .X(_08813_));
 sky130_fd_sc_hd__clkbuf_1 _16845_ (.A(_08813_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _16846_ (.A0(net6421),
    .A1(\matmul0.sin[11] ),
    .S(net4287),
    .X(_08814_));
 sky130_fd_sc_hd__clkbuf_1 _16847_ (.A(_08814_),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _16848_ (.A0(\cordic0.sin[12] ),
    .A1(\matmul0.sin[12] ),
    .S(net4287),
    .X(_08815_));
 sky130_fd_sc_hd__clkbuf_1 _16849_ (.A(_08815_),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _16850_ (.A0(\cordic0.sin[13] ),
    .A1(\matmul0.sin[13] ),
    .S(net4287),
    .X(_08816_));
 sky130_fd_sc_hd__clkbuf_1 _16851_ (.A(_08816_),
    .X(_00323_));
 sky130_fd_sc_hd__and2_1 _16852_ (.A(net6457),
    .B(net3668),
    .X(_08817_));
 sky130_fd_sc_hd__clkbuf_1 _16853_ (.A(_08817_),
    .X(_08818_));
 sky130_fd_sc_hd__buf_1 _16854_ (.A(net2196),
    .X(_08819_));
 sky130_fd_sc_hd__mux2_1 _16855_ (.A0(net6082),
    .A1(net6055),
    .S(net6501),
    .X(_08820_));
 sky130_fd_sc_hd__mux2_1 _16856_ (.A0(net6092),
    .A1(net6061),
    .S(net6501),
    .X(_08821_));
 sky130_fd_sc_hd__mux2_1 _16857_ (.A0(net6254),
    .A1(net6195),
    .S(net6498),
    .X(_08822_));
 sky130_fd_sc_hd__mux2_1 _16858_ (.A0(net6277),
    .A1(net6216),
    .S(net6498),
    .X(_08823_));
 sky130_fd_sc_hd__inv_2 _16859_ (.A(net6525),
    .Y(_08824_));
 sky130_fd_sc_hd__inv_2 _16860_ (.A(net6471),
    .Y(_08825_));
 sky130_fd_sc_hd__mux4_1 _16861_ (.A0(_08820_),
    .A1(_08821_),
    .A2(_08822_),
    .A3(_08823_),
    .S0(net4062),
    .S1(_08825_),
    .X(_08826_));
 sky130_fd_sc_hd__mux2_1 _16862_ (.A0(net6167),
    .A1(net6123),
    .S(net6501),
    .X(_08827_));
 sky130_fd_sc_hd__mux2_1 _16863_ (.A0(net6172),
    .A1(net6133),
    .S(net6504),
    .X(_08828_));
 sky130_fd_sc_hd__mux2_1 _16864_ (.A0(_08827_),
    .A1(_08828_),
    .S(net4062),
    .X(_08829_));
 sky130_fd_sc_hd__mux4_1 _16865_ (.A0(net6363),
    .A1(net6344),
    .A2(net6325),
    .A3(net6309),
    .S0(net6518),
    .S1(net6498),
    .X(_08830_));
 sky130_fd_sc_hd__mux2_1 _16866_ (.A0(_08829_),
    .A1(net4061),
    .S(_08825_),
    .X(_08831_));
 sky130_fd_sc_hd__inv_2 _16867_ (.A(net6483),
    .Y(_08832_));
 sky130_fd_sc_hd__mux2_1 _16868_ (.A0(net3364),
    .A1(_08831_),
    .S(net4059),
    .X(_08833_));
 sky130_fd_sc_hd__mux2_1 _16869_ (.A0(net6020),
    .A1(net5997),
    .S(net6523),
    .X(_08834_));
 sky130_fd_sc_hd__or2_1 _16870_ (.A(net6495),
    .B(net6477),
    .X(_08835_));
 sky130_fd_sc_hd__nor2_2 _16871_ (.A(net6468),
    .B(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__mux2_1 _16872_ (.A0(net5992),
    .A1(net4057),
    .S(_08836_),
    .X(_08837_));
 sky130_fd_sc_hd__mux2_1 _16873_ (.A0(net2189),
    .A1(_08837_),
    .S(net6460),
    .X(_08838_));
 sky130_fd_sc_hd__o21ai_1 _16874_ (.A1(net1829),
    .A2(net1828),
    .B1(net8069),
    .Y(_08839_));
 sky130_fd_sc_hd__nor2_1 _16875_ (.A(net7134),
    .B(net1551),
    .Y(_08840_));
 sky130_fd_sc_hd__a22o_1 _16876_ (.A1(net7134),
    .A2(_08839_),
    .B1(_08840_),
    .B2(net1828),
    .X(_00324_));
 sky130_fd_sc_hd__clkbuf_1 _16877_ (.A(net2932),
    .X(_08841_));
 sky130_fd_sc_hd__mux2_1 _16878_ (.A0(net6061),
    .A1(net6019),
    .S(net6501),
    .X(_08842_));
 sky130_fd_sc_hd__mux2_1 _16879_ (.A0(_08820_),
    .A1(_08842_),
    .S(net6525),
    .X(_08843_));
 sky130_fd_sc_hd__mux2_1 _16880_ (.A0(net6216),
    .A1(net6172),
    .S(net6504),
    .X(_08844_));
 sky130_fd_sc_hd__mux2_1 _16881_ (.A0(_08822_),
    .A1(_08844_),
    .S(net6519),
    .X(_08845_));
 sky130_fd_sc_hd__mux2_1 _16882_ (.A0(net6133),
    .A1(net6092),
    .S(net6504),
    .X(_08846_));
 sky130_fd_sc_hd__mux2_1 _16883_ (.A0(_08827_),
    .A1(_08846_),
    .S(net6525),
    .X(_08847_));
 sky130_fd_sc_hd__mux4_1 _16884_ (.A0(net6344),
    .A1(net6325),
    .A2(net6309),
    .A3(net6277),
    .S0(net6518),
    .S1(net6498),
    .X(_08848_));
 sky130_fd_sc_hd__mux4_1 _16885_ (.A0(net3362),
    .A1(_08845_),
    .A2(_08847_),
    .A3(net4056),
    .S0(_08825_),
    .S1(net4059),
    .X(_08849_));
 sky130_fd_sc_hd__inv_2 _16886_ (.A(net6462),
    .Y(_08850_));
 sky130_fd_sc_hd__mux2_1 _16887_ (.A0(net5989),
    .A1(net2612),
    .S(_08850_),
    .X(_08851_));
 sky130_fd_sc_hd__or2b_1 _16888_ (.A(net6368),
    .B_N(net6390),
    .X(_08852_));
 sky130_fd_sc_hd__or2b_1 _16889_ (.A(\cordic0.slte0.opA[14] ),
    .B_N(net6393),
    .X(_08853_));
 sky130_fd_sc_hd__and2b_1 _16890_ (.A_N(net6390),
    .B(net6368),
    .X(_08854_));
 sky130_fd_sc_hd__a21oi_1 _16891_ (.A1(_08852_),
    .A2(_08853_),
    .B1(_08854_),
    .Y(_08855_));
 sky130_fd_sc_hd__or2_1 _16892_ (.A(\cordic0.slte0.opA[17] ),
    .B(_08855_),
    .X(_08856_));
 sky130_fd_sc_hd__inv_2 _16893_ (.A(net6370),
    .Y(_08857_));
 sky130_fd_sc_hd__nor2_1 _16894_ (.A(net6399),
    .B(_08857_),
    .Y(_08858_));
 sky130_fd_sc_hd__o21ba_1 _16895_ (.A1(net6369),
    .A2(_08858_),
    .B1_N(net6396),
    .X(_08859_));
 sky130_fd_sc_hd__a21oi_1 _16896_ (.A1(net6369),
    .A2(_08858_),
    .B1(_08859_),
    .Y(_08860_));
 sky130_fd_sc_hd__and2b_1 _16897_ (.A_N(net6402),
    .B(net6372),
    .X(_08861_));
 sky130_fd_sc_hd__inv_2 _16898_ (.A(\cordic0.slte0.opB[11] ),
    .Y(_08862_));
 sky130_fd_sc_hd__a21o_1 _16899_ (.A1(net6371),
    .A2(_08861_),
    .B1(_08862_),
    .X(_08863_));
 sky130_fd_sc_hd__o21ai_1 _16900_ (.A1(net6371),
    .A2(_08861_),
    .B1(_08863_),
    .Y(_08864_));
 sky130_fd_sc_hd__inv_2 _16901_ (.A(net6372),
    .Y(_08865_));
 sky130_fd_sc_hd__or2b_1 _16902_ (.A(\cordic0.slte0.opA[8] ),
    .B_N(net6407),
    .X(_08866_));
 sky130_fd_sc_hd__o21bai_1 _16903_ (.A1(\cordic0.slte0.opA[9] ),
    .A2(_08866_),
    .B1_N(net6404),
    .Y(_08867_));
 sky130_fd_sc_hd__nand2_1 _16904_ (.A(\cordic0.slte0.opA[9] ),
    .B(_08866_),
    .Y(_08868_));
 sky130_fd_sc_hd__nor2_1 _16905_ (.A(_08862_),
    .B(net6371),
    .Y(_08869_));
 sky130_fd_sc_hd__a221o_1 _16906_ (.A1(net6402),
    .A2(_08865_),
    .B1(_08867_),
    .B2(_08868_),
    .C1(_08869_),
    .X(_08870_));
 sky130_fd_sc_hd__or2b_1 _16907_ (.A(\cordic0.slte0.opA[6] ),
    .B_N(net6413),
    .X(_08871_));
 sky130_fd_sc_hd__nor2_1 _16908_ (.A(net6373),
    .B(_08871_),
    .Y(_08872_));
 sky130_fd_sc_hd__nand2_1 _16909_ (.A(net6373),
    .B(_08871_),
    .Y(_08873_));
 sky130_fd_sc_hd__xor2_1 _16910_ (.A(net6407),
    .B(\cordic0.slte0.opA[8] ),
    .X(_08874_));
 sky130_fd_sc_hd__xor2_1 _16911_ (.A(net6404),
    .B(\cordic0.slte0.opA[9] ),
    .X(_08875_));
 sky130_fd_sc_hd__xor2_1 _16912_ (.A(net6402),
    .B(net6372),
    .X(_08876_));
 sky130_fd_sc_hd__a2111oi_1 _16913_ (.A1(_08862_),
    .A2(net6371),
    .B1(_08874_),
    .C1(_08875_),
    .D1(_08876_),
    .Y(_08877_));
 sky130_fd_sc_hd__o211a_1 _16914_ (.A1(net6410),
    .A2(_08872_),
    .B1(_08873_),
    .C1(net9247),
    .X(_08878_));
 sky130_fd_sc_hd__or2b_1 _16915_ (.A(net6370),
    .B_N(net6399),
    .X(_08879_));
 sky130_fd_sc_hd__o21bai_1 _16916_ (.A1(net6369),
    .A2(_08879_),
    .B1_N(net6396),
    .Y(_08880_));
 sky130_fd_sc_hd__nand2_1 _16917_ (.A(net6369),
    .B(_08879_),
    .Y(_08881_));
 sky130_fd_sc_hd__a211o_1 _16918_ (.A1(_08880_),
    .A2(_08881_),
    .B1(\cordic0.slte0.opA[17] ),
    .C1(_08855_),
    .X(_08882_));
 sky130_fd_sc_hd__a211o_1 _16919_ (.A1(_08864_),
    .A2(_08870_),
    .B1(_08878_),
    .C1(net2611),
    .X(_08883_));
 sky130_fd_sc_hd__inv_2 _16920_ (.A(\cordic0.slte0.opA[4] ),
    .Y(_08884_));
 sky130_fd_sc_hd__inv_2 _16921_ (.A(\cordic0.slte0.opA[3] ),
    .Y(_08885_));
 sky130_fd_sc_hd__o21ai_1 _16922_ (.A1(\cordic0.slte0.opA[1] ),
    .A2(\cordic0.slte0.opA[0] ),
    .B1(\cordic0.slte0.opA[2] ),
    .Y(_08886_));
 sky130_fd_sc_hd__or3_1 _16923_ (.A(\cordic0.slte0.opA[2] ),
    .B(\cordic0.slte0.opA[1] ),
    .C(\cordic0.slte0.opA[0] ),
    .X(_08887_));
 sky130_fd_sc_hd__a21bo_1 _16924_ (.A1(net6420),
    .A2(_08886_),
    .B1_N(_08887_),
    .X(_08888_));
 sky130_fd_sc_hd__o221a_1 _16925_ (.A1(net6418),
    .A2(_08884_),
    .B1(net6419),
    .B2(_08885_),
    .C1(_08888_),
    .X(_08889_));
 sky130_fd_sc_hd__inv_2 _16926_ (.A(\cordic0.slte0.opA[5] ),
    .Y(_08890_));
 sky130_fd_sc_hd__and2b_1 _16927_ (.A_N(\cordic0.slte0.opA[3] ),
    .B(net6419),
    .X(_08891_));
 sky130_fd_sc_hd__a21o_1 _16928_ (.A1(net6418),
    .A2(_08891_),
    .B1(_08884_),
    .X(_08892_));
 sky130_fd_sc_hd__or2_1 _16929_ (.A(net6418),
    .B(_08891_),
    .X(_08893_));
 sky130_fd_sc_hd__a22o_1 _16930_ (.A1(net6416),
    .A2(_08890_),
    .B1(_08892_),
    .B2(_08893_),
    .X(_08894_));
 sky130_fd_sc_hd__xnor2_1 _16931_ (.A(net6410),
    .B(net6373),
    .Y(_08895_));
 sky130_fd_sc_hd__inv_2 _16932_ (.A(net6374),
    .Y(_08896_));
 sky130_fd_sc_hd__or2_1 _16933_ (.A(net6413),
    .B(_08896_),
    .X(_08897_));
 sky130_fd_sc_hd__o211a_1 _16934_ (.A1(net6416),
    .A2(_08890_),
    .B1(_08871_),
    .C1(_08897_),
    .X(_08898_));
 sky130_fd_sc_hd__o2111a_1 _16935_ (.A1(_08889_),
    .A2(_08894_),
    .B1(_08895_),
    .C1(_08898_),
    .D1(net3360),
    .X(_08899_));
 sky130_fd_sc_hd__inv_2 _16936_ (.A(\cordic0.slte0.opA[16] ),
    .Y(_08900_));
 sky130_fd_sc_hd__and2b_1 _16937_ (.A_N(net6393),
    .B(\cordic0.slte0.opA[14] ),
    .X(_08901_));
 sky130_fd_sc_hd__o21ai_1 _16938_ (.A1(_08854_),
    .A2(_08901_),
    .B1(_08852_),
    .Y(_08902_));
 sky130_fd_sc_hd__a21o_1 _16939_ (.A1(net4054),
    .A2(_08902_),
    .B1(\cordic0.slte0.opA[17] ),
    .X(_08903_));
 sky130_fd_sc_hd__o221a_1 _16940_ (.A1(_08856_),
    .A2(_08860_),
    .B1(net2176),
    .B2(net2174),
    .C1(_08903_),
    .X(_08904_));
 sky130_fd_sc_hd__clkbuf_1 _16941_ (.A(net1827),
    .X(_08905_));
 sky130_fd_sc_hd__xnor2_1 _16942_ (.A(net7138),
    .B(net1506),
    .Y(_08906_));
 sky130_fd_sc_hd__nand2_1 _16943_ (.A(net1828),
    .B(_08906_),
    .Y(_08907_));
 sky130_fd_sc_hd__xor2_1 _16944_ (.A(net2177),
    .B(_08907_),
    .X(_08908_));
 sky130_fd_sc_hd__buf_1 _16945_ (.A(net4241),
    .X(_08909_));
 sky130_fd_sc_hd__a21o_1 _16946_ (.A1(net2180),
    .A2(_08908_),
    .B1(net3351),
    .X(_08910_));
 sky130_fd_sc_hd__buf_1 _16947_ (.A(net2284),
    .X(_08911_));
 sky130_fd_sc_hd__or3_1 _16948_ (.A(net7125),
    .B(net1818),
    .C(_08908_),
    .X(_08912_));
 sky130_fd_sc_hd__a21bo_1 _16949_ (.A1(net7125),
    .A2(_08910_),
    .B1_N(_08912_),
    .X(_00325_));
 sky130_fd_sc_hd__inv_2 _16950_ (.A(net7106),
    .Y(_08913_));
 sky130_fd_sc_hd__buf_1 _16951_ (.A(_08913_),
    .X(_08914_));
 sky130_fd_sc_hd__nor2_1 _16952_ (.A(net4246),
    .B(net2197),
    .Y(_08915_));
 sky130_fd_sc_hd__buf_1 _16953_ (.A(net1814),
    .X(_08916_));
 sky130_fd_sc_hd__clkbuf_1 _16954_ (.A(net1495),
    .X(_08917_));
 sky130_fd_sc_hd__o221ai_1 _16955_ (.A1(_08856_),
    .A2(_08860_),
    .B1(net2176),
    .B2(net2174),
    .C1(_08903_),
    .Y(_08918_));
 sky130_fd_sc_hd__nand2_1 _16956_ (.A(_08838_),
    .B(net1808),
    .Y(_08919_));
 sky130_fd_sc_hd__o21bai_1 _16957_ (.A1(net2177),
    .A2(net1825),
    .B1_N(net7138),
    .Y(_08920_));
 sky130_fd_sc_hd__xnor2_1 _16958_ (.A(net2177),
    .B(net1825),
    .Y(_08921_));
 sky130_fd_sc_hd__a22o_1 _16959_ (.A1(net7129),
    .A2(_08920_),
    .B1(_08921_),
    .B2(net7147),
    .X(_08922_));
 sky130_fd_sc_hd__a32o_1 _16960_ (.A1(net7129),
    .A2(net2177),
    .A3(_08919_),
    .B1(_08922_),
    .B2(_08838_),
    .X(_08923_));
 sky130_fd_sc_hd__clkbuf_2 _16961_ (.A(_08850_),
    .X(_08924_));
 sky130_fd_sc_hd__buf_1 _16962_ (.A(_08924_),
    .X(_08925_));
 sky130_fd_sc_hd__mux2_1 _16963_ (.A0(net6055),
    .A1(net5996),
    .S(net6501),
    .X(_08926_));
 sky130_fd_sc_hd__mux2_1 _16964_ (.A0(_08842_),
    .A1(_08926_),
    .S(net6522),
    .X(_08927_));
 sky130_fd_sc_hd__mux2_1 _16965_ (.A0(net6195),
    .A1(net6167),
    .S(net6504),
    .X(_08928_));
 sky130_fd_sc_hd__mux2_1 _16966_ (.A0(_08844_),
    .A1(_08928_),
    .S(net6519),
    .X(_08929_));
 sky130_fd_sc_hd__mux2_1 _16967_ (.A0(net6123),
    .A1(net6082),
    .S(net6501),
    .X(_08930_));
 sky130_fd_sc_hd__mux2_1 _16968_ (.A0(_08846_),
    .A1(_08930_),
    .S(net6525),
    .X(_08931_));
 sky130_fd_sc_hd__mux4_1 _16969_ (.A0(net6325),
    .A1(net6309),
    .A2(net6277),
    .A3(net6254),
    .S0(net6518),
    .S1(net6498),
    .X(_08932_));
 sky130_fd_sc_hd__mux4_1 _16970_ (.A0(_08927_),
    .A1(_08929_),
    .A2(_08931_),
    .A3(net4053),
    .S0(_08825_),
    .S1(net4059),
    .X(_08933_));
 sky130_fd_sc_hd__o21a_1 _16971_ (.A1(_08838_),
    .A2(net2612),
    .B1(net1808),
    .X(_08934_));
 sky130_fd_sc_hd__xnor2_1 _16972_ (.A(net2606),
    .B(_08934_),
    .Y(_08935_));
 sky130_fd_sc_hd__nand2_1 _16973_ (.A(_08925_),
    .B(_08935_),
    .Y(_08936_));
 sky130_fd_sc_hd__nor2_1 _16974_ (.A(net5989),
    .B(_08919_),
    .Y(_08937_));
 sky130_fd_sc_hd__a211o_1 _16975_ (.A1(net5989),
    .A2(net1825),
    .B1(_08937_),
    .C1(_08924_),
    .X(_08938_));
 sky130_fd_sc_hd__and2_1 _16976_ (.A(_08936_),
    .B(_08938_),
    .X(_08939_));
 sky130_fd_sc_hd__xor2_1 _16977_ (.A(_08923_),
    .B(_08939_),
    .X(_08940_));
 sky130_fd_sc_hd__o21a_1 _16978_ (.A1(net1918),
    .A2(net878),
    .B1(net8069),
    .X(_08941_));
 sky130_fd_sc_hd__nor2_1 _16979_ (.A(net3349),
    .B(_08941_),
    .Y(_08942_));
 sky130_fd_sc_hd__a31o_1 _16980_ (.A1(net3349),
    .A2(net1232),
    .A3(net878),
    .B1(_08942_),
    .X(_00326_));
 sky130_fd_sc_hd__and3_1 _16981_ (.A(net6493),
    .B(net6475),
    .C(net6467),
    .X(_08943_));
 sky130_fd_sc_hd__a21o_1 _16982_ (.A1(net6520),
    .A2(net4052),
    .B1(net6460),
    .X(_08944_));
 sky130_fd_sc_hd__and2b_1 _16983_ (.A_N(net6502),
    .B(net6522),
    .X(_08945_));
 sky130_fd_sc_hd__a22o_1 _16984_ (.A1(_08824_),
    .A2(_08926_),
    .B1(net4051),
    .B2(net6019),
    .X(_08946_));
 sky130_fd_sc_hd__mux2_1 _16985_ (.A0(_08828_),
    .A1(_08928_),
    .S(net4062),
    .X(_08947_));
 sky130_fd_sc_hd__mux2_1 _16986_ (.A0(_08821_),
    .A1(_08930_),
    .S(net4062),
    .X(_08948_));
 sky130_fd_sc_hd__mux4_1 _16987_ (.A0(net6309),
    .A1(net6254),
    .A2(net6277),
    .A3(net6216),
    .S0(net6498),
    .S1(net6518),
    .X(_08949_));
 sky130_fd_sc_hd__mux4_1 _16988_ (.A0(_08946_),
    .A1(_08947_),
    .A2(_08948_),
    .A3(net4049),
    .S0(_08825_),
    .S1(net4059),
    .X(_08950_));
 sky130_fd_sc_hd__a22o_1 _16989_ (.A1(net5989),
    .A2(_08944_),
    .B1(net2605),
    .B2(_08924_),
    .X(_08951_));
 sky130_fd_sc_hd__buf_1 _16990_ (.A(net1809),
    .X(_08952_));
 sky130_fd_sc_hd__or2_1 _16991_ (.A(net2612),
    .B(net2606),
    .X(_08953_));
 sky130_fd_sc_hd__inv_2 _16992_ (.A(net5995),
    .Y(_08954_));
 sky130_fd_sc_hd__nand2_1 _16993_ (.A(net6461),
    .B(net4048),
    .Y(_08955_));
 sky130_fd_sc_hd__a21o_1 _16994_ (.A1(_08836_),
    .A2(net4057),
    .B1(_08955_),
    .X(_08956_));
 sky130_fd_sc_hd__o31a_1 _16995_ (.A1(net6460),
    .A2(net2189),
    .A3(_08953_),
    .B1(_08956_),
    .X(_08957_));
 sky130_fd_sc_hd__nand2_1 _16996_ (.A(_08952_),
    .B(net1806),
    .Y(_08958_));
 sky130_fd_sc_hd__xnor2_1 _16997_ (.A(net2173),
    .B(_08958_),
    .Y(_08959_));
 sky130_fd_sc_hd__a21o_1 _16998_ (.A1(_08936_),
    .A2(_08938_),
    .B1(_08923_),
    .X(_08960_));
 sky130_fd_sc_hd__a31o_1 _16999_ (.A1(_08923_),
    .A2(_08936_),
    .A3(_08938_),
    .B1(net7113),
    .X(_08961_));
 sky130_fd_sc_hd__nand2_1 _17000_ (.A(_08960_),
    .B(_08961_),
    .Y(_08962_));
 sky130_fd_sc_hd__xnor2_1 _17001_ (.A(_08959_),
    .B(_08962_),
    .Y(_08963_));
 sky130_fd_sc_hd__o21ai_1 _17002_ (.A1(net1833),
    .A2(_08963_),
    .B1(net8042),
    .Y(_08964_));
 sky130_fd_sc_hd__nor2_1 _17003_ (.A(net7080),
    .B(net1552),
    .Y(_08965_));
 sky130_fd_sc_hd__a22o_1 _17004_ (.A1(net7080),
    .A2(_08964_),
    .B1(_08965_),
    .B2(_08963_),
    .X(_00327_));
 sky130_fd_sc_hd__inv_2 _17005_ (.A(net7065),
    .Y(_08966_));
 sky130_fd_sc_hd__buf_1 _17006_ (.A(net4044),
    .X(_08967_));
 sky130_fd_sc_hd__or2_1 _17007_ (.A(net6480),
    .B(net3364),
    .X(_08968_));
 sky130_fd_sc_hd__buf_1 _17008_ (.A(_08825_),
    .X(_08969_));
 sky130_fd_sc_hd__nor2_1 _17009_ (.A(net6500),
    .B(net3335),
    .Y(_08970_));
 sky130_fd_sc_hd__clkbuf_2 _17010_ (.A(net4060),
    .X(_08971_));
 sky130_fd_sc_hd__a221o_1 _17011_ (.A1(net3335),
    .A2(net3363),
    .B1(net4057),
    .B2(_08970_),
    .C1(_08971_),
    .X(_08972_));
 sky130_fd_sc_hd__or2_1 _17012_ (.A(net6465),
    .B(net4052),
    .X(_08973_));
 sky130_fd_sc_hd__a32o_1 _17013_ (.A1(net3345),
    .A2(_08968_),
    .A3(_08972_),
    .B1(_08973_),
    .B2(net5993),
    .X(_08974_));
 sky130_fd_sc_hd__or2_1 _17014_ (.A(net2173),
    .B(net1806),
    .X(_08975_));
 sky130_fd_sc_hd__and2_1 _17015_ (.A(net1807),
    .B(net1483),
    .X(_08976_));
 sky130_fd_sc_hd__xnor2_2 _17016_ (.A(net1804),
    .B(_08976_),
    .Y(_08977_));
 sky130_fd_sc_hd__a22o_1 _17017_ (.A1(net7086),
    .A2(_08959_),
    .B1(_08961_),
    .B2(_08960_),
    .X(_08978_));
 sky130_fd_sc_hd__or2_1 _17018_ (.A(net7086),
    .B(_08959_),
    .X(_08979_));
 sky130_fd_sc_hd__nand2_2 _17019_ (.A(_08978_),
    .B(_08979_),
    .Y(_08980_));
 sky130_fd_sc_hd__xor2_1 _17020_ (.A(_08977_),
    .B(_08980_),
    .X(_08981_));
 sky130_fd_sc_hd__o21a_1 _17021_ (.A1(net1917),
    .A2(_08981_),
    .B1(net8043),
    .X(_08982_));
 sky130_fd_sc_hd__nor2_1 _17022_ (.A(net7053),
    .B(net1553),
    .Y(_08983_));
 sky130_fd_sc_hd__a2bb2o_1 _17023_ (.A1_N(net3336),
    .A2_N(_08982_),
    .B1(_08983_),
    .B2(_08981_),
    .X(_00328_));
 sky130_fd_sc_hd__inv_2 _17024_ (.A(net7029),
    .Y(_08984_));
 sky130_fd_sc_hd__buf_1 _17025_ (.A(_08984_),
    .X(_08985_));
 sky130_fd_sc_hd__a31o_1 _17026_ (.A1(net6478),
    .A2(net6473),
    .A3(_06503_),
    .B1(net6460),
    .X(_08986_));
 sky130_fd_sc_hd__nor2_1 _17027_ (.A(net4048),
    .B(net4237),
    .Y(_08987_));
 sky130_fd_sc_hd__mux4_1 _17028_ (.A0(net3362),
    .A1(_08845_),
    .A2(_08987_),
    .A3(_08847_),
    .S0(net3335),
    .S1(net6480),
    .X(_08988_));
 sky130_fd_sc_hd__a22o_1 _17029_ (.A1(net5989),
    .A2(_08986_),
    .B1(net2603),
    .B2(_08924_),
    .X(_08989_));
 sky130_fd_sc_hd__buf_1 _17030_ (.A(net1809),
    .X(_08990_));
 sky130_fd_sc_hd__buf_1 _17031_ (.A(net1480),
    .X(_08991_));
 sky130_fd_sc_hd__buf_1 _17032_ (.A(net1225),
    .X(_08992_));
 sky130_fd_sc_hd__buf_1 _17033_ (.A(net1077),
    .X(_08993_));
 sky130_fd_sc_hd__inv_2 _17034_ (.A(_08980_),
    .Y(_08994_));
 sky130_fd_sc_hd__nor2_1 _17035_ (.A(_08976_),
    .B(_08980_),
    .Y(_08995_));
 sky130_fd_sc_hd__or3_1 _17036_ (.A(net3336),
    .B(net1804),
    .C(_08995_),
    .X(_08996_));
 sky130_fd_sc_hd__nand2_1 _17037_ (.A(net7053),
    .B(net967),
    .Y(_08997_));
 sky130_fd_sc_hd__mux2_1 _17038_ (.A0(net7053),
    .A1(_08997_),
    .S(net1804),
    .X(_08998_));
 sky130_fd_sc_hd__a21o_1 _17039_ (.A1(net1483),
    .A2(_08980_),
    .B1(_08998_),
    .X(_08999_));
 sky130_fd_sc_hd__o311a_1 _17040_ (.A1(net7057),
    .A2(net967),
    .A3(_08994_),
    .B1(_08996_),
    .C1(_08999_),
    .X(_09000_));
 sky130_fd_sc_hd__xor2_1 _17041_ (.A(net2171),
    .B(_09000_),
    .X(_09001_));
 sky130_fd_sc_hd__o21a_1 _17042_ (.A1(net1831),
    .A2(_09001_),
    .B1(net8043),
    .X(_09002_));
 sky130_fd_sc_hd__nor2_1 _17043_ (.A(net3328),
    .B(_09002_),
    .Y(_09003_));
 sky130_fd_sc_hd__a31o_1 _17044_ (.A1(net3328),
    .A2(net1231),
    .A3(_09001_),
    .B1(_09003_),
    .X(_00329_));
 sky130_fd_sc_hd__buf_1 _17045_ (.A(net3334),
    .X(_09004_));
 sky130_fd_sc_hd__or2_1 _17046_ (.A(net6474),
    .B(net6462),
    .X(_09005_));
 sky130_fd_sc_hd__buf_1 _17047_ (.A(_09005_),
    .X(_09006_));
 sky130_fd_sc_hd__o22a_1 _17048_ (.A1(net2601),
    .A2(net5993),
    .B1(_08931_),
    .B2(net3326),
    .X(_09007_));
 sky130_fd_sc_hd__or2_1 _17049_ (.A(net6486),
    .B(net6464),
    .X(_09008_));
 sky130_fd_sc_hd__mux2_1 _17050_ (.A0(_08927_),
    .A1(_08929_),
    .S(_08969_),
    .X(_09009_));
 sky130_fd_sc_hd__o221a_1 _17051_ (.A1(_08971_),
    .A2(_09007_),
    .B1(_09008_),
    .B2(_09009_),
    .C1(_08955_),
    .X(_09010_));
 sky130_fd_sc_hd__o31a_1 _17052_ (.A1(net1805),
    .A2(_08975_),
    .A3(net2172),
    .B1(net1807),
    .X(_09011_));
 sky130_fd_sc_hd__xor2_2 _17053_ (.A(net1802),
    .B(_09011_),
    .X(_09012_));
 sky130_fd_sc_hd__o21ai_1 _17054_ (.A1(net1804),
    .A2(net1483),
    .B1(_08952_),
    .Y(_09013_));
 sky130_fd_sc_hd__xnor2_2 _17055_ (.A(net2171),
    .B(_09013_),
    .Y(_09014_));
 sky130_fd_sc_hd__xnor2_1 _17056_ (.A(net7057),
    .B(_08977_),
    .Y(_09015_));
 sky130_fd_sc_hd__o211a_1 _17057_ (.A1(net7039),
    .A2(_09014_),
    .B1(_09015_),
    .C1(_08994_),
    .X(_09016_));
 sky130_fd_sc_hd__xnor2_1 _17058_ (.A(net1807),
    .B(net2171),
    .Y(_09017_));
 sky130_fd_sc_hd__a21o_1 _17059_ (.A1(net3328),
    .A2(_09017_),
    .B1(net3336),
    .X(_09018_));
 sky130_fd_sc_hd__or2_1 _17060_ (.A(_08977_),
    .B(_09018_),
    .X(_09019_));
 sky130_fd_sc_hd__inv_2 _17061_ (.A(_09019_),
    .Y(_09020_));
 sky130_fd_sc_hd__a211o_1 _17062_ (.A1(net7039),
    .A2(_09014_),
    .B1(_09016_),
    .C1(_09020_),
    .X(_09021_));
 sky130_fd_sc_hd__xnor2_1 _17063_ (.A(_09012_),
    .B(_09021_),
    .Y(_09022_));
 sky130_fd_sc_hd__buf_1 _17064_ (.A(net4246),
    .X(_09023_));
 sky130_fd_sc_hd__a21o_1 _17065_ (.A1(net2179),
    .A2(_09022_),
    .B1(net3320),
    .X(_09024_));
 sky130_fd_sc_hd__nor2_1 _17066_ (.A(net1918),
    .B(_09022_),
    .Y(_09025_));
 sky130_fd_sc_hd__inv_2 _17067_ (.A(net7004),
    .Y(_09026_));
 sky130_fd_sc_hd__mux2_1 _17068_ (.A0(_09024_),
    .A1(_09025_),
    .S(_09026_),
    .X(_09027_));
 sky130_fd_sc_hd__clkbuf_1 _17069_ (.A(_09027_),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _17070_ (.A0(_08946_),
    .A1(_08947_),
    .S(net2601),
    .X(_09028_));
 sky130_fd_sc_hd__nor2_1 _17071_ (.A(net3332),
    .B(net6474),
    .Y(_09029_));
 sky130_fd_sc_hd__a22o_1 _17072_ (.A1(net3332),
    .A2(_09028_),
    .B1(net3342),
    .B2(_09029_),
    .X(_09030_));
 sky130_fd_sc_hd__buf_1 _17073_ (.A(net4062),
    .X(_09031_));
 sky130_fd_sc_hd__inv_2 _17074_ (.A(net6494),
    .Y(_09032_));
 sky130_fd_sc_hd__nor2_1 _17075_ (.A(net3313),
    .B(net4040),
    .Y(_09033_));
 sky130_fd_sc_hd__o21ai_1 _17076_ (.A1(net6485),
    .A2(net2598),
    .B1(net6473),
    .Y(_09034_));
 sky130_fd_sc_hd__nand2_1 _17077_ (.A(net2609),
    .B(_09034_),
    .Y(_09035_));
 sky130_fd_sc_hd__a22o_1 _17078_ (.A1(net2609),
    .A2(_09030_),
    .B1(_09035_),
    .B2(net5990),
    .X(_09036_));
 sky130_fd_sc_hd__or4_1 _17079_ (.A(net1805),
    .B(_08975_),
    .C(net2172),
    .D(net1802),
    .X(_09037_));
 sky130_fd_sc_hd__nand2_1 _17080_ (.A(net1221),
    .B(_09037_),
    .Y(_09038_));
 sky130_fd_sc_hd__xnor2_2 _17081_ (.A(net1478),
    .B(_09038_),
    .Y(_09039_));
 sky130_fd_sc_hd__o21bai_1 _17082_ (.A1(_08977_),
    .A2(_09018_),
    .B1_N(_09014_),
    .Y(_09040_));
 sky130_fd_sc_hd__nand2_1 _17083_ (.A(net7008),
    .B(_09012_),
    .Y(_09041_));
 sky130_fd_sc_hd__nand2b_1 _17084_ (.A_N(_09040_),
    .B(_09041_),
    .Y(_09042_));
 sky130_fd_sc_hd__nand3_1 _17085_ (.A(net3328),
    .B(_09019_),
    .C(_09041_),
    .Y(_09043_));
 sky130_fd_sc_hd__a32o_1 _17086_ (.A1(_08978_),
    .A2(_08979_),
    .A3(_09015_),
    .B1(_09042_),
    .B2(_09043_),
    .X(_09044_));
 sky130_fd_sc_hd__or3b_1 _17087_ (.A(net7039),
    .B(_09014_),
    .C_N(_09041_),
    .X(_09045_));
 sky130_fd_sc_hd__o211a_1 _17088_ (.A1(net7008),
    .A2(_09012_),
    .B1(_09044_),
    .C1(_09045_),
    .X(_09046_));
 sky130_fd_sc_hd__xor2_1 _17089_ (.A(_09039_),
    .B(net772),
    .X(_09047_));
 sky130_fd_sc_hd__o21ai_1 _17090_ (.A1(net1829),
    .A2(_09047_),
    .B1(net8050),
    .Y(_09048_));
 sky130_fd_sc_hd__nor2_1 _17091_ (.A(net6981),
    .B(net1551),
    .Y(_09049_));
 sky130_fd_sc_hd__a22o_1 _17092_ (.A1(net6981),
    .A2(_09048_),
    .B1(_09049_),
    .B2(_09047_),
    .X(_00331_));
 sky130_fd_sc_hd__inv_2 _17093_ (.A(net6974),
    .Y(_09050_));
 sky130_fd_sc_hd__clkbuf_1 _17094_ (.A(_09050_),
    .X(_09051_));
 sky130_fd_sc_hd__mux2_1 _17095_ (.A0(_08820_),
    .A1(_08821_),
    .S(_09031_),
    .X(_09052_));
 sky130_fd_sc_hd__mux2_1 _17096_ (.A0(net2595),
    .A1(net3363),
    .S(_08971_),
    .X(_09053_));
 sky130_fd_sc_hd__nor2_1 _17097_ (.A(net6495),
    .B(net6477),
    .Y(_09054_));
 sky130_fd_sc_hd__nand2_1 _17098_ (.A(net2609),
    .B(net4038),
    .Y(_09055_));
 sky130_fd_sc_hd__o22a_1 _17099_ (.A1(net5992),
    .A2(net4038),
    .B1(net4057),
    .B2(_09055_),
    .X(_09056_));
 sky130_fd_sc_hd__o221a_1 _17100_ (.A1(_09053_),
    .A2(net3326),
    .B1(_09056_),
    .B2(net2602),
    .C1(_08955_),
    .X(_09057_));
 sky130_fd_sc_hd__nor2_1 _17101_ (.A(net1478),
    .B(_09037_),
    .Y(_09058_));
 sky130_fd_sc_hd__or2_1 _17102_ (.A(net1505),
    .B(_09058_),
    .X(_09059_));
 sky130_fd_sc_hd__xnor2_1 _17103_ (.A(net1476),
    .B(_09059_),
    .Y(_09060_));
 sky130_fd_sc_hd__a21o_1 _17104_ (.A1(_09039_),
    .A2(net772),
    .B1(net6981),
    .X(_09061_));
 sky130_fd_sc_hd__o21a_1 _17105_ (.A1(_09039_),
    .A2(net772),
    .B1(_09061_),
    .X(_09062_));
 sky130_fd_sc_hd__nor2_1 _17106_ (.A(_09060_),
    .B(_09062_),
    .Y(_09063_));
 sky130_fd_sc_hd__and2_1 _17107_ (.A(_09060_),
    .B(_09062_),
    .X(_09064_));
 sky130_fd_sc_hd__nor2_1 _17108_ (.A(_09063_),
    .B(_09064_),
    .Y(_09065_));
 sky130_fd_sc_hd__o21a_1 _17109_ (.A1(net1818),
    .A2(_09065_),
    .B1(net8049),
    .X(_09066_));
 sky130_fd_sc_hd__nor2_1 _17110_ (.A(net3307),
    .B(_09066_),
    .Y(_09067_));
 sky130_fd_sc_hd__a31o_1 _17111_ (.A1(net3307),
    .A2(net1233),
    .A3(_09065_),
    .B1(_09067_),
    .X(_00332_));
 sky130_fd_sc_hd__buf_1 _17112_ (.A(net1813),
    .X(_09068_));
 sky130_fd_sc_hd__buf_1 _17113_ (.A(net3332),
    .X(_09069_));
 sky130_fd_sc_hd__mux2_1 _17114_ (.A0(net3362),
    .A1(_08847_),
    .S(net2593),
    .X(_09070_));
 sky130_fd_sc_hd__nor2_1 _17115_ (.A(net6470),
    .B(net6462),
    .Y(_09071_));
 sky130_fd_sc_hd__mux2_1 _17116_ (.A0(net5990),
    .A1(net2170),
    .S(_09071_),
    .X(_09072_));
 sky130_fd_sc_hd__inv_2 _17117_ (.A(_09058_),
    .Y(_09073_));
 sky130_fd_sc_hd__o21ai_2 _17118_ (.A1(net1476),
    .A2(_09073_),
    .B1(net1221),
    .Y(_09074_));
 sky130_fd_sc_hd__xnor2_2 _17119_ (.A(_09072_),
    .B(_09074_),
    .Y(_09075_));
 sky130_fd_sc_hd__o21a_1 _17120_ (.A1(_09060_),
    .A2(_09062_),
    .B1(net6961),
    .X(_09076_));
 sky130_fd_sc_hd__or2_1 _17121_ (.A(_09064_),
    .B(_09076_),
    .X(_09077_));
 sky130_fd_sc_hd__xnor2_1 _17122_ (.A(_09075_),
    .B(_09077_),
    .Y(_09078_));
 sky130_fd_sc_hd__a21o_1 _17123_ (.A1(_09068_),
    .A2(_09078_),
    .B1(net3350),
    .X(_09079_));
 sky130_fd_sc_hd__or3_1 _17124_ (.A(net6936),
    .B(net1819),
    .C(_09078_),
    .X(_09080_));
 sky130_fd_sc_hd__a21bo_1 _17125_ (.A1(net6932),
    .A2(_09079_),
    .B1_N(_09080_),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _17126_ (.A0(net3344),
    .A1(_08931_),
    .S(net2593),
    .X(_09081_));
 sky130_fd_sc_hd__buf_1 _17127_ (.A(_09071_),
    .X(_09082_));
 sky130_fd_sc_hd__mux2_1 _17128_ (.A0(net5990),
    .A1(net2169),
    .S(_09082_),
    .X(_09083_));
 sky130_fd_sc_hd__or3_1 _17129_ (.A(net1476),
    .B(_09073_),
    .C(_09072_),
    .X(_09084_));
 sky130_fd_sc_hd__nand2_1 _17130_ (.A(net1221),
    .B(_09084_),
    .Y(_09085_));
 sky130_fd_sc_hd__xnor2_2 _17131_ (.A(_09083_),
    .B(_09085_),
    .Y(_09086_));
 sky130_fd_sc_hd__a21o_1 _17132_ (.A1(_09075_),
    .A2(_09077_),
    .B1(net6932),
    .X(_09087_));
 sky130_fd_sc_hd__o21a_1 _17133_ (.A1(_09075_),
    .A2(_09077_),
    .B1(_09087_),
    .X(_09088_));
 sky130_fd_sc_hd__xnor2_1 _17134_ (.A(_09086_),
    .B(_09088_),
    .Y(_09089_));
 sky130_fd_sc_hd__a21o_1 _17135_ (.A1(net2181),
    .A2(_09089_),
    .B1(net3322),
    .X(_09090_));
 sky130_fd_sc_hd__or3_1 _17136_ (.A(net6914),
    .B(net1819),
    .C(_09089_),
    .X(_09091_));
 sky130_fd_sc_hd__a21bo_1 _17137_ (.A1(net6914),
    .A2(_09090_),
    .B1_N(_09091_),
    .X(_00334_));
 sky130_fd_sc_hd__inv_2 _17138_ (.A(net6906),
    .Y(_09092_));
 sky130_fd_sc_hd__clkbuf_1 _17139_ (.A(_09092_),
    .X(_09093_));
 sky130_fd_sc_hd__a22o_1 _17140_ (.A1(net5988),
    .A2(net2597),
    .B1(net3343),
    .B2(net3305),
    .X(_09094_));
 sky130_fd_sc_hd__nor2_1 _17141_ (.A(net6484),
    .B(net3325),
    .Y(_09095_));
 sky130_fd_sc_hd__buf_2 _17142_ (.A(_09095_),
    .X(_09096_));
 sky130_fd_sc_hd__buf_1 _17143_ (.A(net4047),
    .X(_09097_));
 sky130_fd_sc_hd__nor2_1 _17144_ (.A(_09097_),
    .B(net3305),
    .Y(_09098_));
 sky130_fd_sc_hd__a221o_1 _17145_ (.A1(net6483),
    .A2(_09094_),
    .B1(_09096_),
    .B2(net3341),
    .C1(_09098_),
    .X(_09099_));
 sky130_fd_sc_hd__nor2_1 _17146_ (.A(_09083_),
    .B(_09084_),
    .Y(_09100_));
 sky130_fd_sc_hd__or2_1 _17147_ (.A(net1504),
    .B(net822),
    .X(_09101_));
 sky130_fd_sc_hd__xnor2_2 _17148_ (.A(net1801),
    .B(_09101_),
    .Y(_09102_));
 sky130_fd_sc_hd__and2_1 _17149_ (.A(net6914),
    .B(_09086_),
    .X(_09103_));
 sky130_fd_sc_hd__a2111o_1 _17150_ (.A1(net6932),
    .A2(_09075_),
    .B1(_09076_),
    .C1(_09103_),
    .D1(_09064_),
    .X(_09104_));
 sky130_fd_sc_hd__or3_1 _17151_ (.A(net6932),
    .B(_09075_),
    .C(_09103_),
    .X(_09105_));
 sky130_fd_sc_hd__o211a_1 _17152_ (.A1(net6914),
    .A2(_09086_),
    .B1(_09104_),
    .C1(_09105_),
    .X(_09106_));
 sky130_fd_sc_hd__xor2_1 _17153_ (.A(_09102_),
    .B(net527),
    .X(_09107_));
 sky130_fd_sc_hd__o21a_1 _17154_ (.A1(net2199),
    .A2(_09107_),
    .B1(net8048),
    .X(_09108_));
 sky130_fd_sc_hd__nor2_1 _17155_ (.A(net3301),
    .B(_09108_),
    .Y(_09109_));
 sky130_fd_sc_hd__a31o_1 _17156_ (.A1(net3301),
    .A2(net1234),
    .A3(_09107_),
    .B1(_09109_),
    .X(_00335_));
 sky130_fd_sc_hd__nor2_1 _17157_ (.A(net4039),
    .B(_09097_),
    .Y(_09110_));
 sky130_fd_sc_hd__a31o_1 _17158_ (.A1(net4039),
    .A2(net4058),
    .A3(net3305),
    .B1(_09110_),
    .X(_09111_));
 sky130_fd_sc_hd__a22o_1 _17159_ (.A1(net2595),
    .A2(_09095_),
    .B1(_09111_),
    .B2(net6484),
    .X(_09112_));
 sky130_fd_sc_hd__or2_1 _17160_ (.A(_09098_),
    .B(_09112_),
    .X(_09113_));
 sky130_fd_sc_hd__inv_2 _17161_ (.A(net822),
    .Y(_09114_));
 sky130_fd_sc_hd__o21ai_1 _17162_ (.A1(net1801),
    .A2(_09114_),
    .B1(net1076),
    .Y(_09115_));
 sky130_fd_sc_hd__xnor2_1 _17163_ (.A(_09113_),
    .B(_09115_),
    .Y(_09116_));
 sky130_fd_sc_hd__a21o_1 _17164_ (.A1(_09102_),
    .A2(net527),
    .B1(net6901),
    .X(_09117_));
 sky130_fd_sc_hd__o21ai_1 _17165_ (.A1(_09102_),
    .A2(net527),
    .B1(_09117_),
    .Y(_09118_));
 sky130_fd_sc_hd__xnor2_1 _17166_ (.A(net670),
    .B(_09118_),
    .Y(_09119_));
 sky130_fd_sc_hd__a21oi_1 _17167_ (.A1(_09068_),
    .A2(_09119_),
    .B1(net6891),
    .Y(_09120_));
 sky130_fd_sc_hd__o211a_1 _17168_ (.A1(net1921),
    .A2(_09119_),
    .B1(net8048),
    .C1(net6891),
    .X(_09121_));
 sky130_fd_sc_hd__nor2_1 _17169_ (.A(_09120_),
    .B(_09121_),
    .Y(_00336_));
 sky130_fd_sc_hd__mux2_1 _17170_ (.A0(net5997),
    .A1(net3361),
    .S(_09096_),
    .X(_09122_));
 sky130_fd_sc_hd__or3_1 _17171_ (.A(net1801),
    .B(_09114_),
    .C(_09113_),
    .X(_09123_));
 sky130_fd_sc_hd__nand2_1 _17172_ (.A(net1076),
    .B(_09123_),
    .Y(_09124_));
 sky130_fd_sc_hd__xnor2_1 _17173_ (.A(_09122_),
    .B(_09124_),
    .Y(_09125_));
 sky130_fd_sc_hd__and2_1 _17174_ (.A(net6891),
    .B(net670),
    .X(_09126_));
 sky130_fd_sc_hd__a211o_1 _17175_ (.A1(net6901),
    .A2(_09102_),
    .B1(net527),
    .C1(_09126_),
    .X(_09127_));
 sky130_fd_sc_hd__or3_1 _17176_ (.A(net6901),
    .B(_09102_),
    .C(_09126_),
    .X(_09128_));
 sky130_fd_sc_hd__o211a_1 _17177_ (.A1(net6891),
    .A2(net670),
    .B1(_09127_),
    .C1(_09128_),
    .X(_09129_));
 sky130_fd_sc_hd__xnor2_1 _17178_ (.A(net618),
    .B(_09129_),
    .Y(_09130_));
 sky130_fd_sc_hd__a21o_1 _17179_ (.A1(net1475),
    .A2(_09130_),
    .B1(net3323),
    .X(_09131_));
 sky130_fd_sc_hd__or3_1 _17180_ (.A(net6850),
    .B(net1820),
    .C(_09130_),
    .X(_09132_));
 sky130_fd_sc_hd__a21bo_1 _17181_ (.A1(net6850),
    .A2(_09131_),
    .B1_N(_09132_),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _17182_ (.A0(net5997),
    .A1(net3344),
    .S(_09096_),
    .X(_09133_));
 sky130_fd_sc_hd__o21ai_1 _17183_ (.A1(_09122_),
    .A2(_09123_),
    .B1(net1076),
    .Y(_09134_));
 sky130_fd_sc_hd__xor2_1 _17184_ (.A(_09133_),
    .B(_09134_),
    .X(_09135_));
 sky130_fd_sc_hd__a21o_1 _17185_ (.A1(net618),
    .A2(_09129_),
    .B1(net6850),
    .X(_09136_));
 sky130_fd_sc_hd__o21ai_1 _17186_ (.A1(net618),
    .A2(_09129_),
    .B1(_09136_),
    .Y(_09137_));
 sky130_fd_sc_hd__xnor2_1 _17187_ (.A(net617),
    .B(_09137_),
    .Y(_09138_));
 sky130_fd_sc_hd__nor2_1 _17188_ (.A(net1922),
    .B(_09138_),
    .Y(_09139_));
 sky130_fd_sc_hd__a21o_1 _17189_ (.A1(net2932),
    .A2(_09138_),
    .B1(net4245),
    .X(_09140_));
 sky130_fd_sc_hd__mux2_1 _17190_ (.A0(_09139_),
    .A1(_09140_),
    .S(net6839),
    .X(_09141_));
 sky130_fd_sc_hd__clkbuf_1 _17191_ (.A(_09141_),
    .X(_00338_));
 sky130_fd_sc_hd__o31a_1 _17192_ (.A1(_09122_),
    .A2(_09123_),
    .A3(_09133_),
    .B1(net1076),
    .X(_09142_));
 sky130_fd_sc_hd__nand2_1 _17193_ (.A(net2592),
    .B(net3305),
    .Y(_09143_));
 sky130_fd_sc_hd__or2_1 _17194_ (.A(net2597),
    .B(_09143_),
    .X(_09144_));
 sky130_fd_sc_hd__a22o_1 _17195_ (.A1(net3343),
    .A2(_09096_),
    .B1(_09144_),
    .B2(net5988),
    .X(_09145_));
 sky130_fd_sc_hd__xor2_2 _17196_ (.A(_09142_),
    .B(_09145_),
    .X(_09146_));
 sky130_fd_sc_hd__inv_2 _17197_ (.A(net617),
    .Y(_09147_));
 sky130_fd_sc_hd__a221o_1 _17198_ (.A1(net6850),
    .A2(net618),
    .B1(_09147_),
    .B2(net6841),
    .C1(_09129_),
    .X(_09148_));
 sky130_fd_sc_hd__nor2_1 _17199_ (.A(net6850),
    .B(net618),
    .Y(_09149_));
 sky130_fd_sc_hd__a21bo_1 _17200_ (.A1(net617),
    .A2(_09149_),
    .B1_N(net6841),
    .X(_09150_));
 sky130_fd_sc_hd__o21ai_1 _17201_ (.A1(net617),
    .A2(_09149_),
    .B1(_09150_),
    .Y(_09151_));
 sky130_fd_sc_hd__nand2_1 _17202_ (.A(_09148_),
    .B(_09151_),
    .Y(_09152_));
 sky130_fd_sc_hd__xor2_1 _17203_ (.A(_09146_),
    .B(_09152_),
    .X(_09153_));
 sky130_fd_sc_hd__a21o_1 _17204_ (.A1(net1815),
    .A2(_09153_),
    .B1(net4245),
    .X(_09154_));
 sky130_fd_sc_hd__nor2_1 _17205_ (.A(net1922),
    .B(_09153_),
    .Y(_09155_));
 sky130_fd_sc_hd__inv_2 _17206_ (.A(net6810),
    .Y(_09156_));
 sky130_fd_sc_hd__clkbuf_1 _17207_ (.A(net4036),
    .X(_09157_));
 sky130_fd_sc_hd__clkbuf_1 _17208_ (.A(net3285),
    .X(_09158_));
 sky130_fd_sc_hd__mux2_1 _17209_ (.A0(_09154_),
    .A1(_09155_),
    .S(net2587),
    .X(_09159_));
 sky130_fd_sc_hd__clkbuf_1 _17210_ (.A(_09159_),
    .X(_00339_));
 sky130_fd_sc_hd__a31o_1 _17211_ (.A1(_09146_),
    .A2(_09148_),
    .A3(_09151_),
    .B1(net6819),
    .X(_09160_));
 sky130_fd_sc_hd__a21o_1 _17212_ (.A1(_09148_),
    .A2(_09151_),
    .B1(_09146_),
    .X(_09161_));
 sky130_fd_sc_hd__and2_1 _17213_ (.A(_09160_),
    .B(_09161_),
    .X(_09162_));
 sky130_fd_sc_hd__a21oi_2 _17214_ (.A1(net966),
    .A2(_09145_),
    .B1(_09142_),
    .Y(_09163_));
 sky130_fd_sc_hd__nor2_1 _17215_ (.A(_08835_),
    .B(_09006_),
    .Y(_09164_));
 sky130_fd_sc_hd__mux2_2 _17216_ (.A0(net5998),
    .A1(_08834_),
    .S(net2583),
    .X(_09165_));
 sky130_fd_sc_hd__xnor2_1 _17217_ (.A(_09163_),
    .B(_09165_),
    .Y(_09166_));
 sky130_fd_sc_hd__xnor2_1 _17218_ (.A(_09162_),
    .B(_09166_),
    .Y(_09167_));
 sky130_fd_sc_hd__a21o_1 _17219_ (.A1(net2187),
    .A2(_09167_),
    .B1(net3324),
    .X(_09168_));
 sky130_fd_sc_hd__or3_1 _17220_ (.A(net6788),
    .B(net1821),
    .C(_09167_),
    .X(_09169_));
 sky130_fd_sc_hd__a21bo_1 _17221_ (.A1(net6788),
    .A2(_09168_),
    .B1_N(_09169_),
    .X(_00340_));
 sky130_fd_sc_hd__buf_1 _17222_ (.A(net3290),
    .X(_09170_));
 sky130_fd_sc_hd__nor2_1 _17223_ (.A(net6806),
    .B(_09165_),
    .Y(_09171_));
 sky130_fd_sc_hd__inv_2 _17224_ (.A(_09165_),
    .Y(_09172_));
 sky130_fd_sc_hd__nand2_1 _17225_ (.A(net6806),
    .B(_09163_),
    .Y(_09173_));
 sky130_fd_sc_hd__o211a_1 _17226_ (.A1(net6791),
    .A2(_09172_),
    .B1(_09173_),
    .C1(_09162_),
    .X(_09174_));
 sky130_fd_sc_hd__and4_1 _17227_ (.A(net6791),
    .B(net966),
    .C(_09163_),
    .D(_09165_),
    .X(_09175_));
 sky130_fd_sc_hd__inv_2 _17228_ (.A(net6799),
    .Y(_09176_));
 sky130_fd_sc_hd__buf_1 _17229_ (.A(_09176_),
    .X(_09177_));
 sky130_fd_sc_hd__or2_1 _17230_ (.A(net3280),
    .B(_09165_),
    .X(_09178_));
 sky130_fd_sc_hd__nand2_1 _17231_ (.A(net3280),
    .B(net1502),
    .Y(_09179_));
 sky130_fd_sc_hd__a21oi_1 _17232_ (.A1(_09178_),
    .A2(_09179_),
    .B1(_09162_),
    .Y(_09180_));
 sky130_fd_sc_hd__a2111o_1 _17233_ (.A1(_09163_),
    .A2(_09171_),
    .B1(_09174_),
    .C1(_09175_),
    .D1(_09180_),
    .X(_09181_));
 sky130_fd_sc_hd__xnor2_1 _17234_ (.A(_09170_),
    .B(_09181_),
    .Y(_09182_));
 sky130_fd_sc_hd__a21o_1 _17235_ (.A1(net2186),
    .A2(_09182_),
    .B1(_09023_),
    .X(_09183_));
 sky130_fd_sc_hd__or3_1 _17236_ (.A(net6759),
    .B(_08911_),
    .C(_09182_),
    .X(_09184_));
 sky130_fd_sc_hd__a21bo_1 _17237_ (.A1(net6759),
    .A2(_09183_),
    .B1_N(_09184_),
    .X(_00341_));
 sky130_fd_sc_hd__buf_1 _17238_ (.A(net2957),
    .X(_09185_));
 sky130_fd_sc_hd__inv_2 _17239_ (.A(\svm0.state[1] ),
    .Y(_09186_));
 sky130_fd_sc_hd__inv_2 _17240_ (.A(\svm0.state[0] ),
    .Y(_09187_));
 sky130_fd_sc_hd__mux2_1 _17241_ (.A0(net3387),
    .A1(_09186_),
    .S(_09187_),
    .X(_09188_));
 sky130_fd_sc_hd__buf_1 _17242_ (.A(_09188_),
    .X(_09189_));
 sky130_fd_sc_hd__buf_1 _17243_ (.A(net2161),
    .X(_09190_));
 sky130_fd_sc_hd__a22o_1 _17244_ (.A1(net2165),
    .A2(net325),
    .B1(net1800),
    .B2(net9155),
    .X(_00342_));
 sky130_fd_sc_hd__a22o_1 _17245_ (.A1(net2165),
    .A2(net288),
    .B1(net1800),
    .B2(net9054),
    .X(_00343_));
 sky130_fd_sc_hd__a22o_1 _17246_ (.A1(net2165),
    .A2(net285),
    .B1(net1800),
    .B2(net9204),
    .X(_00344_));
 sky130_fd_sc_hd__a22o_1 _17247_ (.A1(net2165),
    .A2(net224),
    .B1(net1800),
    .B2(net9167),
    .X(_00345_));
 sky130_fd_sc_hd__a22o_1 _17248_ (.A1(net2164),
    .A2(net257),
    .B1(net1799),
    .B2(net9140),
    .X(_00346_));
 sky130_fd_sc_hd__a22o_1 _17249_ (.A1(net2164),
    .A2(net192),
    .B1(net1799),
    .B2(net9132),
    .X(_00347_));
 sky130_fd_sc_hd__a22o_1 _17250_ (.A1(net2164),
    .A2(net221),
    .B1(net1799),
    .B2(net9090),
    .X(_00348_));
 sky130_fd_sc_hd__a22o_1 _17251_ (.A1(net2164),
    .A2(net190),
    .B1(net1799),
    .B2(net9219),
    .X(_00349_));
 sky130_fd_sc_hd__a22o_1 _17252_ (.A1(_09185_),
    .A2(net218),
    .B1(_09190_),
    .B2(net9099),
    .X(_00350_));
 sky130_fd_sc_hd__a22o_1 _17253_ (.A1(_09185_),
    .A2(net187),
    .B1(_09190_),
    .B2(net9080),
    .X(_00351_));
 sky130_fd_sc_hd__a22o_1 _17254_ (.A1(net2958),
    .A2(net174),
    .B1(net2163),
    .B2(net9165),
    .X(_00352_));
 sky130_fd_sc_hd__a22o_1 _17255_ (.A1(net2958),
    .A2(net157),
    .B1(net2161),
    .B2(net9176),
    .X(_00353_));
 sky130_fd_sc_hd__a22o_1 _17256_ (.A1(net2959),
    .A2(net158),
    .B1(net2162),
    .B2(net9141),
    .X(_00354_));
 sky130_fd_sc_hd__a22o_1 _17257_ (.A1(net2959),
    .A2(net155),
    .B1(net2162),
    .B2(net9129),
    .X(_00355_));
 sky130_fd_sc_hd__a22o_1 _17258_ (.A1(net2960),
    .A2(net154),
    .B1(_09189_),
    .B2(net9096),
    .X(_00356_));
 sky130_fd_sc_hd__a32o_1 _17259_ (.A1(net7606),
    .A2(net2960),
    .A3(net153),
    .B1(net2163),
    .B2(net9214),
    .X(_00357_));
 sky130_fd_sc_hd__buf_1 _17260_ (.A(net2981),
    .X(_09191_));
 sky130_fd_sc_hd__mux2_1 _17261_ (.A0(net3387),
    .A1(_09187_),
    .S(_09186_),
    .X(_09192_));
 sky130_fd_sc_hd__clkbuf_1 _17262_ (.A(_09192_),
    .X(_09193_));
 sky130_fd_sc_hd__clkbuf_1 _17263_ (.A(net2156),
    .X(_09194_));
 sky130_fd_sc_hd__a22o_1 _17264_ (.A1(net2160),
    .A2(net323),
    .B1(net1798),
    .B2(net9089),
    .X(_00358_));
 sky130_fd_sc_hd__a22o_1 _17265_ (.A1(net2160),
    .A2(net287),
    .B1(net1798),
    .B2(net9108),
    .X(_00359_));
 sky130_fd_sc_hd__a22o_1 _17266_ (.A1(net2160),
    .A2(net284),
    .B1(net1798),
    .B2(\svm0.tA[2] ),
    .X(_00360_));
 sky130_fd_sc_hd__a22o_1 _17267_ (.A1(net2160),
    .A2(net223),
    .B1(net1797),
    .B2(\svm0.tA[3] ),
    .X(_00361_));
 sky130_fd_sc_hd__a22o_1 _17268_ (.A1(net2160),
    .A2(net256),
    .B1(net1797),
    .B2(net9186),
    .X(_00362_));
 sky130_fd_sc_hd__a22o_1 _17269_ (.A1(net2159),
    .A2(net191),
    .B1(net1797),
    .B2(net9136),
    .X(_00363_));
 sky130_fd_sc_hd__a22o_1 _17270_ (.A1(net2159),
    .A2(net220),
    .B1(net1797),
    .B2(net9093),
    .X(_00364_));
 sky130_fd_sc_hd__a22o_1 _17271_ (.A1(net2159),
    .A2(net189),
    .B1(net1797),
    .B2(net9220),
    .X(_00365_));
 sky130_fd_sc_hd__a22o_1 _17272_ (.A1(_09191_),
    .A2(net218),
    .B1(net1798),
    .B2(net9100),
    .X(_00366_));
 sky130_fd_sc_hd__a22o_1 _17273_ (.A1(_09191_),
    .A2(net187),
    .B1(net1798),
    .B2(net8971),
    .X(_00367_));
 sky130_fd_sc_hd__a22o_1 _17274_ (.A1(net2982),
    .A2(net174),
    .B1(net2157),
    .B2(net9172),
    .X(_00368_));
 sky130_fd_sc_hd__a22o_1 _17275_ (.A1(net2982),
    .A2(net157),
    .B1(net2157),
    .B2(net9232),
    .X(_00369_));
 sky130_fd_sc_hd__a22o_1 _17276_ (.A1(net2981),
    .A2(net158),
    .B1(net2156),
    .B2(net9143),
    .X(_00370_));
 sky130_fd_sc_hd__a22o_1 _17277_ (.A1(net2983),
    .A2(net155),
    .B1(net2158),
    .B2(net9131),
    .X(_00371_));
 sky130_fd_sc_hd__a22o_1 _17278_ (.A1(net2984),
    .A2(net154),
    .B1(_09193_),
    .B2(net9111),
    .X(_00372_));
 sky130_fd_sc_hd__a32o_1 _17279_ (.A1(net7606),
    .A2(net2983),
    .A3(net153),
    .B1(net2158),
    .B2(net9190),
    .X(_00373_));
 sky130_fd_sc_hd__nor2_1 _17280_ (.A(_08646_),
    .B(net4067),
    .Y(_09195_));
 sky130_fd_sc_hd__inv_2 _17281_ (.A(net6741),
    .Y(_09196_));
 sky130_fd_sc_hd__or4_1 _17282_ (.A(net4035),
    .B(net6738),
    .C(\svm0.counter[3] ),
    .D(net6736),
    .X(_09197_));
 sky130_fd_sc_hd__or4_1 _17283_ (.A(net6732),
    .B(net6716),
    .C(net6708),
    .D(net6745),
    .X(_09198_));
 sky130_fd_sc_hd__or4_1 _17284_ (.A(\svm0.counter[8] ),
    .B(\svm0.counter[11] ),
    .C(\svm0.counter[10] ),
    .D(net6693),
    .X(_09199_));
 sky130_fd_sc_hd__or2_1 _17285_ (.A(_09198_),
    .B(_09199_),
    .X(_09200_));
 sky130_fd_sc_hd__or4_1 _17286_ (.A(net6727),
    .B(net6719),
    .C(_09197_),
    .D(_09200_),
    .X(_09201_));
 sky130_fd_sc_hd__or4_1 _17287_ (.A(net6700),
    .B(net6684),
    .C(net6688),
    .D(_09201_),
    .X(_09202_));
 sky130_fd_sc_hd__nand2_1 _17288_ (.A(_09195_),
    .B(_09202_),
    .Y(_09203_));
 sky130_fd_sc_hd__nand2_1 _17289_ (.A(net6669),
    .B(net1796),
    .Y(_09204_));
 sky130_fd_sc_hd__o21a_1 _17290_ (.A1(net9199),
    .A2(net1924),
    .B1(net1462),
    .X(_00374_));
 sky130_fd_sc_hd__inv_2 _17291_ (.A(net6687),
    .Y(_09205_));
 sky130_fd_sc_hd__or2_1 _17292_ (.A(net7943),
    .B(net7919),
    .X(_09206_));
 sky130_fd_sc_hd__or3_1 _17293_ (.A(net7890),
    .B(net7862),
    .C(_09206_),
    .X(_09207_));
 sky130_fd_sc_hd__or2_1 _17294_ (.A(net7828),
    .B(_09207_),
    .X(_09208_));
 sky130_fd_sc_hd__or2_1 _17295_ (.A(net7806),
    .B(_09208_),
    .X(_09209_));
 sky130_fd_sc_hd__or2_1 _17296_ (.A(net7787),
    .B(_09209_),
    .X(_09210_));
 sky130_fd_sc_hd__or4_1 _17297_ (.A(net7765),
    .B(net7742),
    .C(net7719),
    .D(net1795),
    .X(_09211_));
 sky130_fd_sc_hd__or2_1 _17298_ (.A(net7702),
    .B(_09211_),
    .X(_09212_));
 sky130_fd_sc_hd__or2_1 _17299_ (.A(net7682),
    .B(_09212_),
    .X(_09213_));
 sky130_fd_sc_hd__or3_2 _17300_ (.A(net7661),
    .B(net7643),
    .C(_09213_),
    .X(_09214_));
 sky130_fd_sc_hd__inv_2 _17301_ (.A(net6685),
    .Y(_09215_));
 sky130_fd_sc_hd__o311a_1 _17302_ (.A1(_09205_),
    .A2(net7630),
    .A3(_09214_),
    .B1(net7607),
    .C1(net4031),
    .X(_09216_));
 sky130_fd_sc_hd__nand2_1 _17303_ (.A(_09205_),
    .B(net7630),
    .Y(_09217_));
 sky130_fd_sc_hd__o211ai_1 _17304_ (.A1(net7661),
    .A2(_09213_),
    .B1(_09217_),
    .C1(net7643),
    .Y(_09218_));
 sky130_fd_sc_hd__o21ai_1 _17305_ (.A1(net7661),
    .A2(_09213_),
    .B1(net7643),
    .Y(_09219_));
 sky130_fd_sc_hd__a31oi_1 _17306_ (.A1(_09214_),
    .A2(_09217_),
    .A3(_09219_),
    .B1(net6691),
    .Y(_09220_));
 sky130_fd_sc_hd__nor3_1 _17307_ (.A(net7765),
    .B(net7742),
    .C(net1795),
    .Y(_09221_));
 sky130_fd_sc_hd__o21a_1 _17308_ (.A1(net7765),
    .A2(net1795),
    .B1(net7742),
    .X(_09222_));
 sky130_fd_sc_hd__inv_2 _17309_ (.A(\svm0.counter[8] ),
    .Y(_09223_));
 sky130_fd_sc_hd__xnor2_1 _17310_ (.A(net6709),
    .B(net7719),
    .Y(_09224_));
 sky130_fd_sc_hd__nand2_1 _17311_ (.A(net4024),
    .B(_09224_),
    .Y(_09225_));
 sky130_fd_sc_hd__mux2_1 _17312_ (.A0(_09221_),
    .A1(_09222_),
    .S(_09224_),
    .X(_09226_));
 sky130_fd_sc_hd__nand2_1 _17313_ (.A(net6711),
    .B(_09226_),
    .Y(_09227_));
 sky130_fd_sc_hd__o31a_1 _17314_ (.A1(_09221_),
    .A2(_09222_),
    .A3(_09225_),
    .B1(_09227_),
    .X(_09228_));
 sky130_fd_sc_hd__xor2_1 _17315_ (.A(net6714),
    .B(net7764),
    .X(_09229_));
 sky130_fd_sc_hd__inv_2 _17316_ (.A(net6728),
    .Y(_09230_));
 sky130_fd_sc_hd__nand2_1 _17317_ (.A(net7806),
    .B(_09208_),
    .Y(_09231_));
 sky130_fd_sc_hd__xnor2_1 _17318_ (.A(net6720),
    .B(net7787),
    .Y(_09232_));
 sky130_fd_sc_hd__mux2_1 _17319_ (.A0(_09209_),
    .A1(_09231_),
    .S(_09232_),
    .X(_09233_));
 sky130_fd_sc_hd__nor2_1 _17320_ (.A(net4022),
    .B(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__and4_1 _17321_ (.A(net4022),
    .B(_09209_),
    .C(_09231_),
    .D(_09232_),
    .X(_09235_));
 sky130_fd_sc_hd__xor2_1 _17322_ (.A(net6737),
    .B(net7919),
    .X(_09236_));
 sky130_fd_sc_hd__nor2_1 _17323_ (.A(net4032),
    .B(net7943),
    .Y(_09237_));
 sky130_fd_sc_hd__nor2_1 _17324_ (.A(_04973_),
    .B(_09236_),
    .Y(_09238_));
 sky130_fd_sc_hd__a22o_1 _17325_ (.A1(_09236_),
    .A2(_09237_),
    .B1(_09238_),
    .B2(net4032),
    .X(_09239_));
 sky130_fd_sc_hd__xnor2_1 _17326_ (.A(net6733),
    .B(net7890),
    .Y(_09240_));
 sky130_fd_sc_hd__xnor2_1 _17327_ (.A(_09206_),
    .B(_09240_),
    .Y(_09241_));
 sky130_fd_sc_hd__o211ai_1 _17328_ (.A1(net4028),
    .A2(net7608),
    .B1(_09239_),
    .C1(_09241_),
    .Y(_09242_));
 sky130_fd_sc_hd__inv_2 _17329_ (.A(\svm0.counter[3] ),
    .Y(_09243_));
 sky130_fd_sc_hd__o21ai_1 _17330_ (.A1(net7890),
    .A2(_09206_),
    .B1(net7862),
    .Y(_09244_));
 sky130_fd_sc_hd__xnor2_1 _17331_ (.A(net6730),
    .B(net7828),
    .Y(_09245_));
 sky130_fd_sc_hd__mux2_1 _17332_ (.A0(_09207_),
    .A1(_09244_),
    .S(_09245_),
    .X(_09246_));
 sky130_fd_sc_hd__and4_1 _17333_ (.A(net4017),
    .B(_09207_),
    .C(_09244_),
    .D(_09245_),
    .X(_09247_));
 sky130_fd_sc_hd__o21ba_1 _17334_ (.A1(net4017),
    .A2(_09246_),
    .B1_N(_09247_),
    .X(_09248_));
 sky130_fd_sc_hd__a211oi_1 _17335_ (.A1(_09210_),
    .A2(_09229_),
    .B1(_09242_),
    .C1(_09248_),
    .Y(_09249_));
 sky130_fd_sc_hd__o221ai_2 _17336_ (.A1(_09210_),
    .A2(_09229_),
    .B1(_09234_),
    .B2(_09235_),
    .C1(_09249_),
    .Y(_09250_));
 sky130_fd_sc_hd__or2_1 _17337_ (.A(net6698),
    .B(net7661),
    .X(_09251_));
 sky130_fd_sc_hd__nand2_1 _17338_ (.A(net6698),
    .B(net7661),
    .Y(_09252_));
 sky130_fd_sc_hd__and3_1 _17339_ (.A(_09213_),
    .B(_09251_),
    .C(_09252_),
    .X(_09253_));
 sky130_fd_sc_hd__a21oi_1 _17340_ (.A1(_09251_),
    .A2(_09252_),
    .B1(_09213_),
    .Y(_09254_));
 sky130_fd_sc_hd__or4_1 _17341_ (.A(_09228_),
    .B(net1220),
    .C(_09253_),
    .D(_09254_),
    .X(_09255_));
 sky130_fd_sc_hd__a311o_1 _17342_ (.A1(net6691),
    .A2(_09214_),
    .A3(_09218_),
    .B1(_09220_),
    .C1(_09255_),
    .X(_09256_));
 sky130_fd_sc_hd__inv_2 _17343_ (.A(\svm0.counter[10] ),
    .Y(_09257_));
 sky130_fd_sc_hd__buf_1 _17344_ (.A(net4016),
    .X(_09258_));
 sky130_fd_sc_hd__nand2_1 _17345_ (.A(net7702),
    .B(_09211_),
    .Y(_09259_));
 sky130_fd_sc_hd__xnor2_1 _17346_ (.A(net6703),
    .B(net7682),
    .Y(_09260_));
 sky130_fd_sc_hd__mux2_1 _17347_ (.A0(_09212_),
    .A1(_09259_),
    .S(_09260_),
    .X(_09261_));
 sky130_fd_sc_hd__and4_1 _17348_ (.A(net3278),
    .B(_09212_),
    .C(_09259_),
    .D(_09260_),
    .X(_09262_));
 sky130_fd_sc_hd__o21bai_1 _17349_ (.A1(net3278),
    .A2(_09261_),
    .B1_N(_09262_),
    .Y(_09263_));
 sky130_fd_sc_hd__o21a_1 _17350_ (.A1(net7630),
    .A2(_09214_),
    .B1(_09205_),
    .X(_09264_));
 sky130_fd_sc_hd__a221o_1 _17351_ (.A1(net4031),
    .A2(net7607),
    .B1(_09214_),
    .B2(net7630),
    .C1(_09264_),
    .X(_09265_));
 sky130_fd_sc_hd__and4bb_1 _17352_ (.A_N(_09216_),
    .B_N(_09256_),
    .C(_09263_),
    .D(_09265_),
    .X(_09266_));
 sky130_fd_sc_hd__a21bo_1 _17353_ (.A1(net6658),
    .A2(net771),
    .B1_N(\svm0.rising ),
    .X(_09267_));
 sky130_fd_sc_hd__nand2_1 _17354_ (.A(net1465),
    .B(_09267_),
    .Y(_00375_));
 sky130_fd_sc_hd__nand2_1 _17355_ (.A(net6658),
    .B(net4253),
    .Y(_09268_));
 sky130_fd_sc_hd__a21oi_1 _17356_ (.A1(\svm0.rising ),
    .A2(net771),
    .B1(net1796),
    .Y(_09269_));
 sky130_fd_sc_hd__nor2_1 _17357_ (.A(net3276),
    .B(_09269_),
    .Y(_09270_));
 sky130_fd_sc_hd__and2_1 _17358_ (.A(net7377),
    .B(net669),
    .X(_09271_));
 sky130_fd_sc_hd__buf_1 _17359_ (.A(net3277),
    .X(_09272_));
 sky130_fd_sc_hd__o21ba_1 _17360_ (.A1(net6657),
    .A2(net3389),
    .B1_N(_09269_),
    .X(_09273_));
 sky130_fd_sc_hd__o21ai_1 _17361_ (.A1(net7377),
    .A2(net2579),
    .B1(net667),
    .Y(_09274_));
 sky130_fd_sc_hd__mux2_1 _17362_ (.A0(_09271_),
    .A1(_09274_),
    .S(\svm0.delta[1] ),
    .X(_09275_));
 sky130_fd_sc_hd__clkbuf_1 _17363_ (.A(_09275_),
    .X(_00376_));
 sky130_fd_sc_hd__buf_1 _17364_ (.A(net669),
    .X(_09276_));
 sky130_fd_sc_hd__o21a_1 _17365_ (.A1(net7377),
    .A2(\svm0.delta[1] ),
    .B1(_09276_),
    .X(_09277_));
 sky130_fd_sc_hd__buf_1 _17366_ (.A(net3276),
    .X(_09278_));
 sky130_fd_sc_hd__o31ai_1 _17367_ (.A1(net7377),
    .A2(\svm0.delta[1] ),
    .A3(net2573),
    .B1(net667),
    .Y(_09279_));
 sky130_fd_sc_hd__mux2_1 _17368_ (.A0(_09277_),
    .A1(_09279_),
    .S(\svm0.delta[2] ),
    .X(_09280_));
 sky130_fd_sc_hd__clkbuf_1 _17369_ (.A(_09280_),
    .X(_00377_));
 sky130_fd_sc_hd__inv_2 _17370_ (.A(\svm0.delta[3] ),
    .Y(_09281_));
 sky130_fd_sc_hd__buf_1 _17371_ (.A(net667),
    .X(_09282_));
 sky130_fd_sc_hd__and2_1 _17372_ (.A(_09281_),
    .B(net667),
    .X(_09283_));
 sky130_fd_sc_hd__or3_1 _17373_ (.A(net7377),
    .B(\svm0.delta[1] ),
    .C(net6743),
    .X(_09284_));
 sky130_fd_sc_hd__mux2_1 _17374_ (.A0(\svm0.delta[3] ),
    .A1(_09283_),
    .S(_09284_),
    .X(_09285_));
 sky130_fd_sc_hd__clkbuf_1 _17375_ (.A(_09195_),
    .X(_09286_));
 sky130_fd_sc_hd__a2bb2o_1 _17376_ (.A1_N(_09281_),
    .A2_N(_09282_),
    .B1(_09285_),
    .B2(net2567),
    .X(_00378_));
 sky130_fd_sc_hd__inv_2 _17377_ (.A(\svm0.delta[4] ),
    .Y(_09287_));
 sky130_fd_sc_hd__or2_1 _17378_ (.A(\svm0.delta[3] ),
    .B(_09284_),
    .X(_09288_));
 sky130_fd_sc_hd__or2_1 _17379_ (.A(net2572),
    .B(_09288_),
    .X(_09289_));
 sky130_fd_sc_hd__a21oi_1 _17380_ (.A1(net612),
    .A2(_09289_),
    .B1(_09287_),
    .Y(_09290_));
 sky130_fd_sc_hd__a31o_1 _17381_ (.A1(_09287_),
    .A2(net614),
    .A3(_09288_),
    .B1(_09290_),
    .X(_00379_));
 sky130_fd_sc_hd__inv_2 _17382_ (.A(\svm0.delta[5] ),
    .Y(_09291_));
 sky130_fd_sc_hd__or2_1 _17383_ (.A(\svm0.delta[4] ),
    .B(_09288_),
    .X(_09292_));
 sky130_fd_sc_hd__or2_1 _17384_ (.A(net2572),
    .B(_09292_),
    .X(_09293_));
 sky130_fd_sc_hd__a21oi_1 _17385_ (.A1(net612),
    .A2(_09293_),
    .B1(_09291_),
    .Y(_09294_));
 sky130_fd_sc_hd__a31o_1 _17386_ (.A1(_09291_),
    .A2(net614),
    .A3(_09292_),
    .B1(_09294_),
    .X(_00380_));
 sky130_fd_sc_hd__inv_2 _17387_ (.A(\svm0.delta[6] ),
    .Y(_09295_));
 sky130_fd_sc_hd__or2_1 _17388_ (.A(\svm0.delta[5] ),
    .B(_09292_),
    .X(_09296_));
 sky130_fd_sc_hd__or2_1 _17389_ (.A(net2572),
    .B(_09296_),
    .X(_09297_));
 sky130_fd_sc_hd__a21oi_1 _17390_ (.A1(net612),
    .A2(_09297_),
    .B1(_09295_),
    .Y(_09298_));
 sky130_fd_sc_hd__a31o_1 _17391_ (.A1(_09295_),
    .A2(net614),
    .A3(_09296_),
    .B1(_09298_),
    .X(_00381_));
 sky130_fd_sc_hd__inv_2 _17392_ (.A(\svm0.delta[7] ),
    .Y(_09299_));
 sky130_fd_sc_hd__or2_1 _17393_ (.A(\svm0.delta[6] ),
    .B(_09296_),
    .X(_09300_));
 sky130_fd_sc_hd__or2_1 _17394_ (.A(net2572),
    .B(_09300_),
    .X(_09301_));
 sky130_fd_sc_hd__a21oi_1 _17395_ (.A1(net612),
    .A2(_09301_),
    .B1(_09299_),
    .Y(_09302_));
 sky130_fd_sc_hd__a31o_1 _17396_ (.A1(_09299_),
    .A2(net614),
    .A3(_09300_),
    .B1(_09302_),
    .X(_00382_));
 sky130_fd_sc_hd__inv_2 _17397_ (.A(\svm0.delta[8] ),
    .Y(_09303_));
 sky130_fd_sc_hd__or2_1 _17398_ (.A(\svm0.delta[7] ),
    .B(_09300_),
    .X(_09304_));
 sky130_fd_sc_hd__or2_1 _17399_ (.A(net2573),
    .B(net1461),
    .X(_09305_));
 sky130_fd_sc_hd__a21oi_1 _17400_ (.A1(net613),
    .A2(_09305_),
    .B1(_09303_),
    .Y(_09306_));
 sky130_fd_sc_hd__a31o_1 _17401_ (.A1(_09303_),
    .A2(net616),
    .A3(net1461),
    .B1(_09306_),
    .X(_00383_));
 sky130_fd_sc_hd__inv_2 _17402_ (.A(\svm0.delta[9] ),
    .Y(_09307_));
 sky130_fd_sc_hd__or2_1 _17403_ (.A(\svm0.delta[8] ),
    .B(net1461),
    .X(_09308_));
 sky130_fd_sc_hd__or2_1 _17404_ (.A(net2574),
    .B(_09308_),
    .X(_09309_));
 sky130_fd_sc_hd__a21oi_1 _17405_ (.A1(net613),
    .A2(_09309_),
    .B1(_09307_),
    .Y(_09310_));
 sky130_fd_sc_hd__a31o_1 _17406_ (.A1(_09307_),
    .A2(net616),
    .A3(_09308_),
    .B1(_09310_),
    .X(_00384_));
 sky130_fd_sc_hd__inv_2 _17407_ (.A(\svm0.delta[10] ),
    .Y(_09311_));
 sky130_fd_sc_hd__or2_1 _17408_ (.A(\svm0.delta[9] ),
    .B(_09308_),
    .X(_09312_));
 sky130_fd_sc_hd__or2_1 _17409_ (.A(net2575),
    .B(_09312_),
    .X(_09313_));
 sky130_fd_sc_hd__a21oi_1 _17410_ (.A1(net611),
    .A2(_09313_),
    .B1(_09311_),
    .Y(_09314_));
 sky130_fd_sc_hd__a31o_1 _17411_ (.A1(_09311_),
    .A2(net615),
    .A3(_09312_),
    .B1(_09314_),
    .X(_00385_));
 sky130_fd_sc_hd__inv_2 _17412_ (.A(\svm0.delta[11] ),
    .Y(_09315_));
 sky130_fd_sc_hd__or2_1 _17413_ (.A(\svm0.delta[10] ),
    .B(_09312_),
    .X(_09316_));
 sky130_fd_sc_hd__or2_1 _17414_ (.A(net3276),
    .B(_09316_),
    .X(_09317_));
 sky130_fd_sc_hd__a21oi_1 _17415_ (.A1(net611),
    .A2(_09317_),
    .B1(_09315_),
    .Y(_09318_));
 sky130_fd_sc_hd__a31o_1 _17416_ (.A1(_09315_),
    .A2(net615),
    .A3(_09316_),
    .B1(_09318_),
    .X(_00386_));
 sky130_fd_sc_hd__inv_2 _17417_ (.A(\svm0.delta[12] ),
    .Y(_09319_));
 sky130_fd_sc_hd__or2_1 _17418_ (.A(\svm0.delta[11] ),
    .B(_09316_),
    .X(_09320_));
 sky130_fd_sc_hd__or2_1 _17419_ (.A(net3276),
    .B(_09320_),
    .X(_09321_));
 sky130_fd_sc_hd__a21oi_1 _17420_ (.A1(net611),
    .A2(_09321_),
    .B1(_09319_),
    .Y(_09322_));
 sky130_fd_sc_hd__a31o_1 _17421_ (.A1(_09319_),
    .A2(net615),
    .A3(_09320_),
    .B1(_09322_),
    .X(_00387_));
 sky130_fd_sc_hd__o21a_1 _17422_ (.A1(\svm0.delta[12] ),
    .A2(_09320_),
    .B1(net668),
    .X(_09323_));
 sky130_fd_sc_hd__xnor2_1 _17423_ (.A(net9162),
    .B(_09323_),
    .Y(_09324_));
 sky130_fd_sc_hd__nor2_1 _17424_ (.A(net2615),
    .B(_09324_),
    .Y(_00388_));
 sky130_fd_sc_hd__or3_1 _17425_ (.A(\svm0.delta[12] ),
    .B(net6742),
    .C(_09320_),
    .X(_09325_));
 sky130_fd_sc_hd__and2_1 _17426_ (.A(_09270_),
    .B(_09325_),
    .X(_09326_));
 sky130_fd_sc_hd__o21ai_1 _17427_ (.A1(_09278_),
    .A2(_09325_),
    .B1(net668),
    .Y(_09327_));
 sky130_fd_sc_hd__mux2_1 _17428_ (.A0(_09326_),
    .A1(_09327_),
    .S(\svm0.delta[14] ),
    .X(_09328_));
 sky130_fd_sc_hd__clkbuf_1 _17429_ (.A(_09328_),
    .X(_00389_));
 sky130_fd_sc_hd__o21ai_1 _17430_ (.A1(\svm0.delta[14] ),
    .A2(_09325_),
    .B1(_09273_),
    .Y(_09329_));
 sky130_fd_sc_hd__nand2_1 _17431_ (.A(net9213),
    .B(_09329_),
    .Y(_09330_));
 sky130_fd_sc_hd__or2_1 _17432_ (.A(\svm0.delta[15] ),
    .B(_09329_),
    .X(_09331_));
 sky130_fd_sc_hd__a21oi_1 _17433_ (.A1(_09330_),
    .A2(_09331_),
    .B1(_08648_),
    .Y(_00390_));
 sky130_fd_sc_hd__buf_1 _17434_ (.A(net4067),
    .X(_09332_));
 sky130_fd_sc_hd__o21a_1 _17435_ (.A1(net7376),
    .A2(net3274),
    .B1(net6656),
    .X(_09333_));
 sky130_fd_sc_hd__nor2_1 _17436_ (.A(net4035),
    .B(_09333_),
    .Y(_09334_));
 sky130_fd_sc_hd__a31o_1 _17437_ (.A1(net4035),
    .A2(net7376),
    .A3(net2570),
    .B1(_09334_),
    .X(_00391_));
 sky130_fd_sc_hd__nand2_1 _17438_ (.A(net6741),
    .B(net7376),
    .Y(_09335_));
 sky130_fd_sc_hd__xor2_1 _17439_ (.A(net6744),
    .B(_09335_),
    .X(_09336_));
 sky130_fd_sc_hd__a21o_1 _17440_ (.A1(net4251),
    .A2(_09336_),
    .B1(net3386),
    .X(_09337_));
 sky130_fd_sc_hd__nor2_1 _17441_ (.A(net2578),
    .B(_09336_),
    .Y(_09338_));
 sky130_fd_sc_hd__inv_2 _17442_ (.A(net6738),
    .Y(_09339_));
 sky130_fd_sc_hd__mux2_1 _17443_ (.A0(_09337_),
    .A1(_09338_),
    .S(_09339_),
    .X(_09340_));
 sky130_fd_sc_hd__clkbuf_1 _17444_ (.A(_09340_),
    .X(_00392_));
 sky130_fd_sc_hd__a22o_1 _17445_ (.A1(net6741),
    .A2(net7376),
    .B1(net6744),
    .B2(net6738),
    .X(_09341_));
 sky130_fd_sc_hd__or2_1 _17446_ (.A(net6738),
    .B(net6744),
    .X(_09342_));
 sky130_fd_sc_hd__nand2_1 _17447_ (.A(_09341_),
    .B(_09342_),
    .Y(_09343_));
 sky130_fd_sc_hd__xnor2_1 _17448_ (.A(net6743),
    .B(_09343_),
    .Y(_09344_));
 sky130_fd_sc_hd__o21ai_1 _17449_ (.A1(net3274),
    .A2(_09344_),
    .B1(net6656),
    .Y(_09345_));
 sky130_fd_sc_hd__nor2_1 _17450_ (.A(net6736),
    .B(net2577),
    .Y(_09346_));
 sky130_fd_sc_hd__a22o_1 _17451_ (.A1(net6736),
    .A2(_09345_),
    .B1(_09346_),
    .B2(_09344_),
    .X(_00393_));
 sky130_fd_sc_hd__a31o_1 _17452_ (.A1(net6743),
    .A2(_09341_),
    .A3(_09342_),
    .B1(net6736),
    .X(_09347_));
 sky130_fd_sc_hd__a21o_1 _17453_ (.A1(_09341_),
    .A2(_09342_),
    .B1(net6743),
    .X(_09348_));
 sky130_fd_sc_hd__nand2_1 _17454_ (.A(_09347_),
    .B(_09348_),
    .Y(_09349_));
 sky130_fd_sc_hd__xnor2_1 _17455_ (.A(\svm0.delta[3] ),
    .B(_09349_),
    .Y(_09350_));
 sky130_fd_sc_hd__o21ai_1 _17456_ (.A1(net3274),
    .A2(_09350_),
    .B1(net6662),
    .Y(_09351_));
 sky130_fd_sc_hd__nor2_1 _17457_ (.A(\svm0.counter[3] ),
    .B(net2577),
    .Y(_09352_));
 sky130_fd_sc_hd__a22o_1 _17458_ (.A1(\svm0.counter[3] ),
    .A2(_09351_),
    .B1(_09352_),
    .B2(_09350_),
    .X(_00394_));
 sky130_fd_sc_hd__a31o_1 _17459_ (.A1(\svm0.delta[3] ),
    .A2(_09347_),
    .A3(_09348_),
    .B1(\svm0.counter[3] ),
    .X(_09353_));
 sky130_fd_sc_hd__a21bo_1 _17460_ (.A1(_09281_),
    .A2(_09349_),
    .B1_N(_09353_),
    .X(_09354_));
 sky130_fd_sc_hd__xnor2_1 _17461_ (.A(\svm0.delta[4] ),
    .B(_09354_),
    .Y(_09355_));
 sky130_fd_sc_hd__o21ai_1 _17462_ (.A1(net3273),
    .A2(_09355_),
    .B1(net6661),
    .Y(_09356_));
 sky130_fd_sc_hd__nor2_1 _17463_ (.A(\svm0.counter[4] ),
    .B(net2577),
    .Y(_09357_));
 sky130_fd_sc_hd__a22o_1 _17464_ (.A1(\svm0.counter[4] ),
    .A2(_09356_),
    .B1(_09357_),
    .B2(_09355_),
    .X(_00395_));
 sky130_fd_sc_hd__inv_2 _17465_ (.A(\svm0.counter[4] ),
    .Y(_09358_));
 sky130_fd_sc_hd__a21o_1 _17466_ (.A1(_09287_),
    .A2(_09354_),
    .B1(net4008),
    .X(_09359_));
 sky130_fd_sc_hd__o21a_1 _17467_ (.A1(_09287_),
    .A2(_09354_),
    .B1(_09359_),
    .X(_09360_));
 sky130_fd_sc_hd__and2_1 _17468_ (.A(net4014),
    .B(_09360_),
    .X(_09361_));
 sky130_fd_sc_hd__nor2_1 _17469_ (.A(net4014),
    .B(_09360_),
    .Y(_09362_));
 sky130_fd_sc_hd__nor2_1 _17470_ (.A(_09361_),
    .B(_09362_),
    .Y(_09363_));
 sky130_fd_sc_hd__o21a_1 _17471_ (.A1(net3273),
    .A2(_09363_),
    .B1(net6661),
    .X(_09364_));
 sky130_fd_sc_hd__nor2_1 _17472_ (.A(net4020),
    .B(_09364_),
    .Y(_09365_));
 sky130_fd_sc_hd__a31o_1 _17473_ (.A1(net4020),
    .A2(net2569),
    .A3(_09363_),
    .B1(_09365_),
    .X(_00396_));
 sky130_fd_sc_hd__nand2_1 _17474_ (.A(net4014),
    .B(_09360_),
    .Y(_09366_));
 sky130_fd_sc_hd__a21oi_2 _17475_ (.A1(net6729),
    .A2(_09366_),
    .B1(_09362_),
    .Y(_09367_));
 sky130_fd_sc_hd__xnor2_1 _17476_ (.A(\svm0.delta[6] ),
    .B(_09367_),
    .Y(_09368_));
 sky130_fd_sc_hd__o21ai_1 _17477_ (.A1(net3273),
    .A2(_09368_),
    .B1(net6661),
    .Y(_09369_));
 sky130_fd_sc_hd__nor2_1 _17478_ (.A(net6718),
    .B(net2576),
    .Y(_09370_));
 sky130_fd_sc_hd__a22o_1 _17479_ (.A1(net6718),
    .A2(_09369_),
    .B1(_09370_),
    .B2(_09368_),
    .X(_00397_));
 sky130_fd_sc_hd__o21ba_1 _17480_ (.A1(_09295_),
    .A2(_09367_),
    .B1_N(net6718),
    .X(_09371_));
 sky130_fd_sc_hd__a21o_1 _17481_ (.A1(_09295_),
    .A2(_09367_),
    .B1(_09371_),
    .X(_09372_));
 sky130_fd_sc_hd__xnor2_1 _17482_ (.A(\svm0.delta[7] ),
    .B(_09372_),
    .Y(_09373_));
 sky130_fd_sc_hd__o21ai_1 _17483_ (.A1(net3273),
    .A2(_09373_),
    .B1(net6661),
    .Y(_09374_));
 sky130_fd_sc_hd__nor2_1 _17484_ (.A(net6717),
    .B(net2576),
    .Y(_09375_));
 sky130_fd_sc_hd__a22o_1 _17485_ (.A1(net6717),
    .A2(_09374_),
    .B1(_09375_),
    .B2(_09373_),
    .X(_00398_));
 sky130_fd_sc_hd__inv_2 _17486_ (.A(net6717),
    .Y(_09376_));
 sky130_fd_sc_hd__o21a_1 _17487_ (.A1(_09299_),
    .A2(_09372_),
    .B1(net4005),
    .X(_09377_));
 sky130_fd_sc_hd__a21o_1 _17488_ (.A1(_09299_),
    .A2(_09372_),
    .B1(_09377_),
    .X(_09378_));
 sky130_fd_sc_hd__xnor2_1 _17489_ (.A(\svm0.delta[8] ),
    .B(net770),
    .Y(_09379_));
 sky130_fd_sc_hd__o21a_1 _17490_ (.A1(net2574),
    .A2(_09379_),
    .B1(net6660),
    .X(_09380_));
 sky130_fd_sc_hd__nor2_1 _17491_ (.A(net4027),
    .B(_09380_),
    .Y(_09381_));
 sky130_fd_sc_hd__a31o_1 _17492_ (.A1(net4027),
    .A2(net2567),
    .A3(_09379_),
    .B1(_09381_),
    .X(_00399_));
 sky130_fd_sc_hd__o21a_1 _17493_ (.A1(_09303_),
    .A2(net770),
    .B1(net4027),
    .X(_09382_));
 sky130_fd_sc_hd__a21o_1 _17494_ (.A1(_09303_),
    .A2(net770),
    .B1(_09382_),
    .X(_09383_));
 sky130_fd_sc_hd__xnor2_1 _17495_ (.A(\svm0.delta[9] ),
    .B(_09383_),
    .Y(_09384_));
 sky130_fd_sc_hd__o21ai_1 _17496_ (.A1(net3275),
    .A2(_09384_),
    .B1(net6660),
    .Y(_09385_));
 sky130_fd_sc_hd__nor2_1 _17497_ (.A(net6705),
    .B(net2579),
    .Y(_09386_));
 sky130_fd_sc_hd__a22o_1 _17498_ (.A1(net6705),
    .A2(_09385_),
    .B1(_09386_),
    .B2(_09384_),
    .X(_00400_));
 sky130_fd_sc_hd__o21ba_1 _17499_ (.A1(_09307_),
    .A2(_09383_),
    .B1_N(net6705),
    .X(_09387_));
 sky130_fd_sc_hd__a21o_1 _17500_ (.A1(_09307_),
    .A2(_09383_),
    .B1(_09387_),
    .X(_09388_));
 sky130_fd_sc_hd__xnor2_1 _17501_ (.A(\svm0.delta[10] ),
    .B(_09388_),
    .Y(_09389_));
 sky130_fd_sc_hd__o21a_1 _17502_ (.A1(net4067),
    .A2(_09389_),
    .B1(net6659),
    .X(_09390_));
 sky130_fd_sc_hd__nor2_1 _17503_ (.A(_09258_),
    .B(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__a31o_1 _17504_ (.A1(_09258_),
    .A2(net2571),
    .A3(_09389_),
    .B1(_09391_),
    .X(_00401_));
 sky130_fd_sc_hd__inv_2 _17505_ (.A(net6703),
    .Y(_09392_));
 sky130_fd_sc_hd__clkbuf_2 _17506_ (.A(_09392_),
    .X(_09393_));
 sky130_fd_sc_hd__o21a_1 _17507_ (.A1(_09311_),
    .A2(_09388_),
    .B1(net4016),
    .X(_09394_));
 sky130_fd_sc_hd__a21o_1 _17508_ (.A1(_09311_),
    .A2(_09388_),
    .B1(_09394_),
    .X(_09395_));
 sky130_fd_sc_hd__xnor2_1 _17509_ (.A(\svm0.delta[11] ),
    .B(_09395_),
    .Y(_09396_));
 sky130_fd_sc_hd__o21a_1 _17510_ (.A1(net4067),
    .A2(_09396_),
    .B1(net6659),
    .X(_09397_));
 sky130_fd_sc_hd__nor2_1 _17511_ (.A(net3271),
    .B(_09397_),
    .Y(_09398_));
 sky130_fd_sc_hd__a31o_1 _17512_ (.A1(net3271),
    .A2(net2571),
    .A3(_09396_),
    .B1(_09398_),
    .X(_00402_));
 sky130_fd_sc_hd__o21a_1 _17513_ (.A1(_09315_),
    .A2(_09395_),
    .B1(net3271),
    .X(_09399_));
 sky130_fd_sc_hd__a21o_1 _17514_ (.A1(_09315_),
    .A2(_09395_),
    .B1(_09399_),
    .X(_09400_));
 sky130_fd_sc_hd__xnor2_1 _17515_ (.A(\svm0.delta[12] ),
    .B(_09400_),
    .Y(_09401_));
 sky130_fd_sc_hd__o21ai_1 _17516_ (.A1(net3275),
    .A2(_09401_),
    .B1(net6657),
    .Y(_09402_));
 sky130_fd_sc_hd__nor2_1 _17517_ (.A(net6697),
    .B(_09272_),
    .Y(_09403_));
 sky130_fd_sc_hd__a22o_1 _17518_ (.A1(net6697),
    .A2(_09402_),
    .B1(_09403_),
    .B2(_09401_),
    .X(_00403_));
 sky130_fd_sc_hd__o21ba_1 _17519_ (.A1(_09319_),
    .A2(_09400_),
    .B1_N(net6697),
    .X(_09404_));
 sky130_fd_sc_hd__a21oi_2 _17520_ (.A1(_09319_),
    .A2(_09400_),
    .B1(_09404_),
    .Y(_09405_));
 sky130_fd_sc_hd__xor2_1 _17521_ (.A(net6742),
    .B(_09405_),
    .X(_09406_));
 sky130_fd_sc_hd__o21ai_1 _17522_ (.A1(_09332_),
    .A2(_09406_),
    .B1(net6657),
    .Y(_09407_));
 sky130_fd_sc_hd__nor2_1 _17523_ (.A(net6694),
    .B(_09272_),
    .Y(_09408_));
 sky130_fd_sc_hd__a22o_1 _17524_ (.A1(net6694),
    .A2(_09407_),
    .B1(_09408_),
    .B2(_09406_),
    .X(_00404_));
 sky130_fd_sc_hd__a21o_1 _17525_ (.A1(net6742),
    .A2(_09405_),
    .B1(net6694),
    .X(_09409_));
 sky130_fd_sc_hd__o21a_1 _17526_ (.A1(net6742),
    .A2(_09405_),
    .B1(_09409_),
    .X(_09410_));
 sky130_fd_sc_hd__xnor2_1 _17527_ (.A(\svm0.delta[14] ),
    .B(_09410_),
    .Y(_09411_));
 sky130_fd_sc_hd__a21o_1 _17528_ (.A1(net4253),
    .A2(_09411_),
    .B1(net3388),
    .X(_09412_));
 sky130_fd_sc_hd__or3_1 _17529_ (.A(net6686),
    .B(_09268_),
    .C(_09411_),
    .X(_09413_));
 sky130_fd_sc_hd__a21bo_1 _17530_ (.A1(net6686),
    .A2(_09412_),
    .B1_N(_09413_),
    .X(_00405_));
 sky130_fd_sc_hd__o221a_1 _17531_ (.A1(net6694),
    .A2(net6742),
    .B1(\svm0.delta[14] ),
    .B2(net6686),
    .C1(_09405_),
    .X(_09414_));
 sky130_fd_sc_hd__o211a_1 _17532_ (.A1(net6686),
    .A2(\svm0.delta[14] ),
    .B1(net6742),
    .C1(net6694),
    .X(_09415_));
 sky130_fd_sc_hd__a211o_1 _17533_ (.A1(net6686),
    .A2(\svm0.delta[14] ),
    .B1(_09414_),
    .C1(_09415_),
    .X(_09416_));
 sky130_fd_sc_hd__xnor2_1 _17534_ (.A(\svm0.delta[15] ),
    .B(_09416_),
    .Y(_09417_));
 sky130_fd_sc_hd__a21o_1 _17535_ (.A1(net4253),
    .A2(_09417_),
    .B1(net3388),
    .X(_09418_));
 sky130_fd_sc_hd__or3_1 _17536_ (.A(\svm0.counter[15] ),
    .B(_09268_),
    .C(_09417_),
    .X(_09419_));
 sky130_fd_sc_hd__a21bo_1 _17537_ (.A1(net9041),
    .A2(_09418_),
    .B1_N(_09419_),
    .X(_00406_));
 sky130_fd_sc_hd__xor2_1 _17538_ (.A(net6685),
    .B(\svm0.tC[15] ),
    .X(_09420_));
 sky130_fd_sc_hd__inv_2 _17539_ (.A(\svm0.tC[13] ),
    .Y(_09421_));
 sky130_fd_sc_hd__and2b_1 _17540_ (.A_N(net6687),
    .B(\svm0.tC[14] ),
    .X(_09422_));
 sky130_fd_sc_hd__and2b_1 _17541_ (.A_N(\svm0.tC[14] ),
    .B(net6687),
    .X(_09423_));
 sky130_fd_sc_hd__a211o_1 _17542_ (.A1(net6691),
    .A2(_09421_),
    .B1(_09422_),
    .C1(_09423_),
    .X(_09424_));
 sky130_fd_sc_hd__inv_2 _17543_ (.A(\svm0.tC[12] ),
    .Y(_09425_));
 sky130_fd_sc_hd__inv_2 _17544_ (.A(net6692),
    .Y(_09426_));
 sky130_fd_sc_hd__o2bb2a_1 _17545_ (.A1_N(_09426_),
    .A2_N(\svm0.tC[13] ),
    .B1(_09425_),
    .B2(net6698),
    .X(_09427_));
 sky130_fd_sc_hd__a21bo_1 _17546_ (.A1(net6698),
    .A2(_09425_),
    .B1_N(_09427_),
    .X(_09428_));
 sky130_fd_sc_hd__nor3_1 _17547_ (.A(_09420_),
    .B(_09424_),
    .C(_09428_),
    .Y(_09429_));
 sky130_fd_sc_hd__and2b_1 _17548_ (.A_N(net6722),
    .B(\svm0.tC[6] ),
    .X(_09430_));
 sky130_fd_sc_hd__and2b_1 _17549_ (.A_N(\svm0.tC[6] ),
    .B(net6722),
    .X(_09431_));
 sky130_fd_sc_hd__nor2_1 _17550_ (.A(_09430_),
    .B(_09431_),
    .Y(_09432_));
 sky130_fd_sc_hd__o221a_1 _17551_ (.A1(net4006),
    .A2(\svm0.tC[7] ),
    .B1(\svm0.tC[5] ),
    .B2(_09230_),
    .C1(_09432_),
    .X(_09433_));
 sky130_fd_sc_hd__a21bo_1 _17552_ (.A1(net4006),
    .A2(\svm0.tC[7] ),
    .B1_N(_09433_),
    .X(_09434_));
 sky130_fd_sc_hd__inv_2 _17553_ (.A(\svm0.tC[5] ),
    .Y(_09435_));
 sky130_fd_sc_hd__o2bb2a_1 _17554_ (.A1_N(\svm0.tC[4] ),
    .A2_N(net4010),
    .B1(net6728),
    .B2(_09435_),
    .X(_09436_));
 sky130_fd_sc_hd__o22a_1 _17555_ (.A1(net4009),
    .A2(\svm0.tC[4] ),
    .B1(\svm0.tC[3] ),
    .B2(net4019),
    .X(_09437_));
 sky130_fd_sc_hd__and3b_1 _17556_ (.A_N(_09434_),
    .B(_09436_),
    .C(_09437_),
    .X(_09438_));
 sky130_fd_sc_hd__and2_1 _17557_ (.A(net3278),
    .B(\svm0.tC[10] ),
    .X(_09439_));
 sky130_fd_sc_hd__nor2_1 _17558_ (.A(net3278),
    .B(\svm0.tC[10] ),
    .Y(_09440_));
 sky130_fd_sc_hd__or2_1 _17559_ (.A(_09439_),
    .B(_09440_),
    .X(_09441_));
 sky130_fd_sc_hd__inv_2 _17560_ (.A(\svm0.tC[9] ),
    .Y(_09442_));
 sky130_fd_sc_hd__a2bb2o_1 _17561_ (.A1_N(_09393_),
    .A2_N(\svm0.tC[11] ),
    .B1(_09442_),
    .B2(net6706),
    .X(_09443_));
 sky130_fd_sc_hd__a211o_1 _17562_ (.A1(_09393_),
    .A2(\svm0.tC[11] ),
    .B1(_09441_),
    .C1(_09443_),
    .X(_09444_));
 sky130_fd_sc_hd__xnor2_1 _17563_ (.A(net6712),
    .B(\svm0.tC[8] ),
    .Y(_09445_));
 sky130_fd_sc_hd__inv_2 _17564_ (.A(\svm0.tC[1] ),
    .Y(_09446_));
 sky130_fd_sc_hd__and2_1 _17565_ (.A(net6739),
    .B(\svm0.tC[0] ),
    .X(_09447_));
 sky130_fd_sc_hd__nor2_1 _17566_ (.A(net6739),
    .B(\svm0.tC[0] ),
    .Y(_09448_));
 sky130_fd_sc_hd__or2_1 _17567_ (.A(net6706),
    .B(_09442_),
    .X(_09449_));
 sky130_fd_sc_hd__o221a_1 _17568_ (.A1(net6737),
    .A2(_09446_),
    .B1(_09447_),
    .B2(_09448_),
    .C1(_09449_),
    .X(_09450_));
 sky130_fd_sc_hd__inv_2 _17569_ (.A(net6734),
    .Y(_09451_));
 sky130_fd_sc_hd__a22o_1 _17570_ (.A1(net4019),
    .A2(\svm0.tC[3] ),
    .B1(\svm0.tC[2] ),
    .B2(net4003),
    .X(_09452_));
 sky130_fd_sc_hd__o22a_1 _17571_ (.A1(net4003),
    .A2(\svm0.tC[2] ),
    .B1(\svm0.tC[1] ),
    .B2(net4012),
    .X(_09453_));
 sky130_fd_sc_hd__and2b_1 _17572_ (.A_N(_09452_),
    .B(_09453_),
    .X(_09454_));
 sky130_fd_sc_hd__and4b_1 _17573_ (.A_N(_09444_),
    .B(_09445_),
    .C(_09450_),
    .D(_09454_),
    .X(_09455_));
 sky130_fd_sc_hd__a211o_1 _17574_ (.A1(net4012),
    .A2(\svm0.tC[1] ),
    .B1(\svm0.tC[0] ),
    .C1(net4033),
    .X(_09456_));
 sky130_fd_sc_hd__a21o_1 _17575_ (.A1(_09453_),
    .A2(_09456_),
    .B1(_09452_),
    .X(_09457_));
 sky130_fd_sc_hd__a21o_1 _17576_ (.A1(\svm0.tC[7] ),
    .A2(_09430_),
    .B1(net4006),
    .X(_09458_));
 sky130_fd_sc_hd__or2_1 _17577_ (.A(\svm0.tC[7] ),
    .B(_09430_),
    .X(_09459_));
 sky130_fd_sc_hd__a2bb2o_1 _17578_ (.A1_N(_09434_),
    .A2_N(_09436_),
    .B1(_09458_),
    .B2(_09459_),
    .X(_09460_));
 sky130_fd_sc_hd__a21oi_1 _17579_ (.A1(_09457_),
    .A2(_09438_),
    .B1(_09460_),
    .Y(_09461_));
 sky130_fd_sc_hd__o21ba_1 _17580_ (.A1(net6712),
    .A2(_09461_),
    .B1_N(\svm0.tC[8] ),
    .X(_09462_));
 sky130_fd_sc_hd__a21o_1 _17581_ (.A1(net6712),
    .A2(_09461_),
    .B1(_09462_),
    .X(_09463_));
 sky130_fd_sc_hd__a21oi_1 _17582_ (.A1(_09449_),
    .A2(_09463_),
    .B1(_09444_),
    .Y(_09464_));
 sky130_fd_sc_hd__a31o_1 _17583_ (.A1(net3278),
    .A2(\svm0.tC[11] ),
    .A3(\svm0.tC[10] ),
    .B1(_09393_),
    .X(_09465_));
 sky130_fd_sc_hd__o21a_1 _17584_ (.A1(\svm0.tC[11] ),
    .A2(_09439_),
    .B1(_09465_),
    .X(_09466_));
 sky130_fd_sc_hd__o21ai_1 _17585_ (.A1(net965),
    .A2(_09466_),
    .B1(net2155),
    .Y(_09467_));
 sky130_fd_sc_hd__a21o_1 _17586_ (.A1(\svm0.tC[15] ),
    .A2(_09422_),
    .B1(net4031),
    .X(_09468_));
 sky130_fd_sc_hd__o21ai_1 _17587_ (.A1(\svm0.tC[15] ),
    .A2(_09422_),
    .B1(_09468_),
    .Y(_09469_));
 sky130_fd_sc_hd__o311a_1 _17588_ (.A1(_09420_),
    .A2(_09424_),
    .A3(_09427_),
    .B1(net877),
    .C1(_09469_),
    .X(_09470_));
 sky130_fd_sc_hd__a31o_1 _17589_ (.A1(net2154),
    .A2(net1794),
    .A3(net1460),
    .B1(net820),
    .X(_09471_));
 sky130_fd_sc_hd__a32o_1 _17590_ (.A1(\svm0.calc_ready ),
    .A2(net2568),
    .A3(net769),
    .B1(net9000),
    .B2(net3384),
    .X(_00407_));
 sky130_fd_sc_hd__and2b_1 _17591_ (.A_N(net6689),
    .B(\svm0.tB[14] ),
    .X(_09472_));
 sky130_fd_sc_hd__and2b_1 _17592_ (.A_N(\svm0.tB[14] ),
    .B(net6689),
    .X(_09473_));
 sky130_fd_sc_hd__nor2_1 _17593_ (.A(_09472_),
    .B(_09473_),
    .Y(_09474_));
 sky130_fd_sc_hd__o221a_1 _17594_ (.A1(net4030),
    .A2(\svm0.tB[15] ),
    .B1(\svm0.tB[13] ),
    .B2(_09426_),
    .C1(_09474_),
    .X(_09475_));
 sky130_fd_sc_hd__a21boi_1 _17595_ (.A1(net4030),
    .A2(\svm0.tB[15] ),
    .B1_N(_09475_),
    .Y(_09476_));
 sky130_fd_sc_hd__and2b_1 _17596_ (.A_N(net6721),
    .B(\svm0.tB[6] ),
    .X(_09477_));
 sky130_fd_sc_hd__and2b_1 _17597_ (.A_N(\svm0.tB[6] ),
    .B(net6721),
    .X(_09478_));
 sky130_fd_sc_hd__nor2_1 _17598_ (.A(_09477_),
    .B(_09478_),
    .Y(_09479_));
 sky130_fd_sc_hd__o221a_1 _17599_ (.A1(net4006),
    .A2(\svm0.tB[7] ),
    .B1(\svm0.tB[5] ),
    .B2(net4023),
    .C1(_09479_),
    .X(_09480_));
 sky130_fd_sc_hd__a21boi_1 _17600_ (.A1(net4006),
    .A2(\svm0.tB[7] ),
    .B1_N(_09480_),
    .Y(_09481_));
 sky130_fd_sc_hd__o221a_1 _17601_ (.A1(net4009),
    .A2(\svm0.tB[4] ),
    .B1(\svm0.tB[3] ),
    .B2(net4018),
    .C1(_09481_),
    .X(_09482_));
 sky130_fd_sc_hd__and2_1 _17602_ (.A(net4015),
    .B(\svm0.tB[10] ),
    .X(_09483_));
 sky130_fd_sc_hd__nor2_1 _17603_ (.A(net4015),
    .B(\svm0.tB[10] ),
    .Y(_09484_));
 sky130_fd_sc_hd__or2_1 _17604_ (.A(_09483_),
    .B(_09484_),
    .X(_09485_));
 sky130_fd_sc_hd__inv_2 _17605_ (.A(\svm0.tB[9] ),
    .Y(_09486_));
 sky130_fd_sc_hd__a2bb2o_1 _17606_ (.A1_N(_09392_),
    .A2_N(\svm0.tB[11] ),
    .B1(_09486_),
    .B2(net6706),
    .X(_09487_));
 sky130_fd_sc_hd__a211o_1 _17607_ (.A1(_09393_),
    .A2(\svm0.tB[11] ),
    .B1(_09485_),
    .C1(_09487_),
    .X(_09488_));
 sky130_fd_sc_hd__o2bb2a_1 _17608_ (.A1_N(\svm0.tB[8] ),
    .A2_N(net4025),
    .B1(net6706),
    .B2(_09486_),
    .X(_09489_));
 sky130_fd_sc_hd__inv_2 _17609_ (.A(net6747),
    .Y(_09490_));
 sky130_fd_sc_hd__xnor2_1 _17610_ (.A(net6701),
    .B(\svm0.tB[12] ),
    .Y(_09491_));
 sky130_fd_sc_hd__o221a_1 _17611_ (.A1(net6695),
    .A2(_09490_),
    .B1(\svm0.tB[8] ),
    .B2(net4025),
    .C1(_09491_),
    .X(_09492_));
 sky130_fd_sc_hd__and3b_1 _17612_ (.A_N(_09488_),
    .B(_09489_),
    .C(_09492_),
    .X(_09493_));
 sky130_fd_sc_hd__a22o_1 _17613_ (.A1(net4023),
    .A2(\svm0.tB[5] ),
    .B1(\svm0.tB[4] ),
    .B2(net4009),
    .X(_09494_));
 sky130_fd_sc_hd__or2_1 _17614_ (.A(net6734),
    .B(\svm0.tB[2] ),
    .X(_09495_));
 sky130_fd_sc_hd__nand2_1 _17615_ (.A(net6734),
    .B(\svm0.tB[2] ),
    .Y(_09496_));
 sky130_fd_sc_hd__nand2_1 _17616_ (.A(net6739),
    .B(\svm0.tB[0] ),
    .Y(_09497_));
 sky130_fd_sc_hd__or2_1 _17617_ (.A(net6739),
    .B(\svm0.tB[0] ),
    .X(_09498_));
 sky130_fd_sc_hd__a22o_1 _17618_ (.A1(_09495_),
    .A2(_09496_),
    .B1(_09497_),
    .B2(_09498_),
    .X(_09499_));
 sky130_fd_sc_hd__and2_1 _17619_ (.A(net4012),
    .B(\svm0.tB[1] ),
    .X(_09500_));
 sky130_fd_sc_hd__a21oi_1 _17620_ (.A1(net4018),
    .A2(\svm0.tB[3] ),
    .B1(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__or2_1 _17621_ (.A(net4012),
    .B(\svm0.tB[1] ),
    .X(_09502_));
 sky130_fd_sc_hd__and4bb_1 _17622_ (.A_N(_09494_),
    .B_N(_09499_),
    .C(_09501_),
    .D(_09502_),
    .X(_09503_));
 sky130_fd_sc_hd__o21a_1 _17623_ (.A1(net4033),
    .A2(\svm0.tB[0] ),
    .B1(_09502_),
    .X(_09504_));
 sky130_fd_sc_hd__o22a_1 _17624_ (.A1(_09451_),
    .A2(\svm0.tB[2] ),
    .B1(_09504_),
    .B2(_09500_),
    .X(_09505_));
 sky130_fd_sc_hd__a221o_1 _17625_ (.A1(net4018),
    .A2(\svm0.tB[3] ),
    .B1(\svm0.tB[2] ),
    .B2(_09451_),
    .C1(_09505_),
    .X(_09506_));
 sky130_fd_sc_hd__a21o_1 _17626_ (.A1(\svm0.tB[7] ),
    .A2(_09477_),
    .B1(net4006),
    .X(_09507_));
 sky130_fd_sc_hd__o21a_1 _17627_ (.A1(\svm0.tB[7] ),
    .A2(_09477_),
    .B1(_09507_),
    .X(_09508_));
 sky130_fd_sc_hd__a221o_1 _17628_ (.A1(_09482_),
    .A2(_09506_),
    .B1(_09494_),
    .B2(_09481_),
    .C1(_09508_),
    .X(_09509_));
 sky130_fd_sc_hd__a31o_1 _17629_ (.A1(net3279),
    .A2(\svm0.tB[11] ),
    .A3(\svm0.tB[10] ),
    .B1(_09393_),
    .X(_09510_));
 sky130_fd_sc_hd__or2_1 _17630_ (.A(\svm0.tB[11] ),
    .B(_09483_),
    .X(_09511_));
 sky130_fd_sc_hd__o2bb2a_1 _17631_ (.A1_N(_09510_),
    .A2_N(_09511_),
    .B1(_09488_),
    .B2(_09489_),
    .X(_09512_));
 sky130_fd_sc_hd__o21ba_1 _17632_ (.A1(net6699),
    .A2(_09512_),
    .B1_N(\svm0.tB[12] ),
    .X(_09513_));
 sky130_fd_sc_hd__a21oi_1 _17633_ (.A1(net6699),
    .A2(_09512_),
    .B1(_09513_),
    .Y(_09514_));
 sky130_fd_sc_hd__a221o_1 _17634_ (.A1(net4004),
    .A2(net6747),
    .B1(net1458),
    .B2(_09493_),
    .C1(_09514_),
    .X(_09515_));
 sky130_fd_sc_hd__a21o_1 _17635_ (.A1(\svm0.tB[15] ),
    .A2(_09472_),
    .B1(net4030),
    .X(_09516_));
 sky130_fd_sc_hd__o21a_1 _17636_ (.A1(\svm0.tB[15] ),
    .A2(_09472_),
    .B1(_09516_),
    .X(_09517_));
 sky130_fd_sc_hd__a21oi_1 _17637_ (.A1(net2153),
    .A2(_09515_),
    .B1(net2566),
    .Y(_09518_));
 sky130_fd_sc_hd__a41o_1 _17638_ (.A1(net2153),
    .A2(net1792),
    .A3(_09493_),
    .A4(net2151),
    .B1(_09518_),
    .X(_09519_));
 sky130_fd_sc_hd__a32o_1 _17639_ (.A1(\svm0.calc_ready ),
    .A2(net2568),
    .A3(net876),
    .B1(net8962),
    .B2(net3384),
    .X(_00408_));
 sky130_fd_sc_hd__and2b_1 _17640_ (.A_N(net6689),
    .B(\svm0.tA[14] ),
    .X(_09520_));
 sky130_fd_sc_hd__and2b_1 _17641_ (.A_N(\svm0.tA[14] ),
    .B(net6688),
    .X(_09521_));
 sky130_fd_sc_hd__or2_1 _17642_ (.A(_09520_),
    .B(_09521_),
    .X(_09522_));
 sky130_fd_sc_hd__nor2_1 _17643_ (.A(net4004),
    .B(\svm0.tA[13] ),
    .Y(_09523_));
 sky130_fd_sc_hd__xor2_1 _17644_ (.A(net6684),
    .B(\svm0.tA[15] ),
    .X(_09524_));
 sky130_fd_sc_hd__xor2_1 _17645_ (.A(net6701),
    .B(\svm0.tA[12] ),
    .X(_09525_));
 sky130_fd_sc_hd__and2_1 _17646_ (.A(net4026),
    .B(\svm0.tA[8] ),
    .X(_09526_));
 sky130_fd_sc_hd__nor2_1 _17647_ (.A(net4026),
    .B(\svm0.tA[8] ),
    .Y(_09527_));
 sky130_fd_sc_hd__nand2_1 _17648_ (.A(net6707),
    .B(net6746),
    .Y(_09528_));
 sky130_fd_sc_hd__or2_1 _17649_ (.A(net6707),
    .B(net6746),
    .X(_09529_));
 sky130_fd_sc_hd__or2_1 _17650_ (.A(net6704),
    .B(\svm0.tA[11] ),
    .X(_09530_));
 sky130_fd_sc_hd__nand2_1 _17651_ (.A(net6704),
    .B(\svm0.tA[11] ),
    .Y(_09531_));
 sky130_fd_sc_hd__a22o_1 _17652_ (.A1(_09528_),
    .A2(_09529_),
    .B1(_09530_),
    .B2(_09531_),
    .X(_09532_));
 sky130_fd_sc_hd__or4_1 _17653_ (.A(_09525_),
    .B(_09526_),
    .C(_09527_),
    .D(_09532_),
    .X(_09533_));
 sky130_fd_sc_hd__or4_1 _17654_ (.A(_09522_),
    .B(_09523_),
    .C(_09524_),
    .D(_09533_),
    .X(_09534_));
 sky130_fd_sc_hd__nand2_1 _17655_ (.A(net3279),
    .B(\svm0.tA[10] ),
    .Y(_09535_));
 sky130_fd_sc_hd__or2_1 _17656_ (.A(net3279),
    .B(\svm0.tA[10] ),
    .X(_09536_));
 sky130_fd_sc_hd__nand2_1 _17657_ (.A(net4004),
    .B(\svm0.tA[13] ),
    .Y(_09537_));
 sky130_fd_sc_hd__and4b_1 _17658_ (.A_N(_09534_),
    .B(_09535_),
    .C(_09536_),
    .D(_09537_),
    .X(_09538_));
 sky130_fd_sc_hd__and2b_1 _17659_ (.A_N(net6723),
    .B(\svm0.tA[6] ),
    .X(_09539_));
 sky130_fd_sc_hd__and2b_1 _17660_ (.A_N(\svm0.tA[6] ),
    .B(net6725),
    .X(_09540_));
 sky130_fd_sc_hd__nor2_1 _17661_ (.A(_09539_),
    .B(_09540_),
    .Y(_09541_));
 sky130_fd_sc_hd__o221a_1 _17662_ (.A1(net4007),
    .A2(\svm0.tA[7] ),
    .B1(\svm0.tA[5] ),
    .B2(net4021),
    .C1(_09541_),
    .X(_09542_));
 sky130_fd_sc_hd__a21boi_1 _17663_ (.A1(net4007),
    .A2(\svm0.tA[7] ),
    .B1_N(_09542_),
    .Y(_09543_));
 sky130_fd_sc_hd__xor2_1 _17664_ (.A(\svm0.counter[3] ),
    .B(\svm0.tA[3] ),
    .X(_09544_));
 sky130_fd_sc_hd__inv_2 _17665_ (.A(\svm0.tA[0] ),
    .Y(_09545_));
 sky130_fd_sc_hd__a2bb2o_1 _17666_ (.A1_N(net4013),
    .A2_N(\svm0.tA[1] ),
    .B1(_09545_),
    .B2(net6740),
    .X(_09546_));
 sky130_fd_sc_hd__a22oi_1 _17667_ (.A1(net4021),
    .A2(\svm0.tA[5] ),
    .B1(\svm0.tA[4] ),
    .B2(net4011),
    .Y(_09547_));
 sky130_fd_sc_hd__xnor2_1 _17668_ (.A(net6735),
    .B(\svm0.tA[2] ),
    .Y(_09548_));
 sky130_fd_sc_hd__and4bb_1 _17669_ (.A_N(_09544_),
    .B_N(_09546_),
    .C(_09547_),
    .D(_09548_),
    .X(_09549_));
 sky130_fd_sc_hd__nand2_1 _17670_ (.A(net4013),
    .B(\svm0.tA[1] ),
    .Y(_09550_));
 sky130_fd_sc_hd__o221a_1 _17671_ (.A1(net4011),
    .A2(\svm0.tA[4] ),
    .B1(_09545_),
    .B2(net6740),
    .C1(_09550_),
    .X(_09551_));
 sky130_fd_sc_hd__nor2_1 _17672_ (.A(net4011),
    .B(\svm0.tA[4] ),
    .Y(_09552_));
 sky130_fd_sc_hd__o2bb2a_1 _17673_ (.A1_N(_09550_),
    .A2_N(_09546_),
    .B1(net4002),
    .B2(\svm0.tA[2] ),
    .X(_09553_));
 sky130_fd_sc_hd__a21o_1 _17674_ (.A1(net4002),
    .A2(\svm0.tA[2] ),
    .B1(_09553_),
    .X(_09554_));
 sky130_fd_sc_hd__o21a_1 _17675_ (.A1(\svm0.tA[3] ),
    .A2(_09554_),
    .B1(_09243_),
    .X(_09555_));
 sky130_fd_sc_hd__a21oi_1 _17676_ (.A1(\svm0.tA[3] ),
    .A2(_09554_),
    .B1(_09555_),
    .Y(_09556_));
 sky130_fd_sc_hd__o21ai_1 _17677_ (.A1(_09552_),
    .A2(_09556_),
    .B1(_09547_),
    .Y(_09557_));
 sky130_fd_sc_hd__a21bo_1 _17678_ (.A1(\svm0.tA[7] ),
    .A2(_09539_),
    .B1_N(\svm0.counter[7] ),
    .X(_09558_));
 sky130_fd_sc_hd__or2_1 _17679_ (.A(\svm0.tA[7] ),
    .B(_09539_),
    .X(_09559_));
 sky130_fd_sc_hd__a22o_1 _17680_ (.A1(_09543_),
    .A2(_09557_),
    .B1(_09558_),
    .B2(_09559_),
    .X(_09560_));
 sky130_fd_sc_hd__nand2_1 _17681_ (.A(net1791),
    .B(_09560_),
    .Y(_09561_));
 sky130_fd_sc_hd__a21o_1 _17682_ (.A1(\svm0.tA[15] ),
    .A2(_09520_),
    .B1(net4030),
    .X(_09562_));
 sky130_fd_sc_hd__o21ai_1 _17683_ (.A1(\svm0.tA[15] ),
    .A2(_09520_),
    .B1(_09562_),
    .Y(_09563_));
 sky130_fd_sc_hd__o21ba_1 _17684_ (.A1(net6746),
    .A2(_09526_),
    .B1_N(net6710),
    .X(_09564_));
 sky130_fd_sc_hd__a221o_1 _17685_ (.A1(net4015),
    .A2(\svm0.tA[10] ),
    .B1(net6746),
    .B2(_09526_),
    .C1(_09564_),
    .X(_09565_));
 sky130_fd_sc_hd__a22o_1 _17686_ (.A1(net3272),
    .A2(\svm0.tA[11] ),
    .B1(_09536_),
    .B2(_09565_),
    .X(_09566_));
 sky130_fd_sc_hd__o21ai_1 _17687_ (.A1(net3272),
    .A2(\svm0.tA[11] ),
    .B1(_09566_),
    .Y(_09567_));
 sky130_fd_sc_hd__o21ba_1 _17688_ (.A1(net6701),
    .A2(_09567_),
    .B1_N(\svm0.tA[12] ),
    .X(_09568_));
 sky130_fd_sc_hd__a21o_1 _17689_ (.A1(net6701),
    .A2(_09567_),
    .B1(_09568_),
    .X(_09569_));
 sky130_fd_sc_hd__a2111o_1 _17690_ (.A1(_09537_),
    .A2(_09569_),
    .B1(_09524_),
    .C1(_09523_),
    .D1(_09522_),
    .X(_09570_));
 sky130_fd_sc_hd__and3_1 _17691_ (.A(_09561_),
    .B(net2565),
    .C(net964),
    .X(_09571_));
 sky130_fd_sc_hd__a41o_1 _17692_ (.A1(net1791),
    .A2(_09543_),
    .A3(_09549_),
    .A4(_09551_),
    .B1(_09571_),
    .X(_09572_));
 sky130_fd_sc_hd__a32o_1 _17693_ (.A1(net9244),
    .A2(net2568),
    .A3(_09572_),
    .B1(net9048),
    .B2(net3384),
    .X(_00409_));
 sky130_fd_sc_hd__o211a_1 _17694_ (.A1(\svm0.state[1] ),
    .A2(net5185),
    .B1(_09187_),
    .C1(net3387),
    .X(_00410_));
 sky130_fd_sc_hd__a21o_1 _17695_ (.A1(net2571),
    .A2(_09202_),
    .B1(net1925),
    .X(_00412_));
 sky130_fd_sc_hd__a21bo_1 _17696_ (.A1(net3389),
    .A2(net1796),
    .B1_N(net6655),
    .X(_09573_));
 sky130_fd_sc_hd__nand2_1 _17697_ (.A(_09204_),
    .B(_09573_),
    .Y(_00413_));
 sky130_fd_sc_hd__or3_1 _17698_ (.A(\pid_q.state[0] ),
    .B(net7521),
    .C(net7463),
    .X(_09574_));
 sky130_fd_sc_hd__clkbuf_1 _17699_ (.A(_09574_),
    .X(_09575_));
 sky130_fd_sc_hd__o21a_1 _17700_ (.A1(net7489),
    .A2(net3270),
    .B1(net8864),
    .X(_09576_));
 sky130_fd_sc_hd__buf_1 _17701_ (.A(_09576_),
    .X(_09577_));
 sky130_fd_sc_hd__or2_1 _17702_ (.A(_04869_),
    .B(_09577_),
    .X(_09578_));
 sky130_fd_sc_hd__clkbuf_1 _17703_ (.A(_09578_),
    .X(_09579_));
 sky130_fd_sc_hd__clkbuf_1 _17704_ (.A(net1455),
    .X(_09580_));
 sky130_fd_sc_hd__inv_2 _17705_ (.A(net7496),
    .Y(_09581_));
 sky130_fd_sc_hd__and4b_1 _17706_ (.A_N(_09576_),
    .B(net8864),
    .C(\pid_q.state[4] ),
    .D(_09581_),
    .X(_09582_));
 sky130_fd_sc_hd__clkbuf_1 _17707_ (.A(_09582_),
    .X(_09583_));
 sky130_fd_sc_hd__clkbuf_1 _17708_ (.A(net1788),
    .X(_09584_));
 sky130_fd_sc_hd__a22o_1 _17709_ (.A1(\pid_q.prev_int[0] ),
    .A2(net1218),
    .B1(net1452),
    .B2(net5184),
    .X(_00414_));
 sky130_fd_sc_hd__a22o_1 _17710_ (.A1(\pid_q.prev_int[1] ),
    .A2(net1218),
    .B1(net1452),
    .B2(net5182),
    .X(_00415_));
 sky130_fd_sc_hd__a22o_1 _17711_ (.A1(\pid_q.prev_int[2] ),
    .A2(net1218),
    .B1(net1452),
    .B2(net5180),
    .X(_00416_));
 sky130_fd_sc_hd__a22o_1 _17712_ (.A1(net9207),
    .A2(net1217),
    .B1(net1451),
    .B2(\pid_q.curr_int[3] ),
    .X(_00417_));
 sky130_fd_sc_hd__a22o_1 _17713_ (.A1(net9239),
    .A2(net1217),
    .B1(net1451),
    .B2(\pid_q.curr_int[4] ),
    .X(_00418_));
 sky130_fd_sc_hd__a22o_1 _17714_ (.A1(net9212),
    .A2(net1219),
    .B1(net1453),
    .B2(\pid_q.curr_int[5] ),
    .X(_00419_));
 sky130_fd_sc_hd__a22o_1 _17715_ (.A1(net9211),
    .A2(net1219),
    .B1(net1453),
    .B2(\pid_q.curr_int[6] ),
    .X(_00420_));
 sky130_fd_sc_hd__a22o_1 _17716_ (.A1(net9221),
    .A2(net1216),
    .B1(net1454),
    .B2(net5178),
    .X(_00421_));
 sky130_fd_sc_hd__a22o_1 _17717_ (.A1(net9200),
    .A2(net1216),
    .B1(net1454),
    .B2(\pid_q.curr_int[8] ),
    .X(_00422_));
 sky130_fd_sc_hd__a22o_1 _17718_ (.A1(net9223),
    .A2(net1216),
    .B1(net1453),
    .B2(\pid_q.curr_int[9] ),
    .X(_00423_));
 sky130_fd_sc_hd__a22o_1 _17719_ (.A1(\pid_q.prev_int[10] ),
    .A2(net1455),
    .B1(net1788),
    .B2(net9202),
    .X(_00424_));
 sky130_fd_sc_hd__a22o_1 _17720_ (.A1(net9201),
    .A2(net1456),
    .B1(net1789),
    .B2(net5177),
    .X(_00425_));
 sky130_fd_sc_hd__a22o_1 _17721_ (.A1(net9185),
    .A2(net1456),
    .B1(net1789),
    .B2(net5175),
    .X(_00426_));
 sky130_fd_sc_hd__a22o_1 _17722_ (.A1(net9125),
    .A2(net1456),
    .B1(net1789),
    .B2(net5173),
    .X(_00427_));
 sky130_fd_sc_hd__a22o_1 _17723_ (.A1(net9189),
    .A2(net1457),
    .B1(net1790),
    .B2(net5170),
    .X(_00428_));
 sky130_fd_sc_hd__a22o_1 _17724_ (.A1(net9122),
    .A2(net1457),
    .B1(net1790),
    .B2(net5169),
    .X(_00429_));
 sky130_fd_sc_hd__nor2_1 _17725_ (.A(net6506),
    .B(net1831),
    .Y(_09585_));
 sky130_fd_sc_hd__mux2_1 _17726_ (.A0(net6506),
    .A1(_09585_),
    .S(net8043),
    .X(_09586_));
 sky130_fd_sc_hd__clkbuf_1 _17727_ (.A(_09586_),
    .X(_00430_));
 sky130_fd_sc_hd__nand2_1 _17728_ (.A(net8059),
    .B(net6522),
    .Y(_09587_));
 sky130_fd_sc_hd__xnor2_1 _17729_ (.A(net6502),
    .B(_09587_),
    .Y(_00431_));
 sky130_fd_sc_hd__nand2_1 _17730_ (.A(net8052),
    .B(net2596),
    .Y(_09588_));
 sky130_fd_sc_hd__xnor2_1 _17731_ (.A(net6475),
    .B(_09588_),
    .Y(_00432_));
 sky130_fd_sc_hd__nor2_1 _17732_ (.A(net2590),
    .B(_09588_),
    .Y(_09589_));
 sky130_fd_sc_hd__xnor2_1 _17733_ (.A(net2599),
    .B(_09589_),
    .Y(_00433_));
 sky130_fd_sc_hd__a31o_1 _17734_ (.A1(net6509),
    .A2(net6457),
    .A3(_08943_),
    .B1(net3668),
    .X(_09590_));
 sky130_fd_sc_hd__and3_1 _17735_ (.A(net8052),
    .B(net6509),
    .C(_08943_),
    .X(_09591_));
 sky130_fd_sc_hd__o2bb2a_1 _17736_ (.A1_N(net8052),
    .A2_N(_09590_),
    .B1(_09591_),
    .B2(net6457),
    .X(_00434_));
 sky130_fd_sc_hd__o21a_1 _17737_ (.A1(net6445),
    .A2(net2881),
    .B1(net6447),
    .X(_09592_));
 sky130_fd_sc_hd__or3_1 _17738_ (.A(net6454),
    .B(_06541_),
    .C(_09592_),
    .X(_09593_));
 sky130_fd_sc_hd__o21ai_1 _17739_ (.A1(_06530_),
    .A2(_06646_),
    .B1(_09593_),
    .Y(_00435_));
 sky130_fd_sc_hd__a21oi_1 _17740_ (.A1(net6443),
    .A2(net6650),
    .B1(net6454),
    .Y(_09594_));
 sky130_fd_sc_hd__o21a_1 _17741_ (.A1(_06536_),
    .A2(_09594_),
    .B1(net6449),
    .X(_09595_));
 sky130_fd_sc_hd__a31o_1 _17742_ (.A1(net4235),
    .A2(net6454),
    .A3(_06646_),
    .B1(_09595_),
    .X(_00436_));
 sky130_fd_sc_hd__o21ai_1 _17743_ (.A1(net6453),
    .A2(net6649),
    .B1(net6449),
    .Y(_09596_));
 sky130_fd_sc_hd__a22o_1 _17744_ (.A1(net5370),
    .A2(_06525_),
    .B1(_09596_),
    .B2(net6443),
    .X(_00437_));
 sky130_fd_sc_hd__o21a_1 _17745_ (.A1(net8998),
    .A2(_08819_),
    .B1(net8060),
    .X(_00438_));
 sky130_fd_sc_hd__nand2_1 _17746_ (.A(net8062),
    .B(net2195),
    .Y(_09597_));
 sky130_fd_sc_hd__buf_1 _17747_ (.A(net1786),
    .X(_09598_));
 sky130_fd_sc_hd__and2b_1 _17748_ (.A_N(net7019),
    .B(net6995),
    .X(_09599_));
 sky130_fd_sc_hd__clkbuf_1 _17749_ (.A(_09599_),
    .X(_09600_));
 sky130_fd_sc_hd__xnor2_2 _17750_ (.A(net6974),
    .B(net3268),
    .Y(_09601_));
 sky130_fd_sc_hd__xor2_4 _17751_ (.A(net6908),
    .B(net6948),
    .X(_09602_));
 sky130_fd_sc_hd__xnor2_2 _17752_ (.A(_09601_),
    .B(_09602_),
    .Y(_09603_));
 sky130_fd_sc_hd__and2b_1 _17753_ (.A_N(net7068),
    .B(net7094),
    .X(_09604_));
 sky130_fd_sc_hd__nand2_1 _17754_ (.A(net7105),
    .B(net3998),
    .Y(_09605_));
 sky130_fd_sc_hd__nor2b_1 _17755_ (.A(net7030),
    .B_N(net7022),
    .Y(_09606_));
 sky130_fd_sc_hd__xnor2_1 _17756_ (.A(net6963),
    .B(net6925),
    .Y(_09607_));
 sky130_fd_sc_hd__or2b_1 _17757_ (.A(net6996),
    .B_N(net7028),
    .X(_09608_));
 sky130_fd_sc_hd__nor2_1 _17758_ (.A(net6996),
    .B(net7021),
    .Y(_09609_));
 sky130_fd_sc_hd__a221o_1 _17759_ (.A1(net6996),
    .A2(net3997),
    .B1(_09607_),
    .B2(_09608_),
    .C1(_09609_),
    .X(_09610_));
 sky130_fd_sc_hd__xor2_1 _17760_ (.A(_09605_),
    .B(_09610_),
    .X(_09611_));
 sky130_fd_sc_hd__xnor2_2 _17761_ (.A(_09603_),
    .B(_09611_),
    .Y(_09612_));
 sky130_fd_sc_hd__or2b_1 _17762_ (.A(net7103),
    .B_N(net7121),
    .X(_09613_));
 sky130_fd_sc_hd__nand2b_1 _17763_ (.A_N(net7121),
    .B(net7133),
    .Y(_09614_));
 sky130_fd_sc_hd__buf_1 _17764_ (.A(_09614_),
    .X(_09615_));
 sky130_fd_sc_hd__o22a_1 _17765_ (.A1(net7135),
    .A2(_09613_),
    .B1(net3265),
    .B2(net3346),
    .X(_09616_));
 sky130_fd_sc_hd__inv_2 _17766_ (.A(net7118),
    .Y(_09617_));
 sky130_fd_sc_hd__a21o_1 _17767_ (.A1(net7092),
    .A2(net3996),
    .B1(net7116),
    .X(_09618_));
 sky130_fd_sc_hd__nand2b_1 _17768_ (.A_N(net7123),
    .B(net7104),
    .Y(_09619_));
 sky130_fd_sc_hd__buf_6 _17769_ (.A(_09619_),
    .X(_09620_));
 sky130_fd_sc_hd__a21boi_1 _17770_ (.A1(net7140),
    .A2(_09618_),
    .B1_N(net3261),
    .Y(_09621_));
 sky130_fd_sc_hd__or2b_1 _17771_ (.A(net7092),
    .B_N(net7116),
    .X(_09622_));
 sky130_fd_sc_hd__or2b_1 _17772_ (.A(net7116),
    .B_N(net7092),
    .X(_09623_));
 sky130_fd_sc_hd__nor2b_1 _17773_ (.A(net7133),
    .B_N(net7120),
    .Y(_09624_));
 sky130_fd_sc_hd__a32o_1 _17774_ (.A1(_09622_),
    .A2(_09623_),
    .A3(net3265),
    .B1(net3994),
    .B2(net7092),
    .X(_09625_));
 sky130_fd_sc_hd__nand2_1 _17775_ (.A(net7061),
    .B(_09625_),
    .Y(_09626_));
 sky130_fd_sc_hd__o221a_1 _17776_ (.A1(net7089),
    .A2(_09616_),
    .B1(_09621_),
    .B2(net7061),
    .C1(_09626_),
    .X(_09627_));
 sky130_fd_sc_hd__xnor2_1 _17777_ (.A(_08985_),
    .B(_09627_),
    .Y(_09628_));
 sky130_fd_sc_hd__xnor2_2 _17778_ (.A(_09612_),
    .B(net1448),
    .Y(_09629_));
 sky130_fd_sc_hd__xnor2_4 _17779_ (.A(net6996),
    .B(net3997),
    .Y(_09630_));
 sky130_fd_sc_hd__xnor2_1 _17780_ (.A(_09630_),
    .B(_09607_),
    .Y(_09631_));
 sky130_fd_sc_hd__and2b_1 _17781_ (.A_N(net7090),
    .B(net7104),
    .X(_09632_));
 sky130_fd_sc_hd__nand2_1 _17782_ (.A(net7119),
    .B(_09632_),
    .Y(_09633_));
 sky130_fd_sc_hd__and2_1 _17783_ (.A(net7023),
    .B(net7030),
    .X(_09634_));
 sky130_fd_sc_hd__xnor2_1 _17784_ (.A(net6986),
    .B(net6942),
    .Y(_09635_));
 sky130_fd_sc_hd__or2b_1 _17785_ (.A(net7006),
    .B_N(net7051),
    .X(_09636_));
 sky130_fd_sc_hd__nor2_1 _17786_ (.A(net7022),
    .B(net7036),
    .Y(_09637_));
 sky130_fd_sc_hd__a221o_1 _17787_ (.A1(net4043),
    .A2(net3993),
    .B1(_09635_),
    .B2(net3992),
    .C1(_09637_),
    .X(_09638_));
 sky130_fd_sc_hd__xnor2_1 _17788_ (.A(net3260),
    .B(net3259),
    .Y(_09639_));
 sky130_fd_sc_hd__xnor2_2 _17789_ (.A(net2563),
    .B(_09639_),
    .Y(_09640_));
 sky130_fd_sc_hd__nor2b_2 _17790_ (.A(net7107),
    .B_N(net7081),
    .Y(_09641_));
 sky130_fd_sc_hd__nand2b_1 _17791_ (.A_N(net7133),
    .B(net7120),
    .Y(_09642_));
 sky130_fd_sc_hd__buf_1 _17792_ (.A(_09642_),
    .X(_09643_));
 sky130_fd_sc_hd__nand2b_1 _17793_ (.A_N(net7108),
    .B(net7136),
    .Y(_09644_));
 sky130_fd_sc_hd__xor2_1 _17794_ (.A(net7108),
    .B(net7133),
    .X(_09645_));
 sky130_fd_sc_hd__mux2_1 _17795_ (.A0(_09644_),
    .A1(_09645_),
    .S(net7082),
    .X(_09646_));
 sky130_fd_sc_hd__o221ai_1 _17796_ (.A1(net3991),
    .A2(_09643_),
    .B1(_09646_),
    .B2(net7120),
    .C1(net7051),
    .Y(_09647_));
 sky130_fd_sc_hd__inv_2 _17797_ (.A(net7095),
    .Y(_09648_));
 sky130_fd_sc_hd__clkbuf_1 _17798_ (.A(_09648_),
    .X(_09649_));
 sky130_fd_sc_hd__nand3b_1 _17799_ (.A_N(net7104),
    .B(net7119),
    .C(net7091),
    .Y(_09650_));
 sky130_fd_sc_hd__a21oi_1 _17800_ (.A1(net3263),
    .A2(_09650_),
    .B1(net7132),
    .Y(_09651_));
 sky130_fd_sc_hd__a311o_1 _17801_ (.A1(net3255),
    .A2(net3258),
    .A3(net3266),
    .B1(_09651_),
    .C1(net7061),
    .X(_09652_));
 sky130_fd_sc_hd__and2_1 _17802_ (.A(net2562),
    .B(_09652_),
    .X(_09653_));
 sky130_fd_sc_hd__and3_1 _17803_ (.A(net7061),
    .B(net3262),
    .C(_09613_),
    .X(_09654_));
 sky130_fd_sc_hd__nor2_1 _17804_ (.A(net7061),
    .B(_09613_),
    .Y(_09655_));
 sky130_fd_sc_hd__o21ai_1 _17805_ (.A1(_09654_),
    .A2(_09655_),
    .B1(net7091),
    .Y(_09656_));
 sky130_fd_sc_hd__or3_1 _17806_ (.A(net7060),
    .B(net7090),
    .C(_09620_),
    .X(_09657_));
 sky130_fd_sc_hd__a21bo_1 _17807_ (.A1(_09656_),
    .A2(_09657_),
    .B1_N(net7132),
    .X(_09658_));
 sky130_fd_sc_hd__o21a_1 _17808_ (.A1(_09640_),
    .A2(_09653_),
    .B1(net1781),
    .X(_09659_));
 sky130_fd_sc_hd__inv_2 _17809_ (.A(net6982),
    .Y(_09660_));
 sky130_fd_sc_hd__nand2_1 _17810_ (.A(net6954),
    .B(net6885),
    .Y(_09661_));
 sky130_fd_sc_hd__or2_1 _17811_ (.A(net3988),
    .B(_09661_),
    .X(_09662_));
 sky130_fd_sc_hd__inv_2 _17812_ (.A(net6856),
    .Y(_09663_));
 sky130_fd_sc_hd__nand2_1 _17813_ (.A(net6974),
    .B(net6925),
    .Y(_09664_));
 sky130_fd_sc_hd__xnor2_2 _17814_ (.A(net3977),
    .B(_09664_),
    .Y(_09665_));
 sky130_fd_sc_hd__xor2_2 _17815_ (.A(net3248),
    .B(_09665_),
    .X(_09666_));
 sky130_fd_sc_hd__or2_1 _17816_ (.A(net3259),
    .B(net2563),
    .X(_09667_));
 sky130_fd_sc_hd__and2_1 _17817_ (.A(net3259),
    .B(net2563),
    .X(_09668_));
 sky130_fd_sc_hd__a21o_1 _17818_ (.A1(net3260),
    .A2(_09667_),
    .B1(_09668_),
    .X(_09669_));
 sky130_fd_sc_hd__nand2_1 _17819_ (.A(_09666_),
    .B(_09669_),
    .Y(_09670_));
 sky130_fd_sc_hd__or2_1 _17820_ (.A(_09666_),
    .B(_09669_),
    .X(_09671_));
 sky130_fd_sc_hd__a22o_1 _17821_ (.A1(_09629_),
    .A2(_09659_),
    .B1(_09670_),
    .B2(_09671_),
    .X(_09672_));
 sky130_fd_sc_hd__o21a_1 _17822_ (.A1(_09629_),
    .A2(_09659_),
    .B1(_09672_),
    .X(_09673_));
 sky130_fd_sc_hd__nor2b_1 _17823_ (.A(net6989),
    .B_N(net6965),
    .Y(_09674_));
 sky130_fd_sc_hd__xnor2_2 _17824_ (.A(net6943),
    .B(_09674_),
    .Y(_09675_));
 sky130_fd_sc_hd__xor2_2 _17825_ (.A(net6926),
    .B(net6875),
    .X(_09676_));
 sky130_fd_sc_hd__xor2_1 _17826_ (.A(net3246),
    .B(_09676_),
    .X(_09677_));
 sky130_fd_sc_hd__inv_2 _17827_ (.A(net2561),
    .Y(_09678_));
 sky130_fd_sc_hd__nand2_1 _17828_ (.A(net7122),
    .B(net7139),
    .Y(_09679_));
 sky130_fd_sc_hd__nand2_1 _17829_ (.A(net7065),
    .B(net7032),
    .Y(_09680_));
 sky130_fd_sc_hd__or2b_1 _17830_ (.A(_09679_),
    .B_N(_09680_),
    .X(_09681_));
 sky130_fd_sc_hd__nor2_1 _17831_ (.A(net7060),
    .B(net7027),
    .Y(_09682_));
 sky130_fd_sc_hd__a221o_1 _17832_ (.A1(net7032),
    .A2(_09679_),
    .B1(_09681_),
    .B2(_09648_),
    .C1(net3974),
    .X(_09683_));
 sky130_fd_sc_hd__and2b_1 _17833_ (.A_N(_09600_),
    .B(_09602_),
    .X(_09684_));
 sky130_fd_sc_hd__or2_1 _17834_ (.A(net6974),
    .B(net6995),
    .X(_09685_));
 sky130_fd_sc_hd__o221a_2 _17835_ (.A1(net7019),
    .A2(_09602_),
    .B1(_09684_),
    .B2(_09051_),
    .C1(_09685_),
    .X(_09686_));
 sky130_fd_sc_hd__xor2_1 _17836_ (.A(net2559),
    .B(_09686_),
    .X(_09687_));
 sky130_fd_sc_hd__xnor2_1 _17837_ (.A(_09678_),
    .B(_09687_),
    .Y(_09688_));
 sky130_fd_sc_hd__and2b_1 _17838_ (.A_N(net7059),
    .B(net7028),
    .X(_09689_));
 sky130_fd_sc_hd__xnor2_2 _17839_ (.A(net7020),
    .B(_09689_),
    .Y(_09690_));
 sky130_fd_sc_hd__xnor2_1 _17840_ (.A(_09648_),
    .B(net3261),
    .Y(_09691_));
 sky130_fd_sc_hd__xnor2_1 _17841_ (.A(_09690_),
    .B(net2558),
    .Y(_09692_));
 sky130_fd_sc_hd__o21a_1 _17842_ (.A1(net7104),
    .A2(_09643_),
    .B1(_09620_),
    .X(_09693_));
 sky130_fd_sc_hd__and2b_1 _17843_ (.A_N(net7103),
    .B(net7123),
    .X(_09694_));
 sky130_fd_sc_hd__nand2_1 _17844_ (.A(net7132),
    .B(_09694_),
    .Y(_09695_));
 sky130_fd_sc_hd__nor2b_1 _17845_ (.A(net7094),
    .B_N(net7068),
    .Y(_09696_));
 sky130_fd_sc_hd__xnor2_2 _17846_ (.A(net7027),
    .B(net3970),
    .Y(_09697_));
 sky130_fd_sc_hd__mux2_1 _17847_ (.A0(_09693_),
    .A1(_09695_),
    .S(_09697_),
    .X(_09698_));
 sky130_fd_sc_hd__xor2_1 _17848_ (.A(net2145),
    .B(net2143),
    .X(_09699_));
 sky130_fd_sc_hd__xnor2_1 _17849_ (.A(_09688_),
    .B(_09699_),
    .Y(_09700_));
 sky130_fd_sc_hd__nor2_1 _17850_ (.A(net7043),
    .B(net3347),
    .Y(_09701_));
 sky130_fd_sc_hd__nand2_1 _17851_ (.A(_09622_),
    .B(net3265),
    .Y(_09702_));
 sky130_fd_sc_hd__and2b_1 _17852_ (.A_N(net7130),
    .B(net7146),
    .X(_09703_));
 sky130_fd_sc_hd__nor2_1 _17853_ (.A(net7043),
    .B(net7111),
    .Y(_09704_));
 sky130_fd_sc_hd__o21a_1 _17854_ (.A1(_09703_),
    .A2(_09704_),
    .B1(net3256),
    .X(_09705_));
 sky130_fd_sc_hd__a221o_1 _17855_ (.A1(net7097),
    .A2(_09701_),
    .B1(_09702_),
    .B2(net7033),
    .C1(_09705_),
    .X(_09706_));
 sky130_fd_sc_hd__or3b_1 _17856_ (.A(net7029),
    .B(net7124),
    .C_N(net7140),
    .X(_09707_));
 sky130_fd_sc_hd__o21ai_1 _17857_ (.A1(_08984_),
    .A2(net7105),
    .B1(_09707_),
    .Y(_09708_));
 sky130_fd_sc_hd__xnor2_1 _17858_ (.A(net7028),
    .B(net7105),
    .Y(_09709_));
 sky130_fd_sc_hd__or3_1 _17859_ (.A(net3971),
    .B(net3258),
    .C(_09709_),
    .X(_09710_));
 sky130_fd_sc_hd__nand2_1 _17860_ (.A(net7091),
    .B(net7027),
    .Y(_09711_));
 sky130_fd_sc_hd__o221ai_1 _17861_ (.A1(net7069),
    .A2(_09709_),
    .B1(_09711_),
    .B2(net7105),
    .C1(net3258),
    .Y(_09712_));
 sky130_fd_sc_hd__a22o_1 _17862_ (.A1(net3998),
    .A2(_09708_),
    .B1(_09710_),
    .B2(_09712_),
    .X(_09713_));
 sky130_fd_sc_hd__a21oi_1 _17863_ (.A1(net7064),
    .A2(net2142),
    .B1(_09713_),
    .Y(_09714_));
 sky130_fd_sc_hd__o21a_1 _17864_ (.A1(_08985_),
    .A2(net3258),
    .B1(_09707_),
    .X(_09715_));
 sky130_fd_sc_hd__or3_1 _17865_ (.A(net4043),
    .B(_09632_),
    .C(net3990),
    .X(_09716_));
 sky130_fd_sc_hd__mux2_1 _17866_ (.A0(_09622_),
    .A1(_09623_),
    .S(_08966_),
    .X(_09717_));
 sky130_fd_sc_hd__mux2_1 _17867_ (.A0(net3258),
    .A1(net3266),
    .S(net7031),
    .X(_09718_));
 sky130_fd_sc_hd__o22a_1 _17868_ (.A1(_09715_),
    .A2(_09716_),
    .B1(_09717_),
    .B2(_09718_),
    .X(_09719_));
 sky130_fd_sc_hd__xnor2_1 _17869_ (.A(_09050_),
    .B(net3268),
    .Y(_09720_));
 sky130_fd_sc_hd__xnor2_1 _17870_ (.A(_09720_),
    .B(_09602_),
    .Y(_09721_));
 sky130_fd_sc_hd__a211o_1 _17871_ (.A1(_09605_),
    .A2(net2141),
    .B1(_09721_),
    .C1(_09610_),
    .X(_09722_));
 sky130_fd_sc_hd__nand2_1 _17872_ (.A(_09605_),
    .B(_09610_),
    .Y(_09723_));
 sky130_fd_sc_hd__nor2_1 _17873_ (.A(_09605_),
    .B(_09610_),
    .Y(_09724_));
 sky130_fd_sc_hd__a21oi_1 _17874_ (.A1(_09723_),
    .A2(_09603_),
    .B1(_09724_),
    .Y(_09725_));
 sky130_fd_sc_hd__nor2_1 _17875_ (.A(_09723_),
    .B(_09603_),
    .Y(_09726_));
 sky130_fd_sc_hd__a22o_1 _17876_ (.A1(_09725_),
    .A2(net1780),
    .B1(net2141),
    .B2(_09726_),
    .X(_09727_));
 sky130_fd_sc_hd__o21ba_1 _17877_ (.A1(net1780),
    .A2(_09722_),
    .B1_N(_09727_),
    .X(_09728_));
 sky130_fd_sc_hd__nand2_1 _17878_ (.A(net6908),
    .B(net6948),
    .Y(_09729_));
 sky130_fd_sc_hd__xor2_1 _17879_ (.A(net6844),
    .B(_09729_),
    .X(_09730_));
 sky130_fd_sc_hd__nor2_1 _17880_ (.A(net3977),
    .B(_09664_),
    .Y(_09731_));
 sky130_fd_sc_hd__xnor2_1 _17881_ (.A(net3245),
    .B(_09731_),
    .Y(_09732_));
 sky130_fd_sc_hd__xnor2_1 _17882_ (.A(_09728_),
    .B(_09732_),
    .Y(_09733_));
 sky130_fd_sc_hd__xor2_1 _17883_ (.A(net1214),
    .B(_09733_),
    .X(_09734_));
 sky130_fd_sc_hd__inv_2 _17884_ (.A(net6873),
    .Y(_09735_));
 sky130_fd_sc_hd__nand2_1 _17885_ (.A(net6994),
    .B(net6947),
    .Y(_09736_));
 sky130_fd_sc_hd__xnor2_1 _17886_ (.A(net3964),
    .B(_09736_),
    .Y(_09737_));
 sky130_fd_sc_hd__nand2_1 _17887_ (.A(net6966),
    .B(net7005),
    .Y(_09738_));
 sky130_fd_sc_hd__or3_1 _17888_ (.A(_09092_),
    .B(net3242),
    .C(_09738_),
    .X(_09739_));
 sky130_fd_sc_hd__xnor2_1 _17889_ (.A(net6966),
    .B(net7005),
    .Y(_09740_));
 sky130_fd_sc_hd__or2b_1 _17890_ (.A(net7027),
    .B_N(net7091),
    .X(_09741_));
 sky130_fd_sc_hd__a221o_1 _17891_ (.A1(net7027),
    .A2(net3970),
    .B1(_09740_),
    .B2(_09741_),
    .C1(_09682_),
    .X(_09742_));
 sky130_fd_sc_hd__xnor2_1 _17892_ (.A(_09690_),
    .B(_09635_),
    .Y(_09743_));
 sky130_fd_sc_hd__a21o_1 _17893_ (.A1(_09742_),
    .A2(net2553),
    .B1(_09695_),
    .X(_09744_));
 sky130_fd_sc_hd__o21a_1 _17894_ (.A1(_09742_),
    .A2(net2553),
    .B1(_09744_),
    .X(_09745_));
 sky130_fd_sc_hd__o21ai_1 _17895_ (.A1(_09093_),
    .A2(_09738_),
    .B1(net3242),
    .Y(_09746_));
 sky130_fd_sc_hd__a21boi_2 _17896_ (.A1(_09739_),
    .A2(_09745_),
    .B1_N(_09746_),
    .Y(_09747_));
 sky130_fd_sc_hd__a21o_1 _17897_ (.A1(net3348),
    .A2(net3969),
    .B1(net3995),
    .X(_09748_));
 sky130_fd_sc_hd__o221a_1 _17898_ (.A1(net7132),
    .A2(net3263),
    .B1(_09748_),
    .B2(net7091),
    .C1(_09650_),
    .X(_09749_));
 sky130_fd_sc_hd__xnor2_1 _17899_ (.A(net7060),
    .B(_09749_),
    .Y(_09750_));
 sky130_fd_sc_hd__xnor2_2 _17900_ (.A(_09640_),
    .B(_09750_),
    .Y(_09751_));
 sky130_fd_sc_hd__xnor2_1 _17901_ (.A(_09695_),
    .B(_09742_),
    .Y(_09752_));
 sky130_fd_sc_hd__xnor2_1 _17902_ (.A(net2553),
    .B(_09752_),
    .Y(_09753_));
 sky130_fd_sc_hd__xnor2_4 _17903_ (.A(net7133),
    .B(net2557),
    .Y(_09754_));
 sky130_fd_sc_hd__nand2b_1 _17904_ (.A_N(_09753_),
    .B(_09754_),
    .Y(_09755_));
 sky130_fd_sc_hd__nor2_1 _17905_ (.A(_09751_),
    .B(_09755_),
    .Y(_09756_));
 sky130_fd_sc_hd__nand2_1 _17906_ (.A(_09746_),
    .B(_09739_),
    .Y(_09757_));
 sky130_fd_sc_hd__xor2_1 _17907_ (.A(_09745_),
    .B(_09757_),
    .X(_09758_));
 sky130_fd_sc_hd__nand2_1 _17908_ (.A(_09751_),
    .B(_09755_),
    .Y(_09759_));
 sky130_fd_sc_hd__o21a_1 _17909_ (.A1(_09756_),
    .A2(_09758_),
    .B1(_09759_),
    .X(_09760_));
 sky130_fd_sc_hd__and2_1 _17910_ (.A(_09747_),
    .B(_09760_),
    .X(_09761_));
 sky130_fd_sc_hd__and3_1 _17911_ (.A(net3260),
    .B(_09653_),
    .C(_09667_),
    .X(_09762_));
 sky130_fd_sc_hd__a21o_1 _17912_ (.A1(net2562),
    .A2(_09652_),
    .B1(net3260),
    .X(_09763_));
 sky130_fd_sc_hd__a21oi_1 _17913_ (.A1(net1781),
    .A2(_09763_),
    .B1(_09667_),
    .Y(_09764_));
 sky130_fd_sc_hd__and3_1 _17914_ (.A(net3260),
    .B(net3259),
    .C(net2563),
    .X(_09765_));
 sky130_fd_sc_hd__a22o_1 _17915_ (.A1(_09653_),
    .A2(_09668_),
    .B1(net1781),
    .B2(_09765_),
    .X(_09766_));
 sky130_fd_sc_hd__o31ai_1 _17916_ (.A1(_09762_),
    .A2(_09764_),
    .A3(_09766_),
    .B1(_09666_),
    .Y(_09767_));
 sky130_fd_sc_hd__or4_1 _17917_ (.A(_09762_),
    .B(_09764_),
    .C(_09766_),
    .D(_09666_),
    .X(_09768_));
 sky130_fd_sc_hd__a21o_1 _17918_ (.A1(_09767_),
    .A2(_09768_),
    .B1(_09629_),
    .X(_09769_));
 sky130_fd_sc_hd__nand3_1 _17919_ (.A(_09629_),
    .B(_09767_),
    .C(_09768_),
    .Y(_09770_));
 sky130_fd_sc_hd__o211a_1 _17920_ (.A1(_09747_),
    .A2(_09760_),
    .B1(_09769_),
    .C1(_09770_),
    .X(_09771_));
 sky130_fd_sc_hd__o21a_1 _17921_ (.A1(_09665_),
    .A2(_09669_),
    .B1(net3248),
    .X(_09772_));
 sky130_fd_sc_hd__a21oi_1 _17922_ (.A1(_09665_),
    .A2(_09669_),
    .B1(_09772_),
    .Y(_09773_));
 sky130_fd_sc_hd__o21a_1 _17923_ (.A1(_09761_),
    .A2(_09771_),
    .B1(_09773_),
    .X(_09774_));
 sky130_fd_sc_hd__or3_1 _17924_ (.A(_09761_),
    .B(_09771_),
    .C(_09773_),
    .X(_09775_));
 sky130_fd_sc_hd__o21ai_1 _17925_ (.A1(_09734_),
    .A2(_09774_),
    .B1(_09775_),
    .Y(_09776_));
 sky130_fd_sc_hd__nor2_1 _17926_ (.A(_09761_),
    .B(_09771_),
    .Y(_09777_));
 sky130_fd_sc_hd__inv_2 _17927_ (.A(_09734_),
    .Y(_09778_));
 sky130_fd_sc_hd__inv_2 _17928_ (.A(_09773_),
    .Y(_09779_));
 sky130_fd_sc_hd__nor2_1 _17929_ (.A(net2145),
    .B(net2143),
    .Y(_09780_));
 sky130_fd_sc_hd__nand2_1 _17930_ (.A(net2145),
    .B(net2143),
    .Y(_09781_));
 sky130_fd_sc_hd__o21ai_1 _17931_ (.A1(_09678_),
    .A2(_09780_),
    .B1(_09781_),
    .Y(_09782_));
 sky130_fd_sc_hd__a2bb2o_1 _17932_ (.A1_N(net2559),
    .A2_N(_09782_),
    .B1(_09780_),
    .B2(_09678_),
    .X(_09783_));
 sky130_fd_sc_hd__nand2_1 _17933_ (.A(net2561),
    .B(net2559),
    .Y(_09784_));
 sky130_fd_sc_hd__o211a_1 _17934_ (.A1(net2561),
    .A2(net2559),
    .B1(net2145),
    .C1(net2143),
    .X(_09785_));
 sky130_fd_sc_hd__o21ba_1 _17935_ (.A1(_09780_),
    .A2(_09784_),
    .B1_N(_09785_),
    .X(_09786_));
 sky130_fd_sc_hd__nor2_1 _17936_ (.A(net2561),
    .B(net2559),
    .Y(_09787_));
 sky130_fd_sc_hd__nand2_1 _17937_ (.A(_09780_),
    .B(_09787_),
    .Y(_09788_));
 sky130_fd_sc_hd__o221a_1 _17938_ (.A1(_09781_),
    .A2(_09784_),
    .B1(_09786_),
    .B2(_09686_),
    .C1(_09788_),
    .X(_09789_));
 sky130_fd_sc_hd__a21bo_1 _17939_ (.A1(_09686_),
    .A2(_09783_),
    .B1_N(_09789_),
    .X(_09790_));
 sky130_fd_sc_hd__nor2b_1 _17940_ (.A(net6970),
    .B_N(net6933),
    .Y(_09791_));
 sky130_fd_sc_hd__xnor2_1 _17941_ (.A(net6916),
    .B(_09791_),
    .Y(_09792_));
 sky130_fd_sc_hd__xor2_2 _17942_ (.A(net6912),
    .B(net6851),
    .X(_09793_));
 sky130_fd_sc_hd__xnor2_1 _17943_ (.A(net3240),
    .B(_09793_),
    .Y(_09794_));
 sky130_fd_sc_hd__inv_2 _17944_ (.A(net6941),
    .Y(_09795_));
 sky130_fd_sc_hd__nor2_1 _17945_ (.A(net6978),
    .B(net6951),
    .Y(_09796_));
 sky130_fd_sc_hd__o21bai_1 _17946_ (.A1(net3956),
    .A2(_09676_),
    .B1_N(_09796_),
    .Y(_09797_));
 sky130_fd_sc_hd__nand2_1 _17947_ (.A(net6978),
    .B(net6951),
    .Y(_09798_));
 sky130_fd_sc_hd__a21oi_1 _17948_ (.A1(_09798_),
    .A2(_09676_),
    .B1(net6997),
    .Y(_09799_));
 sky130_fd_sc_hd__nand2_1 _17949_ (.A(net7115),
    .B(net7124),
    .Y(_09800_));
 sky130_fd_sc_hd__a21oi_1 _17950_ (.A1(net7022),
    .A2(_09800_),
    .B1(_09637_),
    .Y(_09801_));
 sky130_fd_sc_hd__o21ai_1 _17951_ (.A1(_09800_),
    .A2(net3993),
    .B1(net4044),
    .Y(_09802_));
 sky130_fd_sc_hd__o211a_1 _17952_ (.A1(_09797_),
    .A2(_09799_),
    .B1(net3239),
    .C1(net3238),
    .X(_09803_));
 sky130_fd_sc_hd__a211oi_1 _17953_ (.A1(net3239),
    .A2(net3238),
    .B1(_09797_),
    .C1(_09799_),
    .Y(_09804_));
 sky130_fd_sc_hd__or3_1 _17954_ (.A(net2552),
    .B(_09803_),
    .C(_09804_),
    .X(_09805_));
 sky130_fd_sc_hd__o21ai_1 _17955_ (.A1(_09803_),
    .A2(_09804_),
    .B1(net2552),
    .Y(_09806_));
 sky130_fd_sc_hd__and2_1 _17956_ (.A(_09805_),
    .B(_09806_),
    .X(_09807_));
 sky130_fd_sc_hd__nand2_1 _17957_ (.A(net7082),
    .B(net7108),
    .Y(_09808_));
 sky130_fd_sc_hd__xnor2_2 _17958_ (.A(net3952),
    .B(_09630_),
    .Y(_09809_));
 sky130_fd_sc_hd__nor2_1 _17959_ (.A(_09696_),
    .B(_09604_),
    .Y(_09810_));
 sky130_fd_sc_hd__xnor2_1 _17960_ (.A(net7141),
    .B(_09810_),
    .Y(_09811_));
 sky130_fd_sc_hd__xnor2_1 _17961_ (.A(_09809_),
    .B(_09811_),
    .Y(_09812_));
 sky130_fd_sc_hd__nor2_1 _17962_ (.A(net7090),
    .B(_09620_),
    .Y(_09813_));
 sky130_fd_sc_hd__nand2_1 _17963_ (.A(_09690_),
    .B(_09633_),
    .Y(_09814_));
 sky130_fd_sc_hd__o31a_1 _17964_ (.A1(_09690_),
    .A2(net3990),
    .A3(_09813_),
    .B1(_09814_),
    .X(_09815_));
 sky130_fd_sc_hd__xor2_1 _17965_ (.A(_09812_),
    .B(net2139),
    .X(_09816_));
 sky130_fd_sc_hd__xnor2_1 _17966_ (.A(_09807_),
    .B(_09816_),
    .Y(_09817_));
 sky130_fd_sc_hd__a21oi_1 _17967_ (.A1(net6924),
    .A2(net6884),
    .B1(_09157_),
    .Y(_09818_));
 sky130_fd_sc_hd__and3_1 _17968_ (.A(net6924),
    .B(net6884),
    .C(net4036),
    .X(_09819_));
 sky130_fd_sc_hd__o2111a_1 _17969_ (.A1(_09818_),
    .A2(_09819_),
    .B1(net6909),
    .C1(net6946),
    .D1(net6845),
    .X(_09820_));
 sky130_fd_sc_hd__a311o_1 _17970_ (.A1(net6909),
    .A2(net6946),
    .A3(net6845),
    .B1(_09818_),
    .C1(_09819_),
    .X(_09821_));
 sky130_fd_sc_hd__or2b_1 _17971_ (.A(_09820_),
    .B_N(_09821_),
    .X(_09822_));
 sky130_fd_sc_hd__xor2_1 _17972_ (.A(_09817_),
    .B(_09822_),
    .X(_09823_));
 sky130_fd_sc_hd__xnor2_1 _17973_ (.A(_09790_),
    .B(net1213),
    .Y(_09824_));
 sky130_fd_sc_hd__or2_1 _17974_ (.A(net3977),
    .B(_09664_),
    .X(_09825_));
 sky130_fd_sc_hd__and3_1 _17975_ (.A(net3245),
    .B(_09825_),
    .C(net1779),
    .X(_09826_));
 sky130_fd_sc_hd__or2_1 _17976_ (.A(net3245),
    .B(net1779),
    .X(_09827_));
 sky130_fd_sc_hd__a21o_1 _17977_ (.A1(net2141),
    .A2(_09612_),
    .B1(net1780),
    .X(_09828_));
 sky130_fd_sc_hd__or2_1 _17978_ (.A(net1214),
    .B(net1447),
    .X(_09829_));
 sky130_fd_sc_hd__o2bb2a_1 _17979_ (.A1_N(net1214),
    .A2_N(_09826_),
    .B1(_09827_),
    .B2(_09829_),
    .X(_09830_));
 sky130_fd_sc_hd__a211o_1 _17980_ (.A1(net3245),
    .A2(net1779),
    .B1(net1447),
    .C1(net1214),
    .X(_09831_));
 sky130_fd_sc_hd__a21o_1 _17981_ (.A1(net1214),
    .A2(net1447),
    .B1(_09827_),
    .X(_09832_));
 sky130_fd_sc_hd__a21o_1 _17982_ (.A1(_09831_),
    .A2(_09832_),
    .B1(_09825_),
    .X(_09833_));
 sky130_fd_sc_hd__nand2_1 _17983_ (.A(_09825_),
    .B(net1779),
    .Y(_09834_));
 sky130_fd_sc_hd__or2_1 _17984_ (.A(_09825_),
    .B(net1779),
    .X(_09835_));
 sky130_fd_sc_hd__nand2_1 _17985_ (.A(net3245),
    .B(_09835_),
    .Y(_09836_));
 sky130_fd_sc_hd__a21boi_1 _17986_ (.A1(_09834_),
    .A2(_09836_),
    .B1_N(net1215),
    .Y(_09837_));
 sky130_fd_sc_hd__o21ai_1 _17987_ (.A1(_09826_),
    .A2(_09837_),
    .B1(net1447),
    .Y(_09838_));
 sky130_fd_sc_hd__and4_1 _17988_ (.A(net963),
    .B(_09830_),
    .C(_09833_),
    .D(_09838_),
    .X(_09839_));
 sky130_fd_sc_hd__a31oi_1 _17989_ (.A1(_09830_),
    .A2(_09833_),
    .A3(_09838_),
    .B1(net963),
    .Y(_09840_));
 sky130_fd_sc_hd__a311o_1 _17990_ (.A1(_09777_),
    .A2(_09778_),
    .A3(_09779_),
    .B1(_09839_),
    .C1(_09840_),
    .X(_09841_));
 sky130_fd_sc_hd__a21o_1 _17991_ (.A1(_09673_),
    .A2(_09776_),
    .B1(_09841_),
    .X(_09842_));
 sky130_fd_sc_hd__and3_2 _17992_ (.A(net6967),
    .B(net7084),
    .C(net7034),
    .X(_09843_));
 sky130_fd_sc_hd__nand2_1 _17993_ (.A(net6940),
    .B(_09843_),
    .Y(_09844_));
 sky130_fd_sc_hd__inv_2 _17994_ (.A(_09843_),
    .Y(_09845_));
 sky130_fd_sc_hd__nor2_1 _17995_ (.A(net6940),
    .B(_09843_),
    .Y(_09846_));
 sky130_fd_sc_hd__or3b_1 _17996_ (.A(net7004),
    .B(_09846_),
    .C_N(net2555),
    .X(_09847_));
 sky130_fd_sc_hd__a211o_1 _17997_ (.A1(net6940),
    .A2(_09845_),
    .B1(net2555),
    .C1(_09026_),
    .X(_09848_));
 sky130_fd_sc_hd__xnor2_2 _17998_ (.A(net7083),
    .B(net7038),
    .Y(_09849_));
 sky130_fd_sc_hd__and3b_1 _17999_ (.A_N(net7135),
    .B(net7118),
    .C(net7109),
    .X(_09850_));
 sky130_fd_sc_hd__a221o_1 _18000_ (.A1(_08913_),
    .A2(_09617_),
    .B1(_09644_),
    .B2(_09849_),
    .C1(_09850_),
    .X(_09851_));
 sky130_fd_sc_hd__a21o_1 _18001_ (.A1(_09847_),
    .A2(_09848_),
    .B1(net3237),
    .X(_09852_));
 sky130_fd_sc_hd__o311a_1 _18002_ (.A1(_09026_),
    .A2(net6940),
    .A3(_09845_),
    .B1(_09852_),
    .C1(net7050),
    .X(_09853_));
 sky130_fd_sc_hd__xnor2_1 _18003_ (.A(_09026_),
    .B(net2555),
    .Y(_09854_));
 sky130_fd_sc_hd__o311a_1 _18004_ (.A1(net3237),
    .A2(_09846_),
    .A3(_09854_),
    .B1(_09844_),
    .C1(net3337),
    .X(_09855_));
 sky130_fd_sc_hd__o22a_1 _18005_ (.A1(net7004),
    .A2(_09844_),
    .B1(_09853_),
    .B2(_09855_),
    .X(_09856_));
 sky130_fd_sc_hd__nand2_1 _18006_ (.A(net3257),
    .B(_09615_),
    .Y(_09857_));
 sky130_fd_sc_hd__xnor2_2 _18007_ (.A(net6990),
    .B(net7035),
    .Y(_09858_));
 sky130_fd_sc_hd__xnor2_2 _18008_ (.A(_09641_),
    .B(_09858_),
    .Y(_09859_));
 sky130_fd_sc_hd__xnor2_4 _18009_ (.A(net7052),
    .B(_09859_),
    .Y(_09860_));
 sky130_fd_sc_hd__or2b_1 _18010_ (.A(net7051),
    .B_N(net7006),
    .X(_09861_));
 sky130_fd_sc_hd__nand2_1 _18011_ (.A(_09636_),
    .B(_09861_),
    .Y(_09862_));
 sky130_fd_sc_hd__nor2_1 _18012_ (.A(net7082),
    .B(_09617_),
    .Y(_09863_));
 sky130_fd_sc_hd__or2_1 _18013_ (.A(net7082),
    .B(net7108),
    .X(_09864_));
 sky130_fd_sc_hd__o221ai_1 _18014_ (.A1(net7118),
    .A2(_09808_),
    .B1(_09862_),
    .B2(_09863_),
    .C1(_09864_),
    .Y(_09865_));
 sky130_fd_sc_hd__nand2_1 _18015_ (.A(_09860_),
    .B(net2550),
    .Y(_09866_));
 sky130_fd_sc_hd__nor2_1 _18016_ (.A(_09860_),
    .B(net2550),
    .Y(_09867_));
 sky130_fd_sc_hd__a21oi_1 _18017_ (.A1(net2551),
    .A2(_09866_),
    .B1(_09867_),
    .Y(_09868_));
 sky130_fd_sc_hd__xnor2_1 _18018_ (.A(_09697_),
    .B(_09740_),
    .Y(_09869_));
 sky130_fd_sc_hd__nand2b_1 _18019_ (.A_N(net7052),
    .B(net7107),
    .Y(_09870_));
 sky130_fd_sc_hd__nor2_1 _18020_ (.A(net7052),
    .B(net7081),
    .Y(_09871_));
 sky130_fd_sc_hd__a221o_1 _18021_ (.A1(net7052),
    .A2(_09641_),
    .B1(_09858_),
    .B2(_09870_),
    .C1(_09871_),
    .X(_09872_));
 sky130_fd_sc_hd__xnor2_2 _18022_ (.A(net7107),
    .B(_09624_),
    .Y(_09873_));
 sky130_fd_sc_hd__xor2_1 _18023_ (.A(_09872_),
    .B(_09873_),
    .X(_09874_));
 sky130_fd_sc_hd__xnor2_2 _18024_ (.A(net2549),
    .B(_09874_),
    .Y(_09875_));
 sky130_fd_sc_hd__inv_2 _18025_ (.A(net6918),
    .Y(_09876_));
 sky130_fd_sc_hd__nand2_1 _18026_ (.A(net6990),
    .B(net7035),
    .Y(_09877_));
 sky130_fd_sc_hd__xnor2_2 _18027_ (.A(net3949),
    .B(_09877_),
    .Y(_09878_));
 sky130_fd_sc_hd__nand2_1 _18028_ (.A(net7013),
    .B(net6936),
    .Y(_09879_));
 sky130_fd_sc_hd__nor2_1 _18029_ (.A(net4043),
    .B(net3943),
    .Y(_09880_));
 sky130_fd_sc_hd__xnor2_2 _18030_ (.A(_09878_),
    .B(net3235),
    .Y(_09881_));
 sky130_fd_sc_hd__xnor2_1 _18031_ (.A(_09875_),
    .B(_09881_),
    .Y(_09882_));
 sky130_fd_sc_hd__xnor2_2 _18032_ (.A(_09868_),
    .B(_09882_),
    .Y(_09883_));
 sky130_fd_sc_hd__nor2_1 _18033_ (.A(_09856_),
    .B(_09883_),
    .Y(_09884_));
 sky130_fd_sc_hd__xnor2_2 _18034_ (.A(_09862_),
    .B(_09851_),
    .Y(_09885_));
 sky130_fd_sc_hd__xnor2_1 _18035_ (.A(net2556),
    .B(_09885_),
    .Y(_09886_));
 sky130_fd_sc_hd__and2_1 _18036_ (.A(net7131),
    .B(_09886_),
    .X(_09887_));
 sky130_fd_sc_hd__mux2_1 _18037_ (.A0(net2555),
    .A1(net7004),
    .S(net3237),
    .X(_09888_));
 sky130_fd_sc_hd__or2_1 _18038_ (.A(net7050),
    .B(net7004),
    .X(_09889_));
 sky130_fd_sc_hd__mux2_1 _18039_ (.A0(_09889_),
    .A1(_09026_),
    .S(net2555),
    .X(_09890_));
 sky130_fd_sc_hd__o2bb2a_2 _18040_ (.A1_N(net7050),
    .A2_N(_09888_),
    .B1(net3237),
    .B2(_09890_),
    .X(_09891_));
 sky130_fd_sc_hd__xnor2_2 _18041_ (.A(net3963),
    .B(_09843_),
    .Y(_09892_));
 sky130_fd_sc_hd__xnor2_4 _18042_ (.A(_09891_),
    .B(_09892_),
    .Y(_09893_));
 sky130_fd_sc_hd__xor2_2 _18043_ (.A(_09860_),
    .B(net2550),
    .X(_09894_));
 sky130_fd_sc_hd__xnor2_2 _18044_ (.A(net2551),
    .B(_09894_),
    .Y(_09895_));
 sky130_fd_sc_hd__o21ba_1 _18045_ (.A1(_09887_),
    .A2(_09893_),
    .B1_N(_09895_),
    .X(_09896_));
 sky130_fd_sc_hd__a21o_1 _18046_ (.A1(_09887_),
    .A2(_09893_),
    .B1(_09896_),
    .X(_09897_));
 sky130_fd_sc_hd__nand2_1 _18047_ (.A(_09856_),
    .B(_09883_),
    .Y(_09898_));
 sky130_fd_sc_hd__o21a_1 _18048_ (.A1(_09884_),
    .A2(_09897_),
    .B1(_09898_),
    .X(_09899_));
 sky130_fd_sc_hd__xor2_2 _18049_ (.A(_09887_),
    .B(_09895_),
    .X(_09900_));
 sky130_fd_sc_hd__xnor2_4 _18050_ (.A(_09893_),
    .B(_09900_),
    .Y(_09901_));
 sky130_fd_sc_hd__xnor2_2 _18051_ (.A(net7078),
    .B(net7112),
    .Y(_09902_));
 sky130_fd_sc_hd__a22o_1 _18052_ (.A1(net7009),
    .A2(net7128),
    .B1(net3969),
    .B2(_09902_),
    .X(_09903_));
 sky130_fd_sc_hd__nor3_1 _18053_ (.A(net7097),
    .B(net3976),
    .C(_09902_),
    .Y(_09904_));
 sky130_fd_sc_hd__a21oi_2 _18054_ (.A1(net7097),
    .A2(_09903_),
    .B1(_09904_),
    .Y(_09905_));
 sky130_fd_sc_hd__a211o_1 _18055_ (.A1(net3348),
    .A2(net3264),
    .B1(net3994),
    .C1(_08966_),
    .X(_09906_));
 sky130_fd_sc_hd__a211o_1 _18056_ (.A1(_08913_),
    .A2(net3257),
    .B1(net3969),
    .C1(net7062),
    .X(_09907_));
 sky130_fd_sc_hd__nand2_1 _18057_ (.A(_09906_),
    .B(_09907_),
    .Y(_09908_));
 sky130_fd_sc_hd__xnor2_4 _18058_ (.A(net6989),
    .B(net7096),
    .Y(_09909_));
 sky130_fd_sc_hd__nand2_1 _18059_ (.A(net7067),
    .B(net7111),
    .Y(_09910_));
 sky130_fd_sc_hd__xor2_1 _18060_ (.A(_09909_),
    .B(_09910_),
    .X(_09911_));
 sky130_fd_sc_hd__xnor2_1 _18061_ (.A(net3330),
    .B(_09911_),
    .Y(_09912_));
 sky130_fd_sc_hd__xnor2_1 _18062_ (.A(_09908_),
    .B(_09912_),
    .Y(_09913_));
 sky130_fd_sc_hd__xor2_2 _18063_ (.A(_09905_),
    .B(_09913_),
    .X(_09914_));
 sky130_fd_sc_hd__nand2_1 _18064_ (.A(net7087),
    .B(\cordic0.vec[1][1] ),
    .Y(_09915_));
 sky130_fd_sc_hd__xnor2_2 _18065_ (.A(net7007),
    .B(_09915_),
    .Y(_09916_));
 sky130_fd_sc_hd__inv_2 _18066_ (.A(_09916_),
    .Y(_09917_));
 sky130_fd_sc_hd__and3_1 _18067_ (.A(net7041),
    .B(net7112),
    .C(net7134),
    .X(_09918_));
 sky130_fd_sc_hd__a21oi_1 _18068_ (.A1(net3256),
    .A2(net7146),
    .B1(net3994),
    .Y(_09919_));
 sky130_fd_sc_hd__xor2_1 _18069_ (.A(_09902_),
    .B(_09919_),
    .X(_09920_));
 sky130_fd_sc_hd__nor2_1 _18070_ (.A(_09918_),
    .B(_09920_),
    .Y(_09921_));
 sky130_fd_sc_hd__nand2_1 _18071_ (.A(_09918_),
    .B(_09920_),
    .Y(_09922_));
 sky130_fd_sc_hd__o21ai_1 _18072_ (.A1(_09917_),
    .A2(_09921_),
    .B1(_09922_),
    .Y(_09923_));
 sky130_fd_sc_hd__and3_1 _18073_ (.A(_09849_),
    .B(_09906_),
    .C(_09907_),
    .X(_09924_));
 sky130_fd_sc_hd__a21oi_1 _18074_ (.A1(_09906_),
    .A2(_09907_),
    .B1(_09849_),
    .Y(_09925_));
 sky130_fd_sc_hd__or2_1 _18075_ (.A(_09924_),
    .B(_09925_),
    .X(_09926_));
 sky130_fd_sc_hd__xnor2_1 _18076_ (.A(net3987),
    .B(net3942),
    .Y(_09927_));
 sky130_fd_sc_hd__o31a_1 _18077_ (.A1(_09905_),
    .A2(_09924_),
    .A3(_09925_),
    .B1(_09927_),
    .X(_09928_));
 sky130_fd_sc_hd__a21oi_1 _18078_ (.A1(_09905_),
    .A2(_09926_),
    .B1(_09928_),
    .Y(_09929_));
 sky130_fd_sc_hd__nand3_1 _18079_ (.A(_09914_),
    .B(_09923_),
    .C(_09929_),
    .Y(_09930_));
 sky130_fd_sc_hd__xnor2_1 _18080_ (.A(net3306),
    .B(_09711_),
    .Y(_09931_));
 sky130_fd_sc_hd__xnor2_2 _18081_ (.A(_09754_),
    .B(_09885_),
    .Y(_09932_));
 sky130_fd_sc_hd__mux2_1 _18082_ (.A0(net3257),
    .A1(net3264),
    .S(_09849_),
    .X(_09933_));
 sky130_fd_sc_hd__nand2_1 _18083_ (.A(net6984),
    .B(net7066),
    .Y(_09934_));
 sky130_fd_sc_hd__o21a_1 _18084_ (.A1(net7062),
    .A2(_09933_),
    .B1(net3940),
    .X(_09935_));
 sky130_fd_sc_hd__mux2_1 _18085_ (.A0(net3969),
    .A1(net3995),
    .S(_09849_),
    .X(_09936_));
 sky130_fd_sc_hd__nand2_1 _18086_ (.A(net7054),
    .B(_09936_),
    .Y(_09937_));
 sky130_fd_sc_hd__mux2_2 _18087_ (.A0(_09935_),
    .A1(_09937_),
    .S(_08914_),
    .X(_09938_));
 sky130_fd_sc_hd__xnor2_2 _18088_ (.A(_09932_),
    .B(_09938_),
    .Y(_09939_));
 sky130_fd_sc_hd__xnor2_1 _18089_ (.A(net2548),
    .B(_09939_),
    .Y(_09940_));
 sky130_fd_sc_hd__a21oi_1 _18090_ (.A1(_09914_),
    .A2(_09923_),
    .B1(_09929_),
    .Y(_09941_));
 sky130_fd_sc_hd__a21oi_1 _18091_ (.A1(_09930_),
    .A2(_09940_),
    .B1(_09941_),
    .Y(_09942_));
 sky130_fd_sc_hd__nand2_1 _18092_ (.A(_09901_),
    .B(_09942_),
    .Y(_09943_));
 sky130_fd_sc_hd__or2_1 _18093_ (.A(_09932_),
    .B(_09938_),
    .X(_09944_));
 sky130_fd_sc_hd__and2_1 _18094_ (.A(_09932_),
    .B(_09938_),
    .X(_09945_));
 sky130_fd_sc_hd__a21oi_1 _18095_ (.A1(net2548),
    .A2(_09944_),
    .B1(_09945_),
    .Y(_09946_));
 sky130_fd_sc_hd__o21ai_1 _18096_ (.A1(_09901_),
    .A2(_09942_),
    .B1(_09946_),
    .Y(_09947_));
 sky130_fd_sc_hd__xor2_1 _18097_ (.A(_09856_),
    .B(_09883_),
    .X(_09948_));
 sky130_fd_sc_hd__xnor2_1 _18098_ (.A(_09897_),
    .B(_09948_),
    .Y(_09949_));
 sky130_fd_sc_hd__a21oi_1 _18099_ (.A1(_09943_),
    .A2(_09947_),
    .B1(net962),
    .Y(_09950_));
 sky130_fd_sc_hd__xnor2_1 _18100_ (.A(_09754_),
    .B(_09753_),
    .Y(_09951_));
 sky130_fd_sc_hd__or2_1 _18101_ (.A(_09872_),
    .B(_09873_),
    .X(_09952_));
 sky130_fd_sc_hd__and2_1 _18102_ (.A(_09872_),
    .B(_09873_),
    .X(_09953_));
 sky130_fd_sc_hd__a21o_1 _18103_ (.A1(net2549),
    .A2(_09952_),
    .B1(_09953_),
    .X(_09954_));
 sky130_fd_sc_hd__xnor2_1 _18104_ (.A(_09092_),
    .B(_09738_),
    .Y(_09955_));
 sky130_fd_sc_hd__nor2_1 _18105_ (.A(net3949),
    .B(_09877_),
    .Y(_09956_));
 sky130_fd_sc_hd__xnor2_1 _18106_ (.A(net3234),
    .B(_09956_),
    .Y(_09957_));
 sky130_fd_sc_hd__inv_2 _18107_ (.A(_09957_),
    .Y(_09958_));
 sky130_fd_sc_hd__xnor2_1 _18108_ (.A(_09954_),
    .B(_09958_),
    .Y(_09959_));
 sky130_fd_sc_hd__xnor2_1 _18109_ (.A(_09951_),
    .B(_09959_),
    .Y(_09960_));
 sky130_fd_sc_hd__o211ai_1 _18110_ (.A1(_09875_),
    .A2(_09881_),
    .B1(_09894_),
    .C1(net2551),
    .Y(_09961_));
 sky130_fd_sc_hd__o21ai_1 _18111_ (.A1(_09860_),
    .A2(net2550),
    .B1(_09881_),
    .Y(_09962_));
 sky130_fd_sc_hd__or3_1 _18112_ (.A(_09860_),
    .B(net2550),
    .C(_09881_),
    .X(_09963_));
 sky130_fd_sc_hd__a21bo_1 _18113_ (.A1(_09962_),
    .A2(_09963_),
    .B1_N(_09875_),
    .X(_09964_));
 sky130_fd_sc_hd__inv_2 _18114_ (.A(net3235),
    .Y(_09965_));
 sky130_fd_sc_hd__o31ai_1 _18115_ (.A1(_09965_),
    .A2(_09860_),
    .A3(net2550),
    .B1(_09878_),
    .Y(_09966_));
 sky130_fd_sc_hd__o21ai_1 _18116_ (.A1(net3235),
    .A2(_09867_),
    .B1(_09966_),
    .Y(_09967_));
 sky130_fd_sc_hd__a21oi_1 _18117_ (.A1(_09961_),
    .A2(_09964_),
    .B1(_09967_),
    .Y(_09968_));
 sky130_fd_sc_hd__nand3_1 _18118_ (.A(_09967_),
    .B(_09961_),
    .C(_09964_),
    .Y(_09969_));
 sky130_fd_sc_hd__and2b_1 _18119_ (.A_N(_09968_),
    .B(_09969_),
    .X(_09970_));
 sky130_fd_sc_hd__xor2_1 _18120_ (.A(_09960_),
    .B(_09970_),
    .X(_09971_));
 sky130_fd_sc_hd__o21ai_1 _18121_ (.A1(_09899_),
    .A2(_09950_),
    .B1(_09971_),
    .Y(_09972_));
 sky130_fd_sc_hd__a21o_1 _18122_ (.A1(net7089),
    .A2(net3263),
    .B1(_09694_),
    .X(_09973_));
 sky130_fd_sc_hd__nand2_1 _18123_ (.A(net7092),
    .B(_09613_),
    .Y(_09974_));
 sky130_fd_sc_hd__a21oi_1 _18124_ (.A1(net3942),
    .A2(_09974_),
    .B1(net7135),
    .Y(_09975_));
 sky130_fd_sc_hd__a221o_1 _18125_ (.A1(net3255),
    .A2(_09748_),
    .B1(_09973_),
    .B2(net7061),
    .C1(_09975_),
    .X(_09976_));
 sky130_fd_sc_hd__nand2_1 _18126_ (.A(net7038),
    .B(_09976_),
    .Y(_09977_));
 sky130_fd_sc_hd__a21o_1 _18127_ (.A1(_09800_),
    .A2(net3265),
    .B1(net3339),
    .X(_09978_));
 sky130_fd_sc_hd__o211a_1 _18128_ (.A1(net3347),
    .A2(net3265),
    .B1(_09978_),
    .C1(net3256),
    .X(_09979_));
 sky130_fd_sc_hd__o211a_1 _18129_ (.A1(net3339),
    .A2(net3262),
    .B1(net3976),
    .C1(net7092),
    .X(_09980_));
 sky130_fd_sc_hd__o32a_1 _18130_ (.A1(net7033),
    .A2(_09979_),
    .A3(_09980_),
    .B1(_09623_),
    .B2(net3976),
    .X(_09981_));
 sky130_fd_sc_hd__or3b_1 _18131_ (.A(_09916_),
    .B(_09921_),
    .C_N(_09922_),
    .X(_09982_));
 sky130_fd_sc_hd__a21bo_1 _18132_ (.A1(_09916_),
    .A2(_09921_),
    .B1_N(_09982_),
    .X(_09983_));
 sky130_fd_sc_hd__o2bb2a_1 _18133_ (.A1_N(_09914_),
    .A2_N(_09983_),
    .B1(_09922_),
    .B2(_09917_),
    .X(_09984_));
 sky130_fd_sc_hd__a211o_1 _18134_ (.A1(_09977_),
    .A2(net1778),
    .B1(_09984_),
    .C1(net962),
    .X(_09985_));
 sky130_fd_sc_hd__nor2_1 _18135_ (.A(_09971_),
    .B(_09899_),
    .Y(_09986_));
 sky130_fd_sc_hd__a21o_1 _18136_ (.A1(_09914_),
    .A2(_09923_),
    .B1(_09929_),
    .X(_09987_));
 sky130_fd_sc_hd__mux2_1 _18137_ (.A0(_09930_),
    .A1(_09987_),
    .S(_09901_),
    .X(_09988_));
 sky130_fd_sc_hd__nand2_1 _18138_ (.A(_09930_),
    .B(_09987_),
    .Y(_09989_));
 sky130_fd_sc_hd__inv_2 _18139_ (.A(_09945_),
    .Y(_09990_));
 sky130_fd_sc_hd__mux2_1 _18140_ (.A0(_09944_),
    .A1(_09990_),
    .S(_09901_),
    .X(_09991_));
 sky130_fd_sc_hd__o221a_1 _18141_ (.A1(_09939_),
    .A2(_09988_),
    .B1(_09989_),
    .B2(_09991_),
    .C1(net2548),
    .X(_09992_));
 sky130_fd_sc_hd__o22a_1 _18142_ (.A1(_09987_),
    .A2(_09944_),
    .B1(_09989_),
    .B2(_09939_),
    .X(_09993_));
 sky130_fd_sc_hd__a31o_1 _18143_ (.A1(_09901_),
    .A2(_09941_),
    .A3(_09945_),
    .B1(net2548),
    .X(_09994_));
 sky130_fd_sc_hd__o21ba_1 _18144_ (.A1(_09901_),
    .A2(_09993_),
    .B1_N(_09994_),
    .X(_09995_));
 sky130_fd_sc_hd__or4_1 _18145_ (.A(_09985_),
    .B(_09986_),
    .C(_09992_),
    .D(_09995_),
    .X(_09996_));
 sky130_fd_sc_hd__a211oi_1 _18146_ (.A1(_09872_),
    .A2(net2549),
    .B1(_09873_),
    .C1(_09958_),
    .Y(_09997_));
 sky130_fd_sc_hd__or2_1 _18147_ (.A(_09872_),
    .B(net2549),
    .X(_09998_));
 sky130_fd_sc_hd__and2_1 _18148_ (.A(_09998_),
    .B(_09957_),
    .X(_09999_));
 sky130_fd_sc_hd__nor2_1 _18149_ (.A(_09954_),
    .B(_09957_),
    .Y(_10000_));
 sky130_fd_sc_hd__o22a_1 _18150_ (.A1(_09951_),
    .A2(_09997_),
    .B1(_09999_),
    .B2(_10000_),
    .X(_10001_));
 sky130_fd_sc_hd__o21ba_1 _18151_ (.A1(_09998_),
    .A2(net3234),
    .B1_N(_09956_),
    .X(_10002_));
 sky130_fd_sc_hd__a21oi_1 _18152_ (.A1(_09998_),
    .A2(net3234),
    .B1(_10002_),
    .Y(_10003_));
 sky130_fd_sc_hd__xor2_1 _18153_ (.A(_09751_),
    .B(_09755_),
    .X(_10004_));
 sky130_fd_sc_hd__xor2_1 _18154_ (.A(_09758_),
    .B(_10004_),
    .X(_10005_));
 sky130_fd_sc_hd__or2_1 _18155_ (.A(_10003_),
    .B(_10005_),
    .X(_10006_));
 sky130_fd_sc_hd__a21o_1 _18156_ (.A1(_09960_),
    .A2(_09969_),
    .B1(_09968_),
    .X(_10007_));
 sky130_fd_sc_hd__a21o_1 _18157_ (.A1(_10003_),
    .A2(_10005_),
    .B1(net1212),
    .X(_10008_));
 sky130_fd_sc_hd__and3_1 _18158_ (.A(_10003_),
    .B(_10005_),
    .C(net1212),
    .X(_10009_));
 sky130_fd_sc_hd__nand2_1 _18159_ (.A(_09769_),
    .B(_09770_),
    .Y(_10010_));
 sky130_fd_sc_hd__xor2_1 _18160_ (.A(_09747_),
    .B(_09760_),
    .X(_10011_));
 sky130_fd_sc_hd__xnor2_1 _18161_ (.A(_10010_),
    .B(_10011_),
    .Y(_10012_));
 sky130_fd_sc_hd__a311oi_1 _18162_ (.A1(_10001_),
    .A2(_10006_),
    .A3(_10008_),
    .B1(_10009_),
    .C1(_10012_),
    .Y(_10013_));
 sky130_fd_sc_hd__xnor2_1 _18163_ (.A(net1212),
    .B(_10001_),
    .Y(_10014_));
 sky130_fd_sc_hd__or3b_1 _18164_ (.A(_10001_),
    .B(_10008_),
    .C_N(_10006_),
    .X(_10015_));
 sky130_fd_sc_hd__o211a_1 _18165_ (.A1(_10006_),
    .A2(_10014_),
    .B1(_10015_),
    .C1(_10012_),
    .X(_10016_));
 sky130_fd_sc_hd__a211o_1 _18166_ (.A1(net819),
    .A2(net818),
    .B1(_10013_),
    .C1(_10016_),
    .X(_10017_));
 sky130_fd_sc_hd__a21o_1 _18167_ (.A1(_10006_),
    .A2(_10008_),
    .B1(_10001_),
    .X(_10018_));
 sky130_fd_sc_hd__o211ai_1 _18168_ (.A1(net1212),
    .A2(_10006_),
    .B1(_10018_),
    .C1(_10012_),
    .Y(_10019_));
 sky130_fd_sc_hd__or2_1 _18169_ (.A(_09840_),
    .B(_09839_),
    .X(_10020_));
 sky130_fd_sc_hd__o31a_1 _18170_ (.A1(_09777_),
    .A2(_09778_),
    .A3(_09779_),
    .B1(_09673_),
    .X(_10021_));
 sky130_fd_sc_hd__a22o_1 _18171_ (.A1(_10020_),
    .A2(_09776_),
    .B1(_10021_),
    .B2(_09841_),
    .X(_10022_));
 sky130_fd_sc_hd__a31o_1 _18172_ (.A1(_09842_),
    .A2(net768),
    .A3(net817),
    .B1(_10022_),
    .X(_10023_));
 sky130_fd_sc_hd__o21ai_1 _18173_ (.A1(_09688_),
    .A2(_09780_),
    .B1(_09781_),
    .Y(_10024_));
 sky130_fd_sc_hd__o21a_1 _18174_ (.A1(_09686_),
    .A2(_09787_),
    .B1(_09784_),
    .X(_10025_));
 sky130_fd_sc_hd__nand2_1 _18175_ (.A(_10025_),
    .B(_09822_),
    .Y(_10026_));
 sky130_fd_sc_hd__or2_1 _18176_ (.A(_10025_),
    .B(_09822_),
    .X(_10027_));
 sky130_fd_sc_hd__o211a_1 _18177_ (.A1(_09817_),
    .A2(_10024_),
    .B1(_10026_),
    .C1(_10027_),
    .X(_10028_));
 sky130_fd_sc_hd__a21o_1 _18178_ (.A1(_09817_),
    .A2(_10024_),
    .B1(_10028_),
    .X(_10029_));
 sky130_fd_sc_hd__nand2_1 _18179_ (.A(net3340),
    .B(net7142),
    .Y(_10030_));
 sky130_fd_sc_hd__nor2_1 _18180_ (.A(net3340),
    .B(net7142),
    .Y(_10031_));
 sky130_fd_sc_hd__xnor2_1 _18181_ (.A(net3346),
    .B(_09630_),
    .Y(_10032_));
 sky130_fd_sc_hd__o21a_1 _18182_ (.A1(_10031_),
    .A2(_10032_),
    .B1(_10030_),
    .X(_10033_));
 sky130_fd_sc_hd__nand2_1 _18183_ (.A(net7063),
    .B(net3254),
    .Y(_10034_));
 sky130_fd_sc_hd__or3b_1 _18184_ (.A(net7142),
    .B(_10034_),
    .C_N(_09630_),
    .X(_10035_));
 sky130_fd_sc_hd__o221a_1 _18185_ (.A1(_10030_),
    .A2(_09630_),
    .B1(_10033_),
    .B2(net3254),
    .C1(_10035_),
    .X(_10036_));
 sky130_fd_sc_hd__xnor2_4 _18186_ (.A(net7032),
    .B(net7124),
    .Y(_10037_));
 sky130_fd_sc_hd__xnor2_4 _18187_ (.A(_10037_),
    .B(net2554),
    .Y(_10038_));
 sky130_fd_sc_hd__xnor2_2 _18188_ (.A(net6847),
    .B(net6875),
    .Y(_10039_));
 sky130_fd_sc_hd__and2b_2 _18189_ (.A_N(net6953),
    .B(net6922),
    .X(_10040_));
 sky130_fd_sc_hd__xnor2_4 _18190_ (.A(net6892),
    .B(_10040_),
    .Y(_10041_));
 sky130_fd_sc_hd__xnor2_1 _18191_ (.A(_10039_),
    .B(_10041_),
    .Y(_10042_));
 sky130_fd_sc_hd__nor2_1 _18192_ (.A(net6927),
    .B(net6945),
    .Y(_10043_));
 sky130_fd_sc_hd__o21bai_1 _18193_ (.A1(net3948),
    .A2(_09793_),
    .B1_N(_10043_),
    .Y(_10044_));
 sky130_fd_sc_hd__nand2_1 _18194_ (.A(net6920),
    .B(net6949),
    .Y(_10045_));
 sky130_fd_sc_hd__a21oi_1 _18195_ (.A1(_09793_),
    .A2(net3936),
    .B1(net6973),
    .Y(_10046_));
 sky130_fd_sc_hd__a21oi_1 _18196_ (.A1(_08984_),
    .A2(net3952),
    .B1(_09609_),
    .Y(_10047_));
 sky130_fd_sc_hd__o21ai_2 _18197_ (.A1(net3997),
    .A2(net3952),
    .B1(net6996),
    .Y(_10048_));
 sky130_fd_sc_hd__o211ai_1 _18198_ (.A1(_10044_),
    .A2(_10046_),
    .B1(net3233),
    .C1(_10048_),
    .Y(_10049_));
 sky130_fd_sc_hd__a211o_1 _18199_ (.A1(net3233),
    .A2(_10048_),
    .B1(_10044_),
    .C1(_10046_),
    .X(_10050_));
 sky130_fd_sc_hd__nand3_1 _18200_ (.A(net2547),
    .B(_10049_),
    .C(_10050_),
    .Y(_10051_));
 sky130_fd_sc_hd__a21o_1 _18201_ (.A1(_10049_),
    .A2(_10050_),
    .B1(net2547),
    .X(_10052_));
 sky130_fd_sc_hd__and2_1 _18202_ (.A(_10051_),
    .B(_10052_),
    .X(_10053_));
 sky130_fd_sc_hd__xnor2_1 _18203_ (.A(_10038_),
    .B(_10053_),
    .Y(_10054_));
 sky130_fd_sc_hd__xnor2_1 _18204_ (.A(_10036_),
    .B(_10054_),
    .Y(_10055_));
 sky130_fd_sc_hd__a31o_1 _18205_ (.A1(net2139),
    .A2(_09805_),
    .A3(_09806_),
    .B1(_09812_),
    .X(_10056_));
 sky130_fd_sc_hd__o21ai_1 _18206_ (.A1(net2139),
    .A2(_09807_),
    .B1(_10056_),
    .Y(_10057_));
 sky130_fd_sc_hd__o21ba_1 _18207_ (.A1(net3956),
    .A2(_09676_),
    .B1_N(_09796_),
    .X(_10058_));
 sky130_fd_sc_hd__a21o_1 _18208_ (.A1(_09798_),
    .A2(_09676_),
    .B1(net6997),
    .X(_10059_));
 sky130_fd_sc_hd__a22o_1 _18209_ (.A1(net3239),
    .A2(net3238),
    .B1(_10058_),
    .B2(_10059_),
    .X(_10060_));
 sky130_fd_sc_hd__and4_1 _18210_ (.A(net3239),
    .B(net3238),
    .C(_10058_),
    .D(_10059_),
    .X(_10061_));
 sky130_fd_sc_hd__a21o_1 _18211_ (.A1(net2552),
    .A2(_10060_),
    .B1(_10061_),
    .X(_10062_));
 sky130_fd_sc_hd__buf_1 _18212_ (.A(net3947),
    .X(_10063_));
 sky130_fd_sc_hd__nand2_1 _18213_ (.A(net6886),
    .B(net6810),
    .Y(_10064_));
 sky130_fd_sc_hd__nand2_1 _18214_ (.A(net6894),
    .B(net6856),
    .Y(_10065_));
 sky130_fd_sc_hd__xnor2_1 _18215_ (.A(_09176_),
    .B(_10065_),
    .Y(_10066_));
 sky130_fd_sc_hd__o21ai_1 _18216_ (.A1(net3232),
    .A2(_10064_),
    .B1(_10066_),
    .Y(_10067_));
 sky130_fd_sc_hd__nor3_1 _18217_ (.A(net3947),
    .B(_10066_),
    .C(_10064_),
    .Y(_10068_));
 sky130_fd_sc_hd__inv_2 _18218_ (.A(net2545),
    .Y(_10069_));
 sky130_fd_sc_hd__nand2_1 _18219_ (.A(net2546),
    .B(_10069_),
    .Y(_10070_));
 sky130_fd_sc_hd__xor2_1 _18220_ (.A(_10062_),
    .B(_10070_),
    .X(_10071_));
 sky130_fd_sc_hd__xnor2_1 _18221_ (.A(_10057_),
    .B(_10071_),
    .Y(_10072_));
 sky130_fd_sc_hd__xnor2_1 _18222_ (.A(_10055_),
    .B(_10072_),
    .Y(_10073_));
 sky130_fd_sc_hd__or2_1 _18223_ (.A(_10029_),
    .B(_10073_),
    .X(_10074_));
 sky130_fd_sc_hd__nand2_1 _18224_ (.A(_10029_),
    .B(_10073_),
    .Y(_10075_));
 sky130_fd_sc_hd__mux2_1 _18225_ (.A0(_09696_),
    .A1(_09604_),
    .S(_10038_),
    .X(_10076_));
 sky130_fd_sc_hd__inv_2 _18226_ (.A(_10038_),
    .Y(_10077_));
 sky130_fd_sc_hd__a21oi_1 _18227_ (.A1(net7094),
    .A2(_10077_),
    .B1(_09809_),
    .Y(_10078_));
 sky130_fd_sc_hd__nor2_1 _18228_ (.A(_10053_),
    .B(_10078_),
    .Y(_10079_));
 sky130_fd_sc_hd__or2b_1 _18229_ (.A(net7144),
    .B_N(_09809_),
    .X(_10080_));
 sky130_fd_sc_hd__mux2_1 _18230_ (.A0(net7063),
    .A1(_10034_),
    .S(_10038_),
    .X(_10081_));
 sky130_fd_sc_hd__a21oi_1 _18231_ (.A1(_10053_),
    .A2(_10080_),
    .B1(_10081_),
    .Y(_10082_));
 sky130_fd_sc_hd__a31o_1 _18232_ (.A1(_10038_),
    .A2(_10051_),
    .A3(_10052_),
    .B1(net7141),
    .X(_10083_));
 sky130_fd_sc_hd__nand2_1 _18233_ (.A(_10077_),
    .B(_09809_),
    .Y(_10084_));
 sky130_fd_sc_hd__a21boi_1 _18234_ (.A1(_10083_),
    .A2(_10084_),
    .B1_N(_09810_),
    .Y(_10085_));
 sky130_fd_sc_hd__a2111o_1 _18235_ (.A1(net7144),
    .A2(_10076_),
    .B1(_10079_),
    .C1(_10082_),
    .D1(_10085_),
    .X(_10086_));
 sky130_fd_sc_hd__o21ai_1 _18236_ (.A1(net7142),
    .A2(net2554),
    .B1(_10037_),
    .Y(_10087_));
 sky130_fd_sc_hd__a21oi_1 _18237_ (.A1(net7142),
    .A2(net2554),
    .B1(net7095),
    .Y(_10088_));
 sky130_fd_sc_hd__nand2_1 _18238_ (.A(_10037_),
    .B(net2564),
    .Y(_10089_));
 sky130_fd_sc_hd__a221o_1 _18239_ (.A1(_10087_),
    .A2(_10088_),
    .B1(_10089_),
    .B2(net7095),
    .C1(net3340),
    .X(_10090_));
 sky130_fd_sc_hd__a211o_1 _18240_ (.A1(_10037_),
    .A2(net2564),
    .B1(_10030_),
    .C1(net3254),
    .X(_10091_));
 sky130_fd_sc_hd__o31a_1 _18241_ (.A1(net7063),
    .A2(_10037_),
    .A3(net2564),
    .B1(_10091_),
    .X(_10092_));
 sky130_fd_sc_hd__nand2_1 _18242_ (.A(_10090_),
    .B(net1777),
    .Y(_10093_));
 sky130_fd_sc_hd__or2_1 _18243_ (.A(net6894),
    .B(net6922),
    .X(_10094_));
 sky130_fd_sc_hd__a21boi_1 _18244_ (.A1(net3956),
    .A2(_10039_),
    .B1_N(_10094_),
    .Y(_10095_));
 sky130_fd_sc_hd__o21ai_1 _18245_ (.A1(_10039_),
    .A2(_10040_),
    .B1(net6911),
    .Y(_10096_));
 sky130_fd_sc_hd__a21o_1 _18246_ (.A1(net7075),
    .A2(net7098),
    .B1(net7014),
    .X(_10097_));
 sky130_fd_sc_hd__and2_1 _18247_ (.A(net3973),
    .B(_10097_),
    .X(_10098_));
 sky130_fd_sc_hd__o31ai_1 _18248_ (.A1(net4044),
    .A2(_09648_),
    .A3(net3267),
    .B1(net6964),
    .Y(_10099_));
 sky130_fd_sc_hd__a22o_1 _18249_ (.A1(_10095_),
    .A2(_10096_),
    .B1(_10098_),
    .B2(net2544),
    .X(_10100_));
 sky130_fd_sc_hd__nand4_1 _18250_ (.A(_10095_),
    .B(_10096_),
    .C(_10098_),
    .D(net2544),
    .Y(_10101_));
 sky130_fd_sc_hd__xnor2_2 _18251_ (.A(net6857),
    .B(net6811),
    .Y(_10102_));
 sky130_fd_sc_hd__nor2b_1 _18252_ (.A(net6920),
    .B_N(net6893),
    .Y(_10103_));
 sky130_fd_sc_hd__xnor2_1 _18253_ (.A(net6872),
    .B(net3932),
    .Y(_10104_));
 sky130_fd_sc_hd__xor2_1 _18254_ (.A(_10102_),
    .B(_10104_),
    .X(_10105_));
 sky130_fd_sc_hd__a21o_1 _18255_ (.A1(_10100_),
    .A2(_10101_),
    .B1(_10105_),
    .X(_10106_));
 sky130_fd_sc_hd__nand3_1 _18256_ (.A(_10105_),
    .B(_10100_),
    .C(_10101_),
    .Y(_10107_));
 sky130_fd_sc_hd__xnor2_2 _18257_ (.A(net7012),
    .B(net7115),
    .Y(_10108_));
 sky130_fd_sc_hd__and3b_1 _18258_ (.A_N(net7032),
    .B(net7124),
    .C(net7064),
    .X(_10109_));
 sky130_fd_sc_hd__a21oi_1 _18259_ (.A1(net3996),
    .A2(net3972),
    .B1(_10109_),
    .Y(_10110_));
 sky130_fd_sc_hd__xnor2_1 _18260_ (.A(_10108_),
    .B(_10110_),
    .Y(_10111_));
 sky130_fd_sc_hd__xnor2_1 _18261_ (.A(net3247),
    .B(_10111_),
    .Y(_10112_));
 sky130_fd_sc_hd__nand3_1 _18262_ (.A(_10106_),
    .B(_10107_),
    .C(net2138),
    .Y(_10113_));
 sky130_fd_sc_hd__a21o_1 _18263_ (.A1(_10106_),
    .A2(_10107_),
    .B1(net2138),
    .X(_10114_));
 sky130_fd_sc_hd__nand3_1 _18264_ (.A(_10093_),
    .B(_10113_),
    .C(_10114_),
    .Y(_10115_));
 sky130_fd_sc_hd__a21o_1 _18265_ (.A1(_10113_),
    .A2(_10114_),
    .B1(_10093_),
    .X(_10116_));
 sky130_fd_sc_hd__nand2_1 _18266_ (.A(net3233),
    .B(_10048_),
    .Y(_10117_));
 sky130_fd_sc_hd__or2_1 _18267_ (.A(_10044_),
    .B(_10046_),
    .X(_10118_));
 sky130_fd_sc_hd__o21a_1 _18268_ (.A1(_10117_),
    .A2(_10118_),
    .B1(net2547),
    .X(_10119_));
 sky130_fd_sc_hd__a21oi_1 _18269_ (.A1(_10117_),
    .A2(_10118_),
    .B1(_10119_),
    .Y(_10120_));
 sky130_fd_sc_hd__nor2_1 _18270_ (.A(_09176_),
    .B(_10065_),
    .Y(_10121_));
 sky130_fd_sc_hd__inv_2 _18271_ (.A(net6760),
    .Y(_10122_));
 sky130_fd_sc_hd__nand2_1 _18272_ (.A(net6832),
    .B(net6881),
    .Y(_10123_));
 sky130_fd_sc_hd__xnor2_1 _18273_ (.A(net3928),
    .B(net3926),
    .Y(_10124_));
 sky130_fd_sc_hd__xnor2_1 _18274_ (.A(_10121_),
    .B(net3228),
    .Y(_10125_));
 sky130_fd_sc_hd__xnor2_1 _18275_ (.A(net1776),
    .B(_10125_),
    .Y(_10126_));
 sky130_fd_sc_hd__nand3_1 _18276_ (.A(_10115_),
    .B(_10116_),
    .C(_10126_),
    .Y(_10127_));
 sky130_fd_sc_hd__a21o_1 _18277_ (.A1(_10115_),
    .A2(_10116_),
    .B1(_10126_),
    .X(_10128_));
 sky130_fd_sc_hd__and3_1 _18278_ (.A(net1074),
    .B(_10127_),
    .C(_10128_),
    .X(_10129_));
 sky130_fd_sc_hd__a21oi_1 _18279_ (.A1(_10127_),
    .A2(_10128_),
    .B1(net1074),
    .Y(_10130_));
 sky130_fd_sc_hd__nor2_1 _18280_ (.A(_10129_),
    .B(_10130_),
    .Y(_10131_));
 sky130_fd_sc_hd__a21oi_1 _18281_ (.A1(net2546),
    .A2(_10062_),
    .B1(net2545),
    .Y(_10132_));
 sky130_fd_sc_hd__or2_1 _18282_ (.A(_10057_),
    .B(_10071_),
    .X(_10133_));
 sky130_fd_sc_hd__and2_1 _18283_ (.A(_10057_),
    .B(_10071_),
    .X(_10134_));
 sky130_fd_sc_hd__a21oi_1 _18284_ (.A1(_10133_),
    .A2(_10055_),
    .B1(_10134_),
    .Y(_10135_));
 sky130_fd_sc_hd__xnor2_1 _18285_ (.A(_10132_),
    .B(_10135_),
    .Y(_10136_));
 sky130_fd_sc_hd__xnor2_1 _18286_ (.A(_10131_),
    .B(_10136_),
    .Y(_10137_));
 sky130_fd_sc_hd__mux2_1 _18287_ (.A0(_10074_),
    .A1(_10075_),
    .S(_10137_),
    .X(_10138_));
 sky130_fd_sc_hd__nand2_1 _18288_ (.A(net963),
    .B(_09834_),
    .Y(_10139_));
 sky130_fd_sc_hd__a21o_1 _18289_ (.A1(net3245),
    .A2(net1215),
    .B1(net1447),
    .X(_10140_));
 sky130_fd_sc_hd__o21ai_1 _18290_ (.A1(net3245),
    .A2(net1215),
    .B1(_10140_),
    .Y(_10141_));
 sky130_fd_sc_hd__o21ai_1 _18291_ (.A1(net963),
    .A2(_09834_),
    .B1(_10141_),
    .Y(_10142_));
 sky130_fd_sc_hd__and3b_1 _18292_ (.A_N(net963),
    .B(_09835_),
    .C(_09829_),
    .X(_10143_));
 sky130_fd_sc_hd__nand2_1 _18293_ (.A(net1215),
    .B(net1447),
    .Y(_10144_));
 sky130_fd_sc_hd__a21oi_1 _18294_ (.A1(net963),
    .A2(_10144_),
    .B1(_09836_),
    .Y(_10145_));
 sky130_fd_sc_hd__a211o_1 _18295_ (.A1(_10139_),
    .A2(_10142_),
    .B1(_10143_),
    .C1(_10145_),
    .X(_10146_));
 sky130_fd_sc_hd__a21oi_2 _18296_ (.A1(_10025_),
    .A2(_09821_),
    .B1(_09820_),
    .Y(_10147_));
 sky130_fd_sc_hd__xnor2_1 _18297_ (.A(net815),
    .B(_10147_),
    .Y(_10148_));
 sky130_fd_sc_hd__and2_1 _18298_ (.A(_10075_),
    .B(_10074_),
    .X(_10149_));
 sky130_fd_sc_hd__or4b_1 _18299_ (.A(net815),
    .B(_10147_),
    .C(_10137_),
    .D_N(_10149_),
    .X(_10150_));
 sky130_fd_sc_hd__nand4_1 _18300_ (.A(net815),
    .B(_10147_),
    .C(_10137_),
    .D(_10149_),
    .Y(_10151_));
 sky130_fd_sc_hd__o211a_1 _18301_ (.A1(_10138_),
    .A2(_10148_),
    .B1(_10150_),
    .C1(_10151_),
    .X(_10152_));
 sky130_fd_sc_hd__a21boi_1 _18302_ (.A1(_10105_),
    .A2(_10100_),
    .B1_N(_10101_),
    .Y(_10153_));
 sky130_fd_sc_hd__nand2_1 _18303_ (.A(net6774),
    .B(net3926),
    .Y(_10154_));
 sky130_fd_sc_hd__nand2_1 _18304_ (.A(net6857),
    .B(net6811),
    .Y(_10155_));
 sky130_fd_sc_hd__xnor2_1 _18305_ (.A(_10154_),
    .B(_10155_),
    .Y(_10156_));
 sky130_fd_sc_hd__xnor2_2 _18306_ (.A(net1775),
    .B(_10156_),
    .Y(_10157_));
 sky130_fd_sc_hd__mux2_1 _18307_ (.A0(_09675_),
    .A1(net3331),
    .S(_10108_),
    .X(_10158_));
 sky130_fd_sc_hd__a211o_1 _18308_ (.A1(_09675_),
    .A2(_10108_),
    .B1(_08967_),
    .C1(net7040),
    .X(_10159_));
 sky130_fd_sc_hd__o21ai_1 _18309_ (.A1(net7071),
    .A2(_10158_),
    .B1(_10159_),
    .Y(_10160_));
 sky130_fd_sc_hd__xnor2_1 _18310_ (.A(net7072),
    .B(_09675_),
    .Y(_10161_));
 sky130_fd_sc_hd__nor3_1 _18311_ (.A(net7046),
    .B(_09675_),
    .C(_10108_),
    .Y(_10162_));
 sky130_fd_sc_hd__a31o_1 _18312_ (.A1(net7040),
    .A2(_10161_),
    .A3(_10108_),
    .B1(_10162_),
    .X(_10163_));
 sky130_fd_sc_hd__a21o_1 _18313_ (.A1(net7126),
    .A2(_10160_),
    .B1(_10163_),
    .X(_10164_));
 sky130_fd_sc_hd__and3_1 _18314_ (.A(_09026_),
    .B(net7034),
    .C(net7110),
    .X(_10165_));
 sky130_fd_sc_hd__a21oi_1 _18315_ (.A1(net3347),
    .A2(_09606_),
    .B1(net3226),
    .Y(_10166_));
 sky130_fd_sc_hd__xnor2_1 _18316_ (.A(net3241),
    .B(_09909_),
    .Y(_10167_));
 sky130_fd_sc_hd__xnor2_1 _18317_ (.A(_10166_),
    .B(_10167_),
    .Y(_10168_));
 sky130_fd_sc_hd__xnor2_2 _18318_ (.A(net6842),
    .B(net6789),
    .Y(_10169_));
 sky130_fd_sc_hd__and2b_1 _18319_ (.A_N(net6903),
    .B(net6887),
    .X(_10170_));
 sky130_fd_sc_hd__xnor2_4 _18320_ (.A(net6852),
    .B(_10170_),
    .Y(_10171_));
 sky130_fd_sc_hd__xor2_2 _18321_ (.A(_10169_),
    .B(_10171_),
    .X(_10172_));
 sky130_fd_sc_hd__a21o_1 _18322_ (.A1(net6892),
    .A2(net6872),
    .B1(_10102_),
    .X(_10173_));
 sky130_fd_sc_hd__nor2_1 _18323_ (.A(net6892),
    .B(net6872),
    .Y(_10174_));
 sky130_fd_sc_hd__a221o_1 _18324_ (.A1(net6872),
    .A2(_10102_),
    .B1(_10173_),
    .B2(net3947),
    .C1(_10174_),
    .X(_10175_));
 sky130_fd_sc_hd__or2b_1 _18325_ (.A(_09680_),
    .B_N(net3955),
    .X(_10176_));
 sky130_fd_sc_hd__a221o_1 _18326_ (.A1(net6945),
    .A2(_09680_),
    .B1(_10176_),
    .B2(net3986),
    .C1(_09796_),
    .X(_10177_));
 sky130_fd_sc_hd__xnor2_1 _18327_ (.A(_10175_),
    .B(net2543),
    .Y(_10178_));
 sky130_fd_sc_hd__xnor2_2 _18328_ (.A(_10172_),
    .B(_10178_),
    .Y(_10179_));
 sky130_fd_sc_hd__xnor2_1 _18329_ (.A(_10168_),
    .B(_10179_),
    .Y(_10180_));
 sky130_fd_sc_hd__xor2_1 _18330_ (.A(_10164_),
    .B(_10180_),
    .X(_10181_));
 sky130_fd_sc_hd__or2b_1 _18331_ (.A(_10093_),
    .B_N(net2138),
    .X(_10182_));
 sky130_fd_sc_hd__a21oi_1 _18332_ (.A1(_10090_),
    .A2(net1777),
    .B1(net2138),
    .Y(_10183_));
 sky130_fd_sc_hd__a31oi_1 _18333_ (.A1(_10106_),
    .A2(_10107_),
    .A3(_10182_),
    .B1(_10183_),
    .Y(_10184_));
 sky130_fd_sc_hd__xnor2_1 _18334_ (.A(net1211),
    .B(net1073),
    .Y(_10185_));
 sky130_fd_sc_hd__xnor2_2 _18335_ (.A(_10157_),
    .B(_10185_),
    .Y(_10186_));
 sky130_fd_sc_hd__nor2_1 _18336_ (.A(_10121_),
    .B(net1776),
    .Y(_10187_));
 sky130_fd_sc_hd__nand2_1 _18337_ (.A(_10121_),
    .B(net1776),
    .Y(_10188_));
 sky130_fd_sc_hd__o21ai_2 _18338_ (.A1(net3228),
    .A2(_10187_),
    .B1(_10188_),
    .Y(_10189_));
 sky130_fd_sc_hd__a21boi_1 _18339_ (.A1(net1074),
    .A2(_10128_),
    .B1_N(_10127_),
    .Y(_10190_));
 sky130_fd_sc_hd__xor2_1 _18340_ (.A(_10189_),
    .B(_10190_),
    .X(_10191_));
 sky130_fd_sc_hd__xnor2_2 _18341_ (.A(_10186_),
    .B(_10191_),
    .Y(_10192_));
 sky130_fd_sc_hd__and2b_1 _18342_ (.A_N(_10135_),
    .B(_10132_),
    .X(_10193_));
 sky130_fd_sc_hd__or2b_1 _18343_ (.A(_10132_),
    .B_N(_10135_),
    .X(_10194_));
 sky130_fd_sc_hd__o21a_1 _18344_ (.A1(_10193_),
    .A2(_10131_),
    .B1(_10194_),
    .X(_10195_));
 sky130_fd_sc_hd__and2_1 _18345_ (.A(_10192_),
    .B(_10195_),
    .X(_10196_));
 sky130_fd_sc_hd__o21a_1 _18346_ (.A1(_10192_),
    .A2(_10193_),
    .B1(_10131_),
    .X(_10197_));
 sky130_fd_sc_hd__a21o_1 _18347_ (.A1(_10192_),
    .A2(_10194_),
    .B1(_10197_),
    .X(_10198_));
 sky130_fd_sc_hd__inv_2 _18348_ (.A(_10075_),
    .Y(_10199_));
 sky130_fd_sc_hd__a21bo_1 _18349_ (.A1(_10147_),
    .A2(_10074_),
    .B1_N(_10075_),
    .X(_10200_));
 sky130_fd_sc_hd__a22o_1 _18350_ (.A1(_10147_),
    .A2(_10199_),
    .B1(_10200_),
    .B2(net815),
    .X(_10201_));
 sky130_fd_sc_hd__o21a_1 _18351_ (.A1(_10192_),
    .A2(_10195_),
    .B1(_10201_),
    .X(_10202_));
 sky130_fd_sc_hd__o32a_1 _18352_ (.A1(net716),
    .A2(net715),
    .A3(_10196_),
    .B1(_10198_),
    .B2(_10202_),
    .X(_10203_));
 sky130_fd_sc_hd__a21o_1 _18353_ (.A1(_10186_),
    .A2(_10189_),
    .B1(_10190_),
    .X(_10204_));
 sky130_fd_sc_hd__o21a_1 _18354_ (.A1(_10186_),
    .A2(_10189_),
    .B1(_10204_),
    .X(_10205_));
 sky130_fd_sc_hd__nand2_1 _18355_ (.A(net6773),
    .B(_10155_),
    .Y(_10206_));
 sky130_fd_sc_hd__inv_2 _18356_ (.A(_10171_),
    .Y(_10207_));
 sky130_fd_sc_hd__nor2_1 _18357_ (.A(_10175_),
    .B(net2543),
    .Y(_10208_));
 sky130_fd_sc_hd__nand2_1 _18358_ (.A(_10175_),
    .B(net2543),
    .Y(_10209_));
 sky130_fd_sc_hd__o21ai_1 _18359_ (.A1(_10207_),
    .A2(_10208_),
    .B1(_10209_),
    .Y(_10210_));
 sky130_fd_sc_hd__nand2_1 _18360_ (.A(net6842),
    .B(net6789),
    .Y(_10211_));
 sky130_fd_sc_hd__xnor2_1 _18361_ (.A(net6789),
    .B(_10171_),
    .Y(_10212_));
 sky130_fd_sc_hd__nor2_1 _18362_ (.A(net6789),
    .B(_10207_),
    .Y(_10213_));
 sky130_fd_sc_hd__mux2_1 _18363_ (.A0(_10212_),
    .A1(_10213_),
    .S(net6842),
    .X(_10214_));
 sky130_fd_sc_hd__a22o_1 _18364_ (.A1(_10208_),
    .A2(_10211_),
    .B1(_10214_),
    .B2(_10209_),
    .X(_10215_));
 sky130_fd_sc_hd__a31o_1 _18365_ (.A1(net6825),
    .A2(net6798),
    .A3(_10210_),
    .B1(_10215_),
    .X(_10216_));
 sky130_fd_sc_hd__xnor2_2 _18366_ (.A(_10206_),
    .B(_10216_),
    .Y(_10217_));
 sky130_fd_sc_hd__and2_1 _18367_ (.A(net6863),
    .B(net6876),
    .X(_10218_));
 sky130_fd_sc_hd__or2_1 _18368_ (.A(_10169_),
    .B(net3924),
    .X(_10219_));
 sky130_fd_sc_hd__nor2_1 _18369_ (.A(net6858),
    .B(net6879),
    .Y(_10220_));
 sky130_fd_sc_hd__a221o_1 _18370_ (.A1(net6858),
    .A2(_10169_),
    .B1(_10219_),
    .B2(net3299),
    .C1(_10220_),
    .X(_10221_));
 sky130_fd_sc_hd__and2b_1 _18371_ (.A_N(net6882),
    .B(net6854),
    .X(_10222_));
 sky130_fd_sc_hd__xnor2_2 _18372_ (.A(net6825),
    .B(_10222_),
    .Y(_10223_));
 sky130_fd_sc_hd__xnor2_2 _18373_ (.A(net6807),
    .B(net6774),
    .Y(_10224_));
 sky130_fd_sc_hd__xor2_1 _18374_ (.A(_10223_),
    .B(_10224_),
    .X(_10225_));
 sky130_fd_sc_hd__nand2_1 _18375_ (.A(net7015),
    .B(net7046),
    .Y(_10226_));
 sky130_fd_sc_hd__nand2_1 _18376_ (.A(net3936),
    .B(_09634_),
    .Y(_10227_));
 sky130_fd_sc_hd__a221o_1 _18377_ (.A1(net6927),
    .A2(_10226_),
    .B1(_10227_),
    .B2(net3311),
    .C1(_10043_),
    .X(_10228_));
 sky130_fd_sc_hd__xnor2_1 _18378_ (.A(_10225_),
    .B(net2541),
    .Y(_10229_));
 sky130_fd_sc_hd__xnor2_1 _18379_ (.A(_10221_),
    .B(_10229_),
    .Y(_10230_));
 sky130_fd_sc_hd__mux2_1 _18380_ (.A0(net7043),
    .A1(_09704_),
    .S(net3241),
    .X(_10231_));
 sky130_fd_sc_hd__nand2_1 _18381_ (.A(net7012),
    .B(_09909_),
    .Y(_10232_));
 sky130_fd_sc_hd__nand2_1 _18382_ (.A(net7045),
    .B(net7111),
    .Y(_10233_));
 sky130_fd_sc_hd__a21o_1 _18383_ (.A1(net3241),
    .A2(_10233_),
    .B1(_09909_),
    .X(_10234_));
 sky130_fd_sc_hd__or2_1 _18384_ (.A(net3241),
    .B(_10233_),
    .X(_10235_));
 sky130_fd_sc_hd__a21o_1 _18385_ (.A1(_10234_),
    .A2(_10235_),
    .B1(net7012),
    .X(_10236_));
 sky130_fd_sc_hd__or3b_1 _18386_ (.A(net3241),
    .B(_09909_),
    .C_N(_09701_),
    .X(_10237_));
 sky130_fd_sc_hd__o211ai_1 _18387_ (.A1(_10231_),
    .A2(_10232_),
    .B1(_10236_),
    .C1(_10237_),
    .Y(_10238_));
 sky130_fd_sc_hd__and3_1 _18388_ (.A(net3986),
    .B(net7014),
    .C(net7098),
    .X(_10239_));
 sky130_fd_sc_hd__a21oi_1 _18389_ (.A1(net3253),
    .A2(net3267),
    .B1(_10239_),
    .Y(_10240_));
 sky130_fd_sc_hd__xnor2_2 _18390_ (.A(net6979),
    .B(net7071),
    .Y(_10241_));
 sky130_fd_sc_hd__xnor2_1 _18391_ (.A(_10041_),
    .B(_10241_),
    .Y(_10242_));
 sky130_fd_sc_hd__xnor2_1 _18392_ (.A(_10240_),
    .B(_10242_),
    .Y(_10243_));
 sky130_fd_sc_hd__xnor2_1 _18393_ (.A(net1773),
    .B(_10243_),
    .Y(_10244_));
 sky130_fd_sc_hd__xnor2_1 _18394_ (.A(net1774),
    .B(_10244_),
    .Y(_10245_));
 sky130_fd_sc_hd__a21bo_1 _18395_ (.A1(_10164_),
    .A2(_10179_),
    .B1_N(_10168_),
    .X(_10246_));
 sky130_fd_sc_hd__o21a_1 _18396_ (.A1(_10164_),
    .A2(_10179_),
    .B1(_10246_),
    .X(_10247_));
 sky130_fd_sc_hd__xor2_1 _18397_ (.A(_10245_),
    .B(net1210),
    .X(_10248_));
 sky130_fd_sc_hd__xnor2_2 _18398_ (.A(_10217_),
    .B(_10248_),
    .Y(_10249_));
 sky130_fd_sc_hd__a31o_1 _18399_ (.A1(net6854),
    .A2(net6811),
    .A3(net6774),
    .B1(net1775),
    .X(_10250_));
 sky130_fd_sc_hd__or2_1 _18400_ (.A(_10155_),
    .B(net1775),
    .X(_10251_));
 sky130_fd_sc_hd__a22o_1 _18401_ (.A1(net3926),
    .A2(_10250_),
    .B1(_10206_),
    .B2(_10251_),
    .X(_10252_));
 sky130_fd_sc_hd__o21ba_1 _18402_ (.A1(net1073),
    .A2(_10157_),
    .B1_N(net1211),
    .X(_10253_));
 sky130_fd_sc_hd__a21oi_2 _18403_ (.A1(net1073),
    .A2(_10157_),
    .B1(_10253_),
    .Y(_10254_));
 sky130_fd_sc_hd__xnor2_1 _18404_ (.A(_10252_),
    .B(_10254_),
    .Y(_10255_));
 sky130_fd_sc_hd__xnor2_1 _18405_ (.A(_10249_),
    .B(_10255_),
    .Y(_10256_));
 sky130_fd_sc_hd__and2b_1 _18406_ (.A_N(_10205_),
    .B(net767),
    .X(_10257_));
 sky130_fd_sc_hd__or2b_1 _18407_ (.A(net767),
    .B_N(_10205_),
    .X(_10258_));
 sky130_fd_sc_hd__and2b_1 _18408_ (.A_N(_10257_),
    .B(_10258_),
    .X(_10259_));
 sky130_fd_sc_hd__xor2_1 _18409_ (.A(_10203_),
    .B(_10259_),
    .X(_10260_));
 sky130_fd_sc_hd__buf_1 _18410_ (.A(net1786),
    .X(_10261_));
 sky130_fd_sc_hd__nor2_1 _18411_ (.A(net606),
    .B(_10261_),
    .Y(_10262_));
 sky130_fd_sc_hd__a31o_1 _18412_ (.A1(net9059),
    .A2(net2289),
    .A3(_09598_),
    .B1(_10262_),
    .X(_00439_));
 sky130_fd_sc_hd__nor2_1 _18413_ (.A(net4245),
    .B(net2932),
    .Y(_10263_));
 sky130_fd_sc_hd__clkbuf_1 _18414_ (.A(net2135),
    .X(_10264_));
 sky130_fd_sc_hd__xnor2_1 _18415_ (.A(_10192_),
    .B(_10195_),
    .Y(_10265_));
 sky130_fd_sc_hd__or4_1 _18416_ (.A(net716),
    .B(net715),
    .C(_10257_),
    .D(_10265_),
    .X(_10266_));
 sky130_fd_sc_hd__o31a_1 _18417_ (.A1(_10202_),
    .A2(_10198_),
    .A3(_10257_),
    .B1(_10258_),
    .X(_10267_));
 sky130_fd_sc_hd__o21ba_1 _18418_ (.A1(_10217_),
    .A2(net1210),
    .B1_N(_10245_),
    .X(_10268_));
 sky130_fd_sc_hd__a21oi_1 _18419_ (.A1(_10217_),
    .A2(net1210),
    .B1(_10268_),
    .Y(_10269_));
 sky130_fd_sc_hd__o21ai_1 _18420_ (.A1(_10172_),
    .A2(_10208_),
    .B1(_10209_),
    .Y(_10270_));
 sky130_fd_sc_hd__a31o_1 _18421_ (.A1(net6825),
    .A2(net6773),
    .A3(net6798),
    .B1(_10270_),
    .X(_10271_));
 sky130_fd_sc_hd__nand2_1 _18422_ (.A(_10155_),
    .B(_10271_),
    .Y(_10272_));
 sky130_fd_sc_hd__nand2_1 _18423_ (.A(net6773),
    .B(_10211_),
    .Y(_10273_));
 sky130_fd_sc_hd__o21ai_1 _18424_ (.A1(_10211_),
    .A2(_10270_),
    .B1(_10273_),
    .Y(_10274_));
 sky130_fd_sc_hd__and2_1 _18425_ (.A(net6826),
    .B(net3983),
    .X(_10275_));
 sky130_fd_sc_hd__clkbuf_2 _18426_ (.A(_10275_),
    .X(_10276_));
 sky130_fd_sc_hd__xnor2_1 _18427_ (.A(net6809),
    .B(_10276_),
    .Y(_10277_));
 sky130_fd_sc_hd__nor2_1 _18428_ (.A(net3929),
    .B(net6801),
    .Y(_10278_));
 sky130_fd_sc_hd__nor2_1 _18429_ (.A(net6785),
    .B(net3283),
    .Y(_10279_));
 sky130_fd_sc_hd__nor2_1 _18430_ (.A(_10278_),
    .B(_10279_),
    .Y(_10280_));
 sky130_fd_sc_hd__xnor2_1 _18431_ (.A(_10277_),
    .B(_10280_),
    .Y(_10281_));
 sky130_fd_sc_hd__nand2_1 _18432_ (.A(net3966),
    .B(_10224_),
    .Y(_10282_));
 sky130_fd_sc_hd__o21ai_1 _18433_ (.A1(_10222_),
    .A2(_10224_),
    .B1(net6827),
    .Y(_10283_));
 sky130_fd_sc_hd__o211a_1 _18434_ (.A1(net6836),
    .A2(net6859),
    .B1(_10282_),
    .C1(_10283_),
    .X(_10284_));
 sky130_fd_sc_hd__nand2_1 _18435_ (.A(net6897),
    .B(net6921),
    .Y(_10285_));
 sky130_fd_sc_hd__a22o_1 _18436_ (.A1(net7000),
    .A2(net7016),
    .B1(net3297),
    .B2(net6956),
    .X(_10286_));
 sky130_fd_sc_hd__o211a_1 _18437_ (.A1(net6956),
    .A2(_10285_),
    .B1(_10286_),
    .C1(net3933),
    .X(_10287_));
 sky130_fd_sc_hd__nor2_1 _18438_ (.A(_10284_),
    .B(_10287_),
    .Y(_10288_));
 sky130_fd_sc_hd__and2_1 _18439_ (.A(_10284_),
    .B(_10287_),
    .X(_10289_));
 sky130_fd_sc_hd__or2_1 _18440_ (.A(_10288_),
    .B(_10289_),
    .X(_10290_));
 sky130_fd_sc_hd__xnor2_1 _18441_ (.A(_10281_),
    .B(_10290_),
    .Y(_10291_));
 sky130_fd_sc_hd__nand2_1 _18442_ (.A(net7014),
    .B(net7099),
    .Y(_10292_));
 sky130_fd_sc_hd__a21o_1 _18443_ (.A1(_10041_),
    .A2(_10292_),
    .B1(_10241_),
    .X(_10293_));
 sky130_fd_sc_hd__o21a_1 _18444_ (.A1(_10041_),
    .A2(_10292_),
    .B1(_10293_),
    .X(_10294_));
 sky130_fd_sc_hd__nor2_1 _18445_ (.A(net7017),
    .B(net7099),
    .Y(_10295_));
 sky130_fd_sc_hd__mux2_1 _18446_ (.A0(net7014),
    .A1(_10295_),
    .S(_10041_),
    .X(_10296_));
 sky130_fd_sc_hd__nand2_1 _18447_ (.A(net6998),
    .B(_10241_),
    .Y(_10297_));
 sky130_fd_sc_hd__or4_1 _18448_ (.A(net7014),
    .B(net3253),
    .C(_10041_),
    .D(_10241_),
    .X(_10298_));
 sky130_fd_sc_hd__o221a_1 _18449_ (.A1(net6998),
    .A2(_10294_),
    .B1(_10296_),
    .B2(_10297_),
    .C1(_10298_),
    .X(_10299_));
 sky130_fd_sc_hd__or2_1 _18450_ (.A(net6988),
    .B(net7076),
    .X(_10300_));
 sky130_fd_sc_hd__mux2_1 _18451_ (.A0(net3941),
    .A1(_10300_),
    .S(net6970),
    .X(_10301_));
 sky130_fd_sc_hd__nor2_1 _18452_ (.A(net3961),
    .B(net7045),
    .Y(_10302_));
 sky130_fd_sc_hd__nor2_1 _18453_ (.A(net6933),
    .B(net3331),
    .Y(_10303_));
 sky130_fd_sc_hd__nor2_2 _18454_ (.A(_10302_),
    .B(_10303_),
    .Y(_10304_));
 sky130_fd_sc_hd__xnor2_1 _18455_ (.A(_10301_),
    .B(_10304_),
    .Y(_10305_));
 sky130_fd_sc_hd__xnor2_1 _18456_ (.A(net3229),
    .B(_10305_),
    .Y(_10306_));
 sky130_fd_sc_hd__xnor2_1 _18457_ (.A(net1766),
    .B(net1440),
    .Y(_10307_));
 sky130_fd_sc_hd__xnor2_1 _18458_ (.A(net1207),
    .B(_10307_),
    .Y(_10308_));
 sky130_fd_sc_hd__nand2_1 _18459_ (.A(_10221_),
    .B(net2541),
    .Y(_10309_));
 sky130_fd_sc_hd__nor2_1 _18460_ (.A(net3925),
    .B(net3225),
    .Y(_10310_));
 sky130_fd_sc_hd__and2_1 _18461_ (.A(net3925),
    .B(net3225),
    .X(_10311_));
 sky130_fd_sc_hd__mux2_1 _18462_ (.A0(_10310_),
    .A1(_10311_),
    .S(net3284),
    .X(_10312_));
 sky130_fd_sc_hd__mux2_1 _18463_ (.A0(_10310_),
    .A1(_10311_),
    .S(net6815),
    .X(_10313_));
 sky130_fd_sc_hd__xnor2_1 _18464_ (.A(net3284),
    .B(net3925),
    .Y(_10314_));
 sky130_fd_sc_hd__nor2_1 _18465_ (.A(_10221_),
    .B(net2541),
    .Y(_10315_));
 sky130_fd_sc_hd__mux2_1 _18466_ (.A0(_10313_),
    .A1(_10314_),
    .S(_10315_),
    .X(_10316_));
 sky130_fd_sc_hd__a21oi_1 _18467_ (.A1(_10309_),
    .A2(_10312_),
    .B1(_10316_),
    .Y(_10317_));
 sky130_fd_sc_hd__or2_1 _18468_ (.A(net3284),
    .B(net3225),
    .X(_10318_));
 sky130_fd_sc_hd__nand2_1 _18469_ (.A(net3284),
    .B(net3225),
    .Y(_10319_));
 sky130_fd_sc_hd__a311o_1 _18470_ (.A1(_10309_),
    .A2(_10318_),
    .A3(_10319_),
    .B1(_10315_),
    .C1(net6771),
    .X(_10320_));
 sky130_fd_sc_hd__or2_1 _18471_ (.A(_10309_),
    .B(_10314_),
    .X(_10321_));
 sky130_fd_sc_hd__o211a_1 _18472_ (.A1(net3930),
    .A2(_10317_),
    .B1(_10320_),
    .C1(_10321_),
    .X(_10322_));
 sky130_fd_sc_hd__or2b_1 _18473_ (.A(net1773),
    .B_N(_10243_),
    .X(_10323_));
 sky130_fd_sc_hd__and2b_1 _18474_ (.A_N(_10243_),
    .B(net1773),
    .X(_10324_));
 sky130_fd_sc_hd__a21o_1 _18475_ (.A1(net1774),
    .A2(_10323_),
    .B1(_10324_),
    .X(_10325_));
 sky130_fd_sc_hd__xor2_1 _18476_ (.A(_10322_),
    .B(net1205),
    .X(_10326_));
 sky130_fd_sc_hd__xnor2_1 _18477_ (.A(_10308_),
    .B(_10326_),
    .Y(_10327_));
 sky130_fd_sc_hd__nand3_1 _18478_ (.A(net1208),
    .B(net1441),
    .C(_10327_),
    .Y(_10328_));
 sky130_fd_sc_hd__a21o_1 _18479_ (.A1(net1208),
    .A2(net1441),
    .B1(_10327_),
    .X(_10329_));
 sky130_fd_sc_hd__nand2_1 _18480_ (.A(_10328_),
    .B(_10329_),
    .Y(_10330_));
 sky130_fd_sc_hd__xnor2_2 _18481_ (.A(net874),
    .B(_10330_),
    .Y(_10331_));
 sky130_fd_sc_hd__a21oi_2 _18482_ (.A1(net663),
    .A2(net659),
    .B1(_10331_),
    .Y(_10332_));
 sky130_fd_sc_hd__and3_1 _18483_ (.A(_10331_),
    .B(net663),
    .C(net659),
    .X(_10333_));
 sky130_fd_sc_hd__nor2_1 _18484_ (.A(_10332_),
    .B(_10333_),
    .Y(_10334_));
 sky130_fd_sc_hd__inv_2 _18485_ (.A(net6378),
    .Y(_10335_));
 sky130_fd_sc_hd__nor2_1 _18486_ (.A(net3923),
    .B(net607),
    .Y(_10336_));
 sky130_fd_sc_hd__a21bo_1 _18487_ (.A1(_10249_),
    .A2(_10254_),
    .B1_N(_10252_),
    .X(_10337_));
 sky130_fd_sc_hd__o21ai_1 _18488_ (.A1(_10249_),
    .A2(_10254_),
    .B1(_10337_),
    .Y(_10338_));
 sky130_fd_sc_hd__inv_2 _18489_ (.A(net765),
    .Y(_10339_));
 sky130_fd_sc_hd__xnor2_1 _18490_ (.A(_10336_),
    .B(_10339_),
    .Y(_10340_));
 sky130_fd_sc_hd__xnor2_1 _18491_ (.A(_10334_),
    .B(_10340_),
    .Y(_10341_));
 sky130_fd_sc_hd__and2_1 _18492_ (.A(_06500_),
    .B(net1787),
    .X(_10342_));
 sky130_fd_sc_hd__clkbuf_1 _18493_ (.A(_10342_),
    .X(_10343_));
 sky130_fd_sc_hd__a22o_1 _18494_ (.A1(net1771),
    .A2(net489),
    .B1(net1203),
    .B2(net9027),
    .X(_00440_));
 sky130_fd_sc_hd__buf_1 _18495_ (.A(net1784),
    .X(_10344_));
 sky130_fd_sc_hd__a21oi_1 _18496_ (.A1(net1208),
    .A2(net1441),
    .B1(_10327_),
    .Y(_10345_));
 sky130_fd_sc_hd__or2_1 _18497_ (.A(net874),
    .B(_10345_),
    .X(_10346_));
 sky130_fd_sc_hd__or2_1 _18498_ (.A(_10284_),
    .B(_10287_),
    .X(_10347_));
 sky130_fd_sc_hd__xnor2_1 _18499_ (.A(net6774),
    .B(net2540),
    .Y(_10348_));
 sky130_fd_sc_hd__nor2_2 _18500_ (.A(net6809),
    .B(_09177_),
    .Y(_10349_));
 sky130_fd_sc_hd__nor2_1 _18501_ (.A(net3286),
    .B(net6799),
    .Y(_10350_));
 sky130_fd_sc_hd__nor2_1 _18502_ (.A(_10349_),
    .B(_10350_),
    .Y(_10351_));
 sky130_fd_sc_hd__a211o_1 _18503_ (.A1(_10347_),
    .A2(_10348_),
    .B1(_10351_),
    .C1(_10289_),
    .X(_10352_));
 sky130_fd_sc_hd__or3b_1 _18504_ (.A(net2540),
    .B(_10290_),
    .C_N(_10351_),
    .X(_10353_));
 sky130_fd_sc_hd__and3_1 _18505_ (.A(net6775),
    .B(_10289_),
    .C(_10351_),
    .X(_10354_));
 sky130_fd_sc_hd__a21oi_1 _18506_ (.A1(net3928),
    .A2(_10288_),
    .B1(_10354_),
    .Y(_10355_));
 sky130_fd_sc_hd__and3_1 _18507_ (.A(_10352_),
    .B(_10353_),
    .C(_10355_),
    .X(_10356_));
 sky130_fd_sc_hd__a21o_1 _18508_ (.A1(net3229),
    .A2(_10304_),
    .B1(net3941),
    .X(_10357_));
 sky130_fd_sc_hd__o21ai_1 _18509_ (.A1(net3229),
    .A2(_10304_),
    .B1(_10357_),
    .Y(_10358_));
 sky130_fd_sc_hd__mux2_1 _18510_ (.A0(_09660_),
    .A1(_10304_),
    .S(net3229),
    .X(_10359_));
 sky130_fd_sc_hd__or3b_1 _18511_ (.A(net6982),
    .B(net7070),
    .C_N(net3229),
    .X(_10360_));
 sky130_fd_sc_hd__o2111a_1 _18512_ (.A1(net7076),
    .A2(_10304_),
    .B1(_10359_),
    .C1(_10360_),
    .D1(net6970),
    .X(_10361_));
 sky130_fd_sc_hd__a21oi_1 _18513_ (.A1(net3308),
    .A2(_10358_),
    .B1(_10361_),
    .Y(_10362_));
 sky130_fd_sc_hd__a22o_1 _18514_ (.A1(net3331),
    .A2(_09791_),
    .B1(_10303_),
    .B2(net6970),
    .X(_10363_));
 sky130_fd_sc_hd__xnor2_2 _18515_ (.A(net7013),
    .B(net6915),
    .Y(_10364_));
 sky130_fd_sc_hd__xor2_1 _18516_ (.A(_10171_),
    .B(_10364_),
    .X(_10365_));
 sky130_fd_sc_hd__xnor2_1 _18517_ (.A(net2130),
    .B(_10365_),
    .Y(_10366_));
 sky130_fd_sc_hd__o22a_1 _18518_ (.A1(net3310),
    .A2(net3989),
    .B1(_10063_),
    .B2(net6872),
    .X(_10367_));
 sky130_fd_sc_hd__a211oi_1 _18519_ (.A1(net6872),
    .A2(net3932),
    .B1(_10367_),
    .C1(_10174_),
    .Y(_10368_));
 sky130_fd_sc_hd__nor2_1 _18520_ (.A(net6817),
    .B(net3929),
    .Y(_10369_));
 sky130_fd_sc_hd__a211o_1 _18521_ (.A1(net6818),
    .A2(net6793),
    .B1(_10369_),
    .C1(net6860),
    .X(_10370_));
 sky130_fd_sc_hd__nand2_1 _18522_ (.A(net6818),
    .B(net3929),
    .Y(_10371_));
 sky130_fd_sc_hd__nand2_2 _18523_ (.A(net3285),
    .B(net6793),
    .Y(_10372_));
 sky130_fd_sc_hd__a21o_1 _18524_ (.A1(_10371_),
    .A2(_10372_),
    .B1(net3981),
    .X(_10373_));
 sky130_fd_sc_hd__a21oi_1 _18525_ (.A1(_10371_),
    .A2(_10372_),
    .B1(net6833),
    .Y(_10374_));
 sky130_fd_sc_hd__a31o_1 _18526_ (.A1(net6833),
    .A2(_10370_),
    .A3(_10373_),
    .B1(_10374_),
    .X(_10375_));
 sky130_fd_sc_hd__xnor2_1 _18527_ (.A(net2129),
    .B(_10375_),
    .Y(_10376_));
 sky130_fd_sc_hd__and2_1 _18528_ (.A(net1765),
    .B(_10376_),
    .X(_10377_));
 sky130_fd_sc_hd__or2_1 _18529_ (.A(net1765),
    .B(_10376_),
    .X(_10378_));
 sky130_fd_sc_hd__and2b_1 _18530_ (.A_N(_10377_),
    .B(_10378_),
    .X(_10379_));
 sky130_fd_sc_hd__xnor2_2 _18531_ (.A(net1197),
    .B(_10379_),
    .Y(_10380_));
 sky130_fd_sc_hd__a21o_1 _18532_ (.A1(net1766),
    .A2(net1440),
    .B1(net1207),
    .X(_10381_));
 sky130_fd_sc_hd__o21ai_1 _18533_ (.A1(net1766),
    .A2(net1440),
    .B1(_10381_),
    .Y(_10382_));
 sky130_fd_sc_hd__xnor2_1 _18534_ (.A(_10380_),
    .B(net961),
    .Y(_10383_));
 sky130_fd_sc_hd__xnor2_2 _18535_ (.A(net1071),
    .B(_10383_),
    .Y(_10384_));
 sky130_fd_sc_hd__o21ba_1 _18536_ (.A1(_10322_),
    .A2(net1205),
    .B1_N(_10308_),
    .X(_10385_));
 sky130_fd_sc_hd__a21oi_1 _18537_ (.A1(_10322_),
    .A2(net1205),
    .B1(_10385_),
    .Y(_10386_));
 sky130_fd_sc_hd__inv_2 _18538_ (.A(net3225),
    .Y(_10387_));
 sky130_fd_sc_hd__o21a_1 _18539_ (.A1(_10387_),
    .A2(net2541),
    .B1(_10221_),
    .X(_10388_));
 sky130_fd_sc_hd__a211o_1 _18540_ (.A1(_10387_),
    .A2(net2541),
    .B1(_10388_),
    .C1(net6815),
    .X(_10389_));
 sky130_fd_sc_hd__a21oi_1 _18541_ (.A1(_10387_),
    .A2(_10309_),
    .B1(net2587),
    .Y(_10390_));
 sky130_fd_sc_hd__clkbuf_1 _18542_ (.A(net3930),
    .X(_10391_));
 sky130_fd_sc_hd__a211oi_1 _18543_ (.A1(net3925),
    .A2(_10389_),
    .B1(_10390_),
    .C1(_10391_),
    .Y(_10392_));
 sky130_fd_sc_hd__xnor2_1 _18544_ (.A(_10386_),
    .B(net1436),
    .Y(_10393_));
 sky130_fd_sc_hd__xnor2_1 _18545_ (.A(_10384_),
    .B(_10393_),
    .Y(_10394_));
 sky130_fd_sc_hd__a21oi_1 _18546_ (.A1(_10328_),
    .A2(_10346_),
    .B1(_10394_),
    .Y(_10395_));
 sky130_fd_sc_hd__and3_1 _18547_ (.A(_10328_),
    .B(_10394_),
    .C(_10346_),
    .X(_10396_));
 sky130_fd_sc_hd__nor2_1 _18548_ (.A(_10395_),
    .B(_10396_),
    .Y(_10397_));
 sky130_fd_sc_hd__o21bai_1 _18549_ (.A1(_10332_),
    .A2(_10339_),
    .B1_N(_10333_),
    .Y(_10398_));
 sky130_fd_sc_hd__a2bb2o_1 _18550_ (.A1_N(net607),
    .A2_N(_10398_),
    .B1(_10339_),
    .B2(_10332_),
    .X(_10399_));
 sky130_fd_sc_hd__mux2_1 _18551_ (.A0(_10398_),
    .A1(_10399_),
    .S(net6379),
    .X(_10400_));
 sky130_fd_sc_hd__a31o_1 _18552_ (.A1(net607),
    .A2(_10333_),
    .A3(net765),
    .B1(_10400_),
    .X(_10401_));
 sky130_fd_sc_hd__xor2_1 _18553_ (.A(_10397_),
    .B(_10401_),
    .X(_10402_));
 sky130_fd_sc_hd__nor2_1 _18554_ (.A(net1438),
    .B(net382),
    .Y(_10403_));
 sky130_fd_sc_hd__a31o_1 _18555_ (.A1(net9088),
    .A2(net2289),
    .A3(_09598_),
    .B1(_10403_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _18556_ (.A0(_10333_),
    .A1(_10332_),
    .S(_10397_),
    .X(_10404_));
 sky130_fd_sc_hd__and3_1 _18557_ (.A(_10334_),
    .B(_10339_),
    .C(_10397_),
    .X(_10405_));
 sky130_fd_sc_hd__a21o_1 _18558_ (.A1(net765),
    .A2(_10404_),
    .B1(_10405_),
    .X(_10406_));
 sky130_fd_sc_hd__nand2_1 _18559_ (.A(net607),
    .B(_10406_),
    .Y(_10407_));
 sky130_fd_sc_hd__a21boi_1 _18560_ (.A1(_10384_),
    .A2(net1436),
    .B1_N(_10386_),
    .Y(_10408_));
 sky130_fd_sc_hd__o21ba_1 _18561_ (.A1(_10384_),
    .A2(net1436),
    .B1_N(_10408_),
    .X(_10409_));
 sky130_fd_sc_hd__a21o_1 _18562_ (.A1(_10328_),
    .A2(_10346_),
    .B1(_10394_),
    .X(_10410_));
 sky130_fd_sc_hd__o21a_1 _18563_ (.A1(_10331_),
    .A2(net765),
    .B1(_10410_),
    .X(_10411_));
 sky130_fd_sc_hd__a31o_1 _18564_ (.A1(_10331_),
    .A2(net765),
    .A3(_10410_),
    .B1(_10396_),
    .X(_10412_));
 sky130_fd_sc_hd__a31o_1 _18565_ (.A1(net663),
    .A2(net659),
    .A3(_10411_),
    .B1(_10412_),
    .X(_10413_));
 sky130_fd_sc_hd__a21o_1 _18566_ (.A1(net1071),
    .A2(_10380_),
    .B1(net961),
    .X(_10414_));
 sky130_fd_sc_hd__o21ai_1 _18567_ (.A1(net1071),
    .A2(_10380_),
    .B1(_10414_),
    .Y(_10415_));
 sky130_fd_sc_hd__or2b_1 _18568_ (.A(_10284_),
    .B_N(net2540),
    .X(_10416_));
 sky130_fd_sc_hd__a32o_1 _18569_ (.A1(net6859),
    .A2(_10282_),
    .A3(_10283_),
    .B1(_10287_),
    .B2(_10416_),
    .X(_10417_));
 sky130_fd_sc_hd__a21o_1 _18570_ (.A1(_10372_),
    .A2(_10417_),
    .B1(_10350_),
    .X(_10418_));
 sky130_fd_sc_hd__nand2_1 _18571_ (.A(net6769),
    .B(net1435),
    .Y(_10419_));
 sky130_fd_sc_hd__o21ai_1 _18572_ (.A1(net1197),
    .A2(_10377_),
    .B1(_10378_),
    .Y(_10420_));
 sky130_fd_sc_hd__mux2_1 _18573_ (.A0(_10171_),
    .A1(net3960),
    .S(_10364_),
    .X(_10421_));
 sky130_fd_sc_hd__a211o_1 _18574_ (.A1(_10171_),
    .A2(_10364_),
    .B1(net3308),
    .C1(net6934),
    .X(_10422_));
 sky130_fd_sc_hd__o21ai_1 _18575_ (.A1(net6972),
    .A2(_10421_),
    .B1(_10422_),
    .Y(_10423_));
 sky130_fd_sc_hd__or2_1 _18576_ (.A(net3308),
    .B(_10171_),
    .X(_10424_));
 sky130_fd_sc_hd__nand2_1 _18577_ (.A(net3308),
    .B(_10171_),
    .Y(_10425_));
 sky130_fd_sc_hd__nor3_1 _18578_ (.A(net6934),
    .B(_10171_),
    .C(_10364_),
    .Y(_10426_));
 sky130_fd_sc_hd__a41o_1 _18579_ (.A1(net6934),
    .A2(_10364_),
    .A3(_10424_),
    .A4(_10425_),
    .B1(_10426_),
    .X(_10427_));
 sky130_fd_sc_hd__a21oi_1 _18580_ (.A1(net7044),
    .A2(_10423_),
    .B1(_10427_),
    .Y(_10428_));
 sky130_fd_sc_hd__or2_1 _18581_ (.A(net7016),
    .B(net6952),
    .X(_10429_));
 sky130_fd_sc_hd__mux2_1 _18582_ (.A0(net3945),
    .A1(_10429_),
    .S(net6919),
    .X(_10430_));
 sky130_fd_sc_hd__xnor2_2 _18583_ (.A(net7000),
    .B(net6895),
    .Y(_10431_));
 sky130_fd_sc_hd__xnor2_1 _18584_ (.A(_10430_),
    .B(_10431_),
    .Y(_10432_));
 sky130_fd_sc_hd__xnor2_1 _18585_ (.A(net3225),
    .B(_10432_),
    .Y(_10433_));
 sky130_fd_sc_hd__nand2_1 _18586_ (.A(net6900),
    .B(net3981),
    .Y(_10434_));
 sky130_fd_sc_hd__a221o_1 _18587_ (.A1(net3953),
    .A2(_10434_),
    .B1(net3924),
    .B2(net3299),
    .C1(_10220_),
    .X(_10435_));
 sky130_fd_sc_hd__nand2_1 _18588_ (.A(net6833),
    .B(net6817),
    .Y(_10436_));
 sky130_fd_sc_hd__o21a_1 _18589_ (.A1(net6792),
    .A2(_10436_),
    .B1(_10372_),
    .X(_10437_));
 sky130_fd_sc_hd__xnor2_1 _18590_ (.A(net6786),
    .B(_10437_),
    .Y(_10438_));
 sky130_fd_sc_hd__xnor2_2 _18591_ (.A(net2539),
    .B(_10438_),
    .Y(_10439_));
 sky130_fd_sc_hd__xor2_1 _18592_ (.A(net2128),
    .B(_10439_),
    .X(_10440_));
 sky130_fd_sc_hd__xnor2_2 _18593_ (.A(net1762),
    .B(_10440_),
    .Y(_10441_));
 sky130_fd_sc_hd__or4_1 _18594_ (.A(net6865),
    .B(net2589),
    .C(net6771),
    .D(net2129),
    .X(_10442_));
 sky130_fd_sc_hd__a21oi_1 _18595_ (.A1(net6771),
    .A2(net2129),
    .B1(net3281),
    .Y(_10443_));
 sky130_fd_sc_hd__o22a_1 _18596_ (.A1(net6771),
    .A2(net2129),
    .B1(_10443_),
    .B2(net6818),
    .X(_10444_));
 sky130_fd_sc_hd__a21o_1 _18597_ (.A1(net6860),
    .A2(net3285),
    .B1(net2129),
    .X(_10445_));
 sky130_fd_sc_hd__nor2_1 _18598_ (.A(net3930),
    .B(net3281),
    .Y(_10446_));
 sky130_fd_sc_hd__o211a_1 _18599_ (.A1(net6860),
    .A2(_10369_),
    .B1(_10371_),
    .C1(net2129),
    .X(_10447_));
 sky130_fd_sc_hd__o2bb2a_1 _18600_ (.A1_N(_10445_),
    .A2_N(_10446_),
    .B1(net6793),
    .B2(_10447_),
    .X(_10448_));
 sky130_fd_sc_hd__mux2_1 _18601_ (.A0(_10444_),
    .A1(_10448_),
    .S(net6831),
    .X(_10449_));
 sky130_fd_sc_hd__nand2_1 _18602_ (.A(_10442_),
    .B(_10449_),
    .Y(_10450_));
 sky130_fd_sc_hd__xor2_1 _18603_ (.A(_10441_),
    .B(net1069),
    .X(_10451_));
 sky130_fd_sc_hd__xnor2_1 _18604_ (.A(net1070),
    .B(_10451_),
    .Y(_10452_));
 sky130_fd_sc_hd__and2_1 _18605_ (.A(net1196),
    .B(_10452_),
    .X(_10453_));
 sky130_fd_sc_hd__nor2_1 _18606_ (.A(net1196),
    .B(_10452_),
    .Y(_10454_));
 sky130_fd_sc_hd__or2_1 _18607_ (.A(_10453_),
    .B(_10454_),
    .X(_10455_));
 sky130_fd_sc_hd__xnor2_2 _18608_ (.A(net814),
    .B(_10455_),
    .Y(_10456_));
 sky130_fd_sc_hd__xnor2_1 _18609_ (.A(net605),
    .B(_10456_),
    .Y(_10457_));
 sky130_fd_sc_hd__xnor2_1 _18610_ (.A(net714),
    .B(_10457_),
    .Y(_10458_));
 sky130_fd_sc_hd__a21o_1 _18611_ (.A1(net6377),
    .A2(net422),
    .B1(_10458_),
    .X(_10459_));
 sky130_fd_sc_hd__nand3_1 _18612_ (.A(net6377),
    .B(net422),
    .C(_10458_),
    .Y(_10460_));
 sky130_fd_sc_hd__a32o_1 _18613_ (.A1(net2134),
    .A2(_10459_),
    .A3(_10460_),
    .B1(net1203),
    .B2(net8966),
    .X(_00442_));
 sky130_fd_sc_hd__o21a_1 _18614_ (.A1(net1196),
    .A2(_10452_),
    .B1(net814),
    .X(_10461_));
 sky130_fd_sc_hd__inv_2 _18615_ (.A(_10439_),
    .Y(_10462_));
 sky130_fd_sc_hd__a21o_1 _18616_ (.A1(net2128),
    .A2(_10462_),
    .B1(net1762),
    .X(_10463_));
 sky130_fd_sc_hd__o21ai_2 _18617_ (.A1(net2128),
    .A2(_10462_),
    .B1(_10463_),
    .Y(_10464_));
 sky130_fd_sc_hd__mux2_1 _18618_ (.A0(net6919),
    .A1(_10223_),
    .S(net3959),
    .X(_10465_));
 sky130_fd_sc_hd__nor2_1 _18619_ (.A(_10431_),
    .B(_10465_),
    .Y(_10466_));
 sky130_fd_sc_hd__a31o_1 _18620_ (.A1(net3230),
    .A2(net6957),
    .A3(_10387_),
    .B1(_10466_),
    .X(_10467_));
 sky130_fd_sc_hd__mux2_1 _18621_ (.A0(net3959),
    .A1(_10429_),
    .S(_10223_),
    .X(_10468_));
 sky130_fd_sc_hd__nor3_1 _18622_ (.A(net6919),
    .B(_10223_),
    .C(_10431_),
    .Y(_10469_));
 sky130_fd_sc_hd__a31o_1 _18623_ (.A1(net6929),
    .A2(_10431_),
    .A3(_10468_),
    .B1(_10469_),
    .X(_10470_));
 sky130_fd_sc_hd__a21oi_1 _18624_ (.A1(net7016),
    .A2(_10467_),
    .B1(_10470_),
    .Y(_10471_));
 sky130_fd_sc_hd__or3_1 _18625_ (.A(net3988),
    .B(net6893),
    .C(net3232),
    .X(_10472_));
 sky130_fd_sc_hd__or3_1 _18626_ (.A(net6999),
    .B(net3296),
    .C(net6920),
    .X(_10473_));
 sky130_fd_sc_hd__nand2_1 _18627_ (.A(_10472_),
    .B(_10473_),
    .Y(_10474_));
 sky130_fd_sc_hd__xnor2_2 _18628_ (.A(net6976),
    .B(net6874),
    .Y(_10475_));
 sky130_fd_sc_hd__xor2_1 _18629_ (.A(_10474_),
    .B(_10475_),
    .X(_10476_));
 sky130_fd_sc_hd__xnor2_1 _18630_ (.A(net2131),
    .B(_10476_),
    .Y(_10477_));
 sky130_fd_sc_hd__or2_1 _18631_ (.A(net6827),
    .B(net3966),
    .X(_10478_));
 sky130_fd_sc_hd__nand2_1 _18632_ (.A(net6829),
    .B(net6862),
    .Y(_10479_));
 sky130_fd_sc_hd__o2bb2a_1 _18633_ (.A1_N(_10478_),
    .A2_N(net3938),
    .B1(net6878),
    .B2(_10479_),
    .X(_10480_));
 sky130_fd_sc_hd__o21ai_1 _18634_ (.A1(net6827),
    .A2(net6862),
    .B1(_10480_),
    .Y(_10481_));
 sky130_fd_sc_hd__o21ai_1 _18635_ (.A1(net6813),
    .A2(net6779),
    .B1(net6795),
    .Y(_10482_));
 sky130_fd_sc_hd__xnor2_2 _18636_ (.A(net2127),
    .B(_10482_),
    .Y(_10483_));
 sky130_fd_sc_hd__xnor2_1 _18637_ (.A(net1431),
    .B(_10483_),
    .Y(_10484_));
 sky130_fd_sc_hd__xnor2_2 _18638_ (.A(net1433),
    .B(_10484_),
    .Y(_10485_));
 sky130_fd_sc_hd__nand2_1 _18639_ (.A(net6830),
    .B(net3282),
    .Y(_10486_));
 sky130_fd_sc_hd__nand2_1 _18640_ (.A(net2538),
    .B(net2539),
    .Y(_10487_));
 sky130_fd_sc_hd__mux2_1 _18641_ (.A0(net6792),
    .A1(net6769),
    .S(net2539),
    .X(_10488_));
 sky130_fd_sc_hd__inv_2 _18642_ (.A(_10488_),
    .Y(_10489_));
 sky130_fd_sc_hd__or4_1 _18643_ (.A(net6770),
    .B(net6792),
    .C(net2539),
    .D(_10436_),
    .X(_10490_));
 sky130_fd_sc_hd__o221a_1 _18644_ (.A1(net3223),
    .A2(_10487_),
    .B1(_10489_),
    .B2(net6817),
    .C1(_10490_),
    .X(_10491_));
 sky130_fd_sc_hd__xnor2_1 _18645_ (.A(_10485_),
    .B(_10491_),
    .Y(_10492_));
 sky130_fd_sc_hd__xnor2_2 _18646_ (.A(_10464_),
    .B(_10492_),
    .Y(_10493_));
 sky130_fd_sc_hd__o21ba_1 _18647_ (.A1(_10441_),
    .A2(net1069),
    .B1_N(net1070),
    .X(_10494_));
 sky130_fd_sc_hd__a21o_1 _18648_ (.A1(_10441_),
    .A2(net1069),
    .B1(_10494_),
    .X(_10495_));
 sky130_fd_sc_hd__a22o_1 _18649_ (.A1(net2589),
    .A2(net2129),
    .B1(_10445_),
    .B2(net6831),
    .X(_10496_));
 sky130_fd_sc_hd__and2_1 _18650_ (.A(_10446_),
    .B(_10496_),
    .X(_10497_));
 sky130_fd_sc_hd__xnor2_1 _18651_ (.A(_10495_),
    .B(net1195),
    .Y(_10498_));
 sky130_fd_sc_hd__xnor2_1 _18652_ (.A(_10493_),
    .B(_10498_),
    .Y(_10499_));
 sky130_fd_sc_hd__o21a_1 _18653_ (.A1(_10453_),
    .A2(_10461_),
    .B1(_10499_),
    .X(_10500_));
 sky130_fd_sc_hd__or3_1 _18654_ (.A(_10453_),
    .B(_10499_),
    .C(_10461_),
    .X(_10501_));
 sky130_fd_sc_hd__and2b_1 _18655_ (.A_N(_10500_),
    .B(_10501_),
    .X(_10502_));
 sky130_fd_sc_hd__nand2_1 _18656_ (.A(net605),
    .B(_10456_),
    .Y(_10503_));
 sky130_fd_sc_hd__or2_1 _18657_ (.A(net605),
    .B(_10456_),
    .X(_10504_));
 sky130_fd_sc_hd__clkinvlp_2 _18658_ (.A(_10504_),
    .Y(_10505_));
 sky130_fd_sc_hd__o21ai_1 _18659_ (.A1(net714),
    .A2(_10505_),
    .B1(_10503_),
    .Y(_10506_));
 sky130_fd_sc_hd__a21o_1 _18660_ (.A1(net422),
    .A2(_10503_),
    .B1(_10505_),
    .X(_10507_));
 sky130_fd_sc_hd__a221o_1 _18661_ (.A1(net422),
    .A2(_10505_),
    .B1(_10507_),
    .B2(net714),
    .C1(net3923),
    .X(_10508_));
 sky130_fd_sc_hd__o21ai_1 _18662_ (.A1(net6379),
    .A2(_10506_),
    .B1(_10508_),
    .Y(_10509_));
 sky130_fd_sc_hd__o31a_1 _18663_ (.A1(net422),
    .A2(net714),
    .A3(_10503_),
    .B1(_10509_),
    .X(_10510_));
 sky130_fd_sc_hd__xnor2_1 _18664_ (.A(_10502_),
    .B(_10510_),
    .Y(_10511_));
 sky130_fd_sc_hd__nor2_1 _18665_ (.A(net1437),
    .B(net246),
    .Y(_10512_));
 sky130_fd_sc_hd__a31o_1 _18666_ (.A1(net9075),
    .A2(net2287),
    .A3(net1450),
    .B1(_10512_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _18667_ (.A0(_10503_),
    .A1(_10504_),
    .S(_10502_),
    .X(_10513_));
 sky130_fd_sc_hd__nand2_1 _18668_ (.A(net714),
    .B(_10502_),
    .Y(_10514_));
 sky130_fd_sc_hd__o22a_1 _18669_ (.A1(net714),
    .A2(_10513_),
    .B1(_10514_),
    .B2(_10457_),
    .X(_10515_));
 sky130_fd_sc_hd__nor2_1 _18670_ (.A(_10407_),
    .B(_10515_),
    .Y(_10516_));
 sky130_fd_sc_hd__nor2_1 _18671_ (.A(net3923),
    .B(_10516_),
    .Y(_10517_));
 sky130_fd_sc_hd__a21oi_1 _18672_ (.A1(_10501_),
    .A2(_10506_),
    .B1(_10500_),
    .Y(_10518_));
 sky130_fd_sc_hd__o21a_1 _18673_ (.A1(net1431),
    .A2(_10483_),
    .B1(net1433),
    .X(_10519_));
 sky130_fd_sc_hd__a21o_1 _18674_ (.A1(net1431),
    .A2(_10483_),
    .B1(_10519_),
    .X(_10520_));
 sky130_fd_sc_hd__mux2_1 _18675_ (.A0(net6893),
    .A1(net2131),
    .S(net3231),
    .X(_10521_));
 sky130_fd_sc_hd__inv_2 _18676_ (.A(_10103_),
    .Y(_10522_));
 sky130_fd_sc_hd__mux2_1 _18677_ (.A0(_10521_),
    .A1(_10522_),
    .S(_10475_),
    .X(_10523_));
 sky130_fd_sc_hd__o31a_1 _18678_ (.A1(net6893),
    .A2(net3231),
    .A3(net2131),
    .B1(_10523_),
    .X(_10524_));
 sky130_fd_sc_hd__nor2_1 _18679_ (.A(net3231),
    .B(net2131),
    .Y(_10525_));
 sky130_fd_sc_hd__and2_1 _18680_ (.A(net3231),
    .B(net2131),
    .X(_10526_));
 sky130_fd_sc_hd__or4b_1 _18681_ (.A(net3296),
    .B(_10525_),
    .C(_10526_),
    .D_N(_10475_),
    .X(_10527_));
 sky130_fd_sc_hd__or3_1 _18682_ (.A(net6893),
    .B(net2131),
    .C(_10475_),
    .X(_10528_));
 sky130_fd_sc_hd__o211a_1 _18683_ (.A1(net3988),
    .A2(_10524_),
    .B1(_10527_),
    .C1(_10528_),
    .X(_10529_));
 sky130_fd_sc_hd__nand2_1 _18684_ (.A(net6896),
    .B(net6877),
    .Y(_10530_));
 sky130_fd_sc_hd__nor2_1 _18685_ (.A(net6838),
    .B(net3287),
    .Y(_10531_));
 sky130_fd_sc_hd__xor2_1 _18686_ (.A(_10530_),
    .B(_10531_),
    .X(_10532_));
 sky130_fd_sc_hd__xnor2_2 _18687_ (.A(net6796),
    .B(_10532_),
    .Y(_10533_));
 sky130_fd_sc_hd__xor2_2 _18688_ (.A(net6955),
    .B(net6867),
    .X(_10534_));
 sky130_fd_sc_hd__mux2_1 _18689_ (.A0(net6877),
    .A1(net6896),
    .S(net6975),
    .X(_10535_));
 sky130_fd_sc_hd__xnor2_1 _18690_ (.A(_10534_),
    .B(_10535_),
    .Y(_10536_));
 sky130_fd_sc_hd__xnor2_1 _18691_ (.A(_10533_),
    .B(_10536_),
    .Y(_10537_));
 sky130_fd_sc_hd__nand2_1 _18692_ (.A(net6863),
    .B(net2588),
    .Y(_10538_));
 sky130_fd_sc_hd__nor2_1 _18693_ (.A(net6829),
    .B(net6809),
    .Y(_10539_));
 sky130_fd_sc_hd__a221o_1 _18694_ (.A1(net6820),
    .A2(_10276_),
    .B1(_10285_),
    .B2(_10538_),
    .C1(_10539_),
    .X(_10540_));
 sky130_fd_sc_hd__nand2_1 _18695_ (.A(net6778),
    .B(net1760),
    .Y(_10541_));
 sky130_fd_sc_hd__or2_1 _18696_ (.A(net6778),
    .B(net1760),
    .X(_10542_));
 sky130_fd_sc_hd__nand2_1 _18697_ (.A(_10541_),
    .B(_10542_),
    .Y(_10543_));
 sky130_fd_sc_hd__xor2_1 _18698_ (.A(net1430),
    .B(_10543_),
    .X(_10544_));
 sky130_fd_sc_hd__xnor2_1 _18699_ (.A(net1066),
    .B(_10544_),
    .Y(_10545_));
 sky130_fd_sc_hd__nor2_1 _18700_ (.A(net2588),
    .B(net6785),
    .Y(_10546_));
 sky130_fd_sc_hd__nor2_1 _18701_ (.A(net3282),
    .B(net2127),
    .Y(_10547_));
 sky130_fd_sc_hd__mux2_1 _18702_ (.A0(net6779),
    .A1(net2126),
    .S(_10547_),
    .X(_10548_));
 sky130_fd_sc_hd__nor2_1 _18703_ (.A(_10545_),
    .B(_10548_),
    .Y(_10549_));
 sky130_fd_sc_hd__nand2_1 _18704_ (.A(_10545_),
    .B(_10548_),
    .Y(_10550_));
 sky130_fd_sc_hd__and2b_1 _18705_ (.A_N(_10549_),
    .B(_10550_),
    .X(_10551_));
 sky130_fd_sc_hd__xnor2_2 _18706_ (.A(_10520_),
    .B(_10551_),
    .Y(_10552_));
 sky130_fd_sc_hd__a2bb2o_1 _18707_ (.A1_N(net6792),
    .A2_N(net2539),
    .B1(_10487_),
    .B2(net6812),
    .X(_10553_));
 sky130_fd_sc_hd__nand2_1 _18708_ (.A(net6772),
    .B(_10553_),
    .Y(_10554_));
 sky130_fd_sc_hd__nor2_1 _18709_ (.A(_10485_),
    .B(_10491_),
    .Y(_10555_));
 sky130_fd_sc_hd__nand2_1 _18710_ (.A(_10485_),
    .B(_10491_),
    .Y(_10556_));
 sky130_fd_sc_hd__o21ai_1 _18711_ (.A1(_10464_),
    .A2(_10555_),
    .B1(_10556_),
    .Y(_10557_));
 sky130_fd_sc_hd__and2_1 _18712_ (.A(_10554_),
    .B(_10557_),
    .X(_10558_));
 sky130_fd_sc_hd__nor2_1 _18713_ (.A(_10554_),
    .B(_10557_),
    .Y(_10559_));
 sky130_fd_sc_hd__nor2_1 _18714_ (.A(_10558_),
    .B(_10559_),
    .Y(_10560_));
 sky130_fd_sc_hd__xnor2_2 _18715_ (.A(_10552_),
    .B(_10560_),
    .Y(_10561_));
 sky130_fd_sc_hd__a21bo_1 _18716_ (.A1(_10493_),
    .A2(net1195),
    .B1_N(_10495_),
    .X(_10562_));
 sky130_fd_sc_hd__o21ai_1 _18717_ (.A1(_10493_),
    .A2(net1195),
    .B1(_10562_),
    .Y(_10563_));
 sky130_fd_sc_hd__or2_1 _18718_ (.A(_10561_),
    .B(net764),
    .X(_10564_));
 sky130_fd_sc_hd__nand2_1 _18719_ (.A(_10561_),
    .B(net764),
    .Y(_10565_));
 sky130_fd_sc_hd__nand2_1 _18720_ (.A(_10564_),
    .B(_10565_),
    .Y(_10566_));
 sky130_fd_sc_hd__xor2_1 _18721_ (.A(net421),
    .B(_10566_),
    .X(_10567_));
 sky130_fd_sc_hd__xnor2_1 _18722_ (.A(_10517_),
    .B(_10567_),
    .Y(_10568_));
 sky130_fd_sc_hd__a22o_1 _18723_ (.A1(net9016),
    .A2(net1203),
    .B1(_10568_),
    .B2(net1771),
    .X(_00444_));
 sky130_fd_sc_hd__nor2_1 _18724_ (.A(_10552_),
    .B(_10559_),
    .Y(_10569_));
 sky130_fd_sc_hd__inv_2 _18725_ (.A(net1066),
    .Y(_10570_));
 sky130_fd_sc_hd__a21o_1 _18726_ (.A1(_10570_),
    .A2(net1430),
    .B1(_10543_),
    .X(_10571_));
 sky130_fd_sc_hd__o21a_1 _18727_ (.A1(_10570_),
    .A2(net1430),
    .B1(_10571_),
    .X(_10572_));
 sky130_fd_sc_hd__nand2_1 _18728_ (.A(net6877),
    .B(_10534_),
    .Y(_10573_));
 sky130_fd_sc_hd__or2_1 _18729_ (.A(net6877),
    .B(_10534_),
    .X(_10574_));
 sky130_fd_sc_hd__mux2_1 _18730_ (.A0(net6877),
    .A1(_10533_),
    .S(_10534_),
    .X(_10575_));
 sky130_fd_sc_hd__o211a_1 _18731_ (.A1(_10533_),
    .A2(_10534_),
    .B1(_10573_),
    .C1(net6896),
    .X(_10576_));
 sky130_fd_sc_hd__a21o_1 _18732_ (.A1(net3298),
    .A2(_10575_),
    .B1(_10576_),
    .X(_10577_));
 sky130_fd_sc_hd__a32o_1 _18733_ (.A1(_10533_),
    .A2(_10573_),
    .A3(_10574_),
    .B1(_10577_),
    .B2(net6975),
    .X(_10578_));
 sky130_fd_sc_hd__xnor2_2 _18734_ (.A(net6784),
    .B(_10349_),
    .Y(_10579_));
 sky130_fd_sc_hd__or2_1 _18735_ (.A(net6955),
    .B(net6878),
    .X(_10580_));
 sky130_fd_sc_hd__mux2_1 _18736_ (.A0(net3985),
    .A1(_10580_),
    .S(net6855),
    .X(_10581_));
 sky130_fd_sc_hd__nor2_1 _18737_ (.A(net3231),
    .B(net6826),
    .Y(_10582_));
 sky130_fd_sc_hd__and2_1 _18738_ (.A(net3231),
    .B(net6826),
    .X(_10583_));
 sky130_fd_sc_hd__nor2_1 _18739_ (.A(_10582_),
    .B(_10583_),
    .Y(_10584_));
 sky130_fd_sc_hd__xor2_1 _18740_ (.A(_10581_),
    .B(_10584_),
    .X(_10585_));
 sky130_fd_sc_hd__xnor2_1 _18741_ (.A(_10579_),
    .B(_10585_),
    .Y(_10586_));
 sky130_fd_sc_hd__nor2_1 _18742_ (.A(net6813),
    .B(net6796),
    .Y(_10587_));
 sky130_fd_sc_hd__a221o_1 _18743_ (.A1(_10530_),
    .A2(_10486_),
    .B1(_10531_),
    .B2(net6796),
    .C1(_10587_),
    .X(_10588_));
 sky130_fd_sc_hd__nand2_1 _18744_ (.A(net6781),
    .B(net2125),
    .Y(_10589_));
 sky130_fd_sc_hd__or2_1 _18745_ (.A(net6781),
    .B(net2125),
    .X(_10590_));
 sky130_fd_sc_hd__and2_1 _18746_ (.A(_10589_),
    .B(_10590_),
    .X(_10591_));
 sky130_fd_sc_hd__xor2_1 _18747_ (.A(net1429),
    .B(_10591_),
    .X(_10592_));
 sky130_fd_sc_hd__xnor2_2 _18748_ (.A(net1065),
    .B(_10592_),
    .Y(_10593_));
 sky130_fd_sc_hd__xor2_1 _18749_ (.A(_10541_),
    .B(_10593_),
    .X(_10594_));
 sky130_fd_sc_hd__xnor2_1 _18750_ (.A(_10572_),
    .B(_10594_),
    .Y(_10595_));
 sky130_fd_sc_hd__o21ai_2 _18751_ (.A1(_10520_),
    .A2(_10549_),
    .B1(_10550_),
    .Y(_10596_));
 sky130_fd_sc_hd__nand2_1 _18752_ (.A(net6779),
    .B(net6795),
    .Y(_10597_));
 sky130_fd_sc_hd__nor2_1 _18753_ (.A(_10597_),
    .B(net2127),
    .Y(_10598_));
 sky130_fd_sc_hd__xnor2_1 _18754_ (.A(_10596_),
    .B(_10598_),
    .Y(_10599_));
 sky130_fd_sc_hd__xor2_1 _18755_ (.A(_10595_),
    .B(_10599_),
    .X(_10600_));
 sky130_fd_sc_hd__o21ai_1 _18756_ (.A1(_10558_),
    .A2(_10569_),
    .B1(_10600_),
    .Y(_10601_));
 sky130_fd_sc_hd__or3_1 _18757_ (.A(_10558_),
    .B(_10600_),
    .C(_10569_),
    .X(_10602_));
 sky130_fd_sc_hd__and2_1 _18758_ (.A(_10601_),
    .B(_10602_),
    .X(_10603_));
 sky130_fd_sc_hd__nor2_1 _18759_ (.A(net421),
    .B(_10565_),
    .Y(_10604_));
 sky130_fd_sc_hd__a21o_1 _18760_ (.A1(_10516_),
    .A2(net764),
    .B1(_10561_),
    .X(_10605_));
 sky130_fd_sc_hd__o21ai_1 _18761_ (.A1(_10516_),
    .A2(net764),
    .B1(_10605_),
    .Y(_10606_));
 sky130_fd_sc_hd__a2bb2o_1 _18762_ (.A1_N(_10516_),
    .A2_N(_10564_),
    .B1(_10606_),
    .B2(net421),
    .X(_10607_));
 sky130_fd_sc_hd__inv_2 _18763_ (.A(net714),
    .Y(_10608_));
 sky130_fd_sc_hd__and2_1 _18764_ (.A(_10501_),
    .B(_10564_),
    .X(_10609_));
 sky130_fd_sc_hd__o211a_1 _18765_ (.A1(_10608_),
    .A2(_10456_),
    .B1(_10609_),
    .C1(net605),
    .X(_10610_));
 sky130_fd_sc_hd__a32o_1 _18766_ (.A1(_10608_),
    .A2(_10456_),
    .A3(_10609_),
    .B1(_10564_),
    .B2(_10500_),
    .X(_10611_));
 sky130_fd_sc_hd__or2_1 _18767_ (.A(_10610_),
    .B(_10611_),
    .X(_10612_));
 sky130_fd_sc_hd__a21o_1 _18768_ (.A1(_10561_),
    .A2(net764),
    .B1(net526),
    .X(_10613_));
 sky130_fd_sc_hd__mux2_1 _18769_ (.A0(_10607_),
    .A1(_10613_),
    .S(_10335_),
    .X(_10614_));
 sky130_fd_sc_hd__a21oi_1 _18770_ (.A1(_10516_),
    .A2(_10604_),
    .B1(_10614_),
    .Y(_10615_));
 sky130_fd_sc_hd__xnor2_1 _18771_ (.A(_10603_),
    .B(_10615_),
    .Y(_10616_));
 sky130_fd_sc_hd__nor2_1 _18772_ (.A(net1437),
    .B(net180),
    .Y(_10617_));
 sky130_fd_sc_hd__a31o_1 _18773_ (.A1(net9064),
    .A2(net2287),
    .A3(net1450),
    .B1(_10617_),
    .X(_00445_));
 sky130_fd_sc_hd__or2_1 _18774_ (.A(net764),
    .B(_10600_),
    .X(_10618_));
 sky130_fd_sc_hd__nand2_1 _18775_ (.A(net764),
    .B(_10603_),
    .Y(_10619_));
 sky130_fd_sc_hd__a21bo_1 _18776_ (.A1(_10601_),
    .A2(_10602_),
    .B1_N(net764),
    .X(_10620_));
 sky130_fd_sc_hd__or2b_1 _18777_ (.A(net764),
    .B_N(_10603_),
    .X(_10621_));
 sky130_fd_sc_hd__mux4_1 _18778_ (.A0(_10618_),
    .A1(_10619_),
    .A2(_10620_),
    .A3(_10621_),
    .S0(net421),
    .S1(_10561_),
    .X(_10622_));
 sky130_fd_sc_hd__or3_1 _18779_ (.A(_10407_),
    .B(_10515_),
    .C(_10622_),
    .X(_10623_));
 sky130_fd_sc_hd__nand2_1 _18780_ (.A(_10565_),
    .B(_10601_),
    .Y(_10624_));
 sky130_fd_sc_hd__o21ai_1 _18781_ (.A1(net526),
    .A2(_10624_),
    .B1(_10602_),
    .Y(_10625_));
 sky130_fd_sc_hd__a21bo_1 _18782_ (.A1(_10572_),
    .A2(_10593_),
    .B1_N(_10541_),
    .X(_10626_));
 sky130_fd_sc_hd__o21a_1 _18783_ (.A1(_10572_),
    .A2(_10593_),
    .B1(_10626_),
    .X(_10627_));
 sky130_fd_sc_hd__a21bo_1 _18784_ (.A1(net1065),
    .A2(net1429),
    .B1_N(_10591_),
    .X(_10628_));
 sky130_fd_sc_hd__o21ai_2 _18785_ (.A1(net1065),
    .A2(net1429),
    .B1(_10628_),
    .Y(_10629_));
 sky130_fd_sc_hd__mux2_1 _18786_ (.A0(net6862),
    .A1(_10579_),
    .S(net3967),
    .X(_10630_));
 sky130_fd_sc_hd__or2_1 _18787_ (.A(_10584_),
    .B(_10630_),
    .X(_10631_));
 sky130_fd_sc_hd__o31a_1 _18788_ (.A1(net6862),
    .A2(net3967),
    .A3(_10579_),
    .B1(_10631_),
    .X(_10632_));
 sky130_fd_sc_hd__mux2_1 _18789_ (.A0(net3967),
    .A1(_10580_),
    .S(_10579_),
    .X(_10633_));
 sky130_fd_sc_hd__nor3_1 _18790_ (.A(net6855),
    .B(_10579_),
    .C(_10584_),
    .Y(_10634_));
 sky130_fd_sc_hd__a31o_1 _18791_ (.A1(net6855),
    .A2(_10584_),
    .A3(_10633_),
    .B1(_10634_),
    .X(_10635_));
 sky130_fd_sc_hd__o21ba_1 _18792_ (.A1(net3957),
    .A2(_10632_),
    .B1_N(_10635_),
    .X(_10636_));
 sky130_fd_sc_hd__mux2_1 _18793_ (.A0(_10582_),
    .A1(_10583_),
    .S(net3983),
    .X(_10637_));
 sky130_fd_sc_hd__xnor2_2 _18794_ (.A(net6897),
    .B(net6808),
    .Y(_10638_));
 sky130_fd_sc_hd__xnor2_1 _18795_ (.A(net3920),
    .B(_10638_),
    .Y(_10639_));
 sky130_fd_sc_hd__xnor2_1 _18796_ (.A(_10637_),
    .B(_10639_),
    .Y(_10640_));
 sky130_fd_sc_hd__nand2_1 _18797_ (.A(net6867),
    .B(net6878),
    .Y(_10641_));
 sky130_fd_sc_hd__a21o_1 _18798_ (.A1(net2588),
    .A2(_10218_),
    .B1(_10546_),
    .X(_10642_));
 sky130_fd_sc_hd__a22o_1 _18799_ (.A1(net6784),
    .A2(_10641_),
    .B1(_10642_),
    .B2(net6800),
    .X(_10643_));
 sky130_fd_sc_hd__nor2_1 _18800_ (.A(_10640_),
    .B(_10643_),
    .Y(_10644_));
 sky130_fd_sc_hd__nand2_1 _18801_ (.A(_10640_),
    .B(_10643_),
    .Y(_10645_));
 sky130_fd_sc_hd__or2b_1 _18802_ (.A(_10644_),
    .B_N(_10645_),
    .X(_10646_));
 sky130_fd_sc_hd__xnor2_2 _18803_ (.A(_10636_),
    .B(_10646_),
    .Y(_10647_));
 sky130_fd_sc_hd__xor2_1 _18804_ (.A(_10589_),
    .B(_10647_),
    .X(_10648_));
 sky130_fd_sc_hd__xnor2_2 _18805_ (.A(_10629_),
    .B(_10648_),
    .Y(_10649_));
 sky130_fd_sc_hd__nor2_1 _18806_ (.A(net3221),
    .B(net1760),
    .Y(_10650_));
 sky130_fd_sc_hd__xor2_1 _18807_ (.A(_10649_),
    .B(_10650_),
    .X(_10651_));
 sky130_fd_sc_hd__xnor2_1 _18808_ (.A(_10627_),
    .B(_10651_),
    .Y(_10652_));
 sky130_fd_sc_hd__a21o_1 _18809_ (.A1(_10596_),
    .A2(_10598_),
    .B1(_10595_),
    .X(_10653_));
 sky130_fd_sc_hd__o21ai_2 _18810_ (.A1(_10596_),
    .A2(_10598_),
    .B1(_10653_),
    .Y(_10654_));
 sky130_fd_sc_hd__xor2_1 _18811_ (.A(_10652_),
    .B(_10654_),
    .X(_10655_));
 sky130_fd_sc_hd__xnor2_1 _18812_ (.A(_10625_),
    .B(_10655_),
    .Y(_10656_));
 sky130_fd_sc_hd__a21oi_1 _18813_ (.A1(net6376),
    .A2(_10623_),
    .B1(_10656_),
    .Y(_10657_));
 sky130_fd_sc_hd__and3_1 _18814_ (.A(net6376),
    .B(_10656_),
    .C(_10623_),
    .X(_10658_));
 sky130_fd_sc_hd__o21a_1 _18815_ (.A1(_10657_),
    .A2(_10658_),
    .B1(net2132),
    .X(_10659_));
 sky130_fd_sc_hd__a31o_1 _18816_ (.A1(net9098),
    .A2(net2288),
    .A3(net1449),
    .B1(_10659_),
    .X(_00446_));
 sky130_fd_sc_hd__inv_2 _18817_ (.A(_10654_),
    .Y(_10660_));
 sky130_fd_sc_hd__o21bai_1 _18818_ (.A1(_10625_),
    .A2(_10660_),
    .B1_N(_10652_),
    .Y(_10661_));
 sky130_fd_sc_hd__a21o_1 _18819_ (.A1(_10627_),
    .A2(_10649_),
    .B1(_10650_),
    .X(_10662_));
 sky130_fd_sc_hd__o21ai_1 _18820_ (.A1(_10627_),
    .A2(_10649_),
    .B1(_10662_),
    .Y(_10663_));
 sky130_fd_sc_hd__and2_1 _18821_ (.A(_10661_),
    .B(_10663_),
    .X(_10664_));
 sky130_fd_sc_hd__nand2_1 _18822_ (.A(_10661_),
    .B(_10663_),
    .Y(_10665_));
 sky130_fd_sc_hd__a21o_1 _18823_ (.A1(_10636_),
    .A2(_10645_),
    .B1(_10644_),
    .X(_10666_));
 sky130_fd_sc_hd__mux2_1 _18824_ (.A0(net6837),
    .A1(net3920),
    .S(net3983),
    .X(_10667_));
 sky130_fd_sc_hd__nor2_1 _18825_ (.A(_10638_),
    .B(_10667_),
    .Y(_10668_));
 sky130_fd_sc_hd__nor2_1 _18826_ (.A(net6826),
    .B(net3920),
    .Y(_10669_));
 sky130_fd_sc_hd__a22o_1 _18827_ (.A1(_10276_),
    .A2(_10638_),
    .B1(_10669_),
    .B2(net6855),
    .X(_10670_));
 sky130_fd_sc_hd__o21ai_1 _18828_ (.A1(_10668_),
    .A2(_10670_),
    .B1(net6921),
    .Y(_10671_));
 sky130_fd_sc_hd__xnor2_1 _18829_ (.A(net6868),
    .B(net3920),
    .Y(_10672_));
 sky130_fd_sc_hd__nand3_1 _18830_ (.A(net6837),
    .B(_10638_),
    .C(_10672_),
    .Y(_10673_));
 sky130_fd_sc_hd__o311a_1 _18831_ (.A1(net6837),
    .A2(net3920),
    .A3(_10638_),
    .B1(_10671_),
    .C1(_10673_),
    .X(_10674_));
 sky130_fd_sc_hd__and3_1 _18832_ (.A(net6896),
    .B(net6829),
    .C(net2588),
    .X(_10675_));
 sky130_fd_sc_hd__a21oi_1 _18833_ (.A1(net3298),
    .A2(_10531_),
    .B1(_10675_),
    .Y(_10676_));
 sky130_fd_sc_hd__xor2_4 _18834_ (.A(net6877),
    .B(net6796),
    .X(_10677_));
 sky130_fd_sc_hd__xnor2_1 _18835_ (.A(net3222),
    .B(_10677_),
    .Y(_10678_));
 sky130_fd_sc_hd__xnor2_2 _18836_ (.A(_10676_),
    .B(_10678_),
    .Y(_10679_));
 sky130_fd_sc_hd__o21ai_4 _18837_ (.A1(net3282),
    .A2(net3922),
    .B1(net6779),
    .Y(_10680_));
 sky130_fd_sc_hd__xnor2_1 _18838_ (.A(_10679_),
    .B(_10680_),
    .Y(_10681_));
 sky130_fd_sc_hd__xnor2_1 _18839_ (.A(net1428),
    .B(_10681_),
    .Y(_10682_));
 sky130_fd_sc_hd__nor2_1 _18840_ (.A(_10641_),
    .B(_10349_),
    .Y(_10683_));
 sky130_fd_sc_hd__or2_1 _18841_ (.A(net3222),
    .B(_10683_),
    .X(_10684_));
 sky130_fd_sc_hd__xnor2_1 _18842_ (.A(_10682_),
    .B(_10684_),
    .Y(_10685_));
 sky130_fd_sc_hd__xnor2_2 _18843_ (.A(_10666_),
    .B(_10685_),
    .Y(_10686_));
 sky130_fd_sc_hd__inv_2 _18844_ (.A(net2125),
    .Y(_10687_));
 sky130_fd_sc_hd__nor2_1 _18845_ (.A(_10629_),
    .B(_10647_),
    .Y(_10688_));
 sky130_fd_sc_hd__nand2_1 _18846_ (.A(_10629_),
    .B(_10647_),
    .Y(_10689_));
 sky130_fd_sc_hd__o22ai_1 _18847_ (.A1(net6781),
    .A2(_10688_),
    .B1(_10689_),
    .B2(_10687_),
    .Y(_10690_));
 sky130_fd_sc_hd__a31o_1 _18848_ (.A1(net6781),
    .A2(_10687_),
    .A3(_10688_),
    .B1(_10690_),
    .X(_10691_));
 sky130_fd_sc_hd__xor2_1 _18849_ (.A(_10686_),
    .B(_10691_),
    .X(_10692_));
 sky130_fd_sc_hd__mux2_1 _18850_ (.A0(_10664_),
    .A1(_10665_),
    .S(net658),
    .X(_10693_));
 sky130_fd_sc_hd__nand2b_1 _18851_ (.A_N(_10623_),
    .B(_10656_),
    .Y(_10694_));
 sky130_fd_sc_hd__nand2_1 _18852_ (.A(net6376),
    .B(_10694_),
    .Y(_10695_));
 sky130_fd_sc_hd__or2_1 _18853_ (.A(net352),
    .B(_10695_),
    .X(_10696_));
 sky130_fd_sc_hd__nand2_1 _18854_ (.A(net352),
    .B(_10695_),
    .Y(_10697_));
 sky130_fd_sc_hd__a21oi_1 _18855_ (.A1(_10696_),
    .A2(_10697_),
    .B1(net1443),
    .Y(_10698_));
 sky130_fd_sc_hd__a31o_1 _18856_ (.A1(net9085),
    .A2(net2288),
    .A3(net1449),
    .B1(_10698_),
    .X(_00447_));
 sky130_fd_sc_hd__nor2_1 _18857_ (.A(net658),
    .B(_10664_),
    .Y(_10699_));
 sky130_fd_sc_hd__nor2_1 _18858_ (.A(_10686_),
    .B(_10688_),
    .Y(_10700_));
 sky130_fd_sc_hd__o2bb2a_1 _18859_ (.A1_N(_10686_),
    .A2_N(_10689_),
    .B1(_10700_),
    .B2(net2125),
    .X(_10701_));
 sky130_fd_sc_hd__o2bb2a_1 _18860_ (.A1_N(_10686_),
    .A2_N(_10688_),
    .B1(_10701_),
    .B2(net3221),
    .X(_10702_));
 sky130_fd_sc_hd__inv_2 _18861_ (.A(_10679_),
    .Y(_10703_));
 sky130_fd_sc_hd__o21a_1 _18862_ (.A1(_10703_),
    .A2(_10680_),
    .B1(net1428),
    .X(_10704_));
 sky130_fd_sc_hd__a21o_1 _18863_ (.A1(_10703_),
    .A2(_10680_),
    .B1(_10704_),
    .X(_10705_));
 sky130_fd_sc_hd__mux2_1 _18864_ (.A0(net6812),
    .A1(net6770),
    .S(_10677_),
    .X(_10706_));
 sky130_fd_sc_hd__o21a_1 _18865_ (.A1(net6770),
    .A2(_10677_),
    .B1(net2589),
    .X(_10707_));
 sky130_fd_sc_hd__mux2_1 _18866_ (.A0(_10706_),
    .A1(_10707_),
    .S(net6834),
    .X(_10708_));
 sky130_fd_sc_hd__and2_1 _18867_ (.A(net6832),
    .B(net3224),
    .X(_10709_));
 sky130_fd_sc_hd__nor2_1 _18868_ (.A(net6832),
    .B(net3224),
    .Y(_10710_));
 sky130_fd_sc_hd__or2_1 _18869_ (.A(_10709_),
    .B(_10710_),
    .X(_10711_));
 sky130_fd_sc_hd__nor3b_1 _18870_ (.A(net2589),
    .B(_10677_),
    .C_N(_10711_),
    .Y(_10712_));
 sky130_fd_sc_hd__a221o_1 _18871_ (.A1(_10369_),
    .A2(_10677_),
    .B1(_10708_),
    .B2(net6898),
    .C1(_10712_),
    .X(_10713_));
 sky130_fd_sc_hd__or2_1 _18872_ (.A(net6881),
    .B(net6814),
    .X(_10714_));
 sky130_fd_sc_hd__mux2_1 _18873_ (.A0(net3934),
    .A1(_10714_),
    .S(net6794),
    .X(_10715_));
 sky130_fd_sc_hd__xnor2_2 _18874_ (.A(net6860),
    .B(_10715_),
    .Y(_10716_));
 sky130_fd_sc_hd__nand2_1 _18875_ (.A(net6770),
    .B(_10436_),
    .Y(_10717_));
 sky130_fd_sc_hd__nor2_1 _18876_ (.A(_10716_),
    .B(_10717_),
    .Y(_10718_));
 sky130_fd_sc_hd__and2_1 _18877_ (.A(_10716_),
    .B(_10717_),
    .X(_10719_));
 sky130_fd_sc_hd__or2_1 _18878_ (.A(_10718_),
    .B(_10719_),
    .X(_10720_));
 sky130_fd_sc_hd__xnor2_1 _18879_ (.A(_10713_),
    .B(_10720_),
    .Y(_10721_));
 sky130_fd_sc_hd__xnor2_1 _18880_ (.A(_10680_),
    .B(net1194),
    .Y(_10722_));
 sky130_fd_sc_hd__xnor2_2 _18881_ (.A(_10705_),
    .B(_10722_),
    .Y(_10723_));
 sky130_fd_sc_hd__o21ai_1 _18882_ (.A1(_10682_),
    .A2(_10683_),
    .B1(net6781),
    .Y(_10724_));
 sky130_fd_sc_hd__a2bb2o_1 _18883_ (.A1_N(net6781),
    .A2_N(_10682_),
    .B1(_10724_),
    .B2(_10666_),
    .X(_10725_));
 sky130_fd_sc_hd__xnor2_1 _18884_ (.A(_10723_),
    .B(net873),
    .Y(_10726_));
 sky130_fd_sc_hd__xnor2_1 _18885_ (.A(net657),
    .B(_10726_),
    .Y(_10727_));
 sky130_fd_sc_hd__xnor2_1 _18886_ (.A(_10699_),
    .B(_10727_),
    .Y(_10728_));
 sky130_fd_sc_hd__or2_1 _18887_ (.A(net352),
    .B(_10694_),
    .X(_10729_));
 sky130_fd_sc_hd__nand2_1 _18888_ (.A(net6376),
    .B(_10729_),
    .Y(_10730_));
 sky130_fd_sc_hd__xor2_1 _18889_ (.A(net302),
    .B(_10730_),
    .X(_10731_));
 sky130_fd_sc_hd__nor2_1 _18890_ (.A(net1437),
    .B(_10731_),
    .Y(_10732_));
 sky130_fd_sc_hd__a31o_1 _18891_ (.A1(net9076),
    .A2(net2287),
    .A3(net1450),
    .B1(_10732_),
    .X(_00448_));
 sky130_fd_sc_hd__or2_1 _18892_ (.A(_10705_),
    .B(net1194),
    .X(_10733_));
 sky130_fd_sc_hd__and2_1 _18893_ (.A(_10705_),
    .B(net1194),
    .X(_10734_));
 sky130_fd_sc_hd__a21oi_1 _18894_ (.A1(_10680_),
    .A2(_10733_),
    .B1(_10734_),
    .Y(_10735_));
 sky130_fd_sc_hd__nand2_1 _18895_ (.A(net3283),
    .B(net3934),
    .Y(_10736_));
 sky130_fd_sc_hd__a22o_1 _18896_ (.A1(net6794),
    .A2(_10714_),
    .B1(_10736_),
    .B2(net6860),
    .X(_10737_));
 sky130_fd_sc_hd__xor2_2 _18897_ (.A(_10711_),
    .B(_10737_),
    .X(_10738_));
 sky130_fd_sc_hd__mux2_1 _18898_ (.A0(_10718_),
    .A1(_10719_),
    .S(_10713_),
    .X(_10739_));
 sky130_fd_sc_hd__xor2_1 _18899_ (.A(_10738_),
    .B(_10739_),
    .X(_10740_));
 sky130_fd_sc_hd__a2bb2o_1 _18900_ (.A1_N(net3922),
    .A2_N(_10597_),
    .B1(_10735_),
    .B2(_10740_),
    .X(_10741_));
 sky130_fd_sc_hd__or2_1 _18901_ (.A(_10735_),
    .B(_10740_),
    .X(_10742_));
 sky130_fd_sc_hd__or2b_1 _18902_ (.A(_10741_),
    .B_N(_10742_),
    .X(_10743_));
 sky130_fd_sc_hd__o221a_1 _18903_ (.A1(net658),
    .A2(_10664_),
    .B1(_10723_),
    .B2(net873),
    .C1(net657),
    .X(_10744_));
 sky130_fd_sc_hd__a21oi_1 _18904_ (.A1(_10723_),
    .A2(net873),
    .B1(_10744_),
    .Y(_10745_));
 sky130_fd_sc_hd__xnor2_1 _18905_ (.A(_10743_),
    .B(_10745_),
    .Y(_10746_));
 sky130_fd_sc_hd__or2_1 _18906_ (.A(net302),
    .B(_10729_),
    .X(_10747_));
 sky130_fd_sc_hd__or3b_1 _18907_ (.A(_10335_),
    .B(net275),
    .C_N(_10747_),
    .X(_10748_));
 sky130_fd_sc_hd__a21bo_1 _18908_ (.A1(net6376),
    .A2(_10747_),
    .B1_N(net275),
    .X(_10749_));
 sky130_fd_sc_hd__a21oi_1 _18909_ (.A1(_10748_),
    .A2(_10749_),
    .B1(net1443),
    .Y(_10750_));
 sky130_fd_sc_hd__a31o_1 _18910_ (.A1(net9062),
    .A2(net2288),
    .A3(net1449),
    .B1(_10750_),
    .X(_00449_));
 sky130_fd_sc_hd__nor2_1 _18911_ (.A(net6876),
    .B(net6814),
    .Y(_10751_));
 sky130_fd_sc_hd__a221oi_1 _18912_ (.A1(_10278_),
    .A2(_10531_),
    .B1(_10751_),
    .B2(net6828),
    .C1(net6864),
    .Y(_10752_));
 sky130_fd_sc_hd__o221a_1 _18913_ (.A1(_10123_),
    .A2(_10371_),
    .B1(_10372_),
    .B2(net6832),
    .C1(net6859),
    .X(_10753_));
 sky130_fd_sc_hd__nor2_1 _18914_ (.A(net6828),
    .B(net6876),
    .Y(_10754_));
 sky130_fd_sc_hd__a22o_1 _18915_ (.A1(net6828),
    .A2(_10279_),
    .B1(_10754_),
    .B2(_10278_),
    .X(_10755_));
 sky130_fd_sc_hd__nand2_1 _18916_ (.A(net6814),
    .B(_10755_),
    .Y(_10756_));
 sky130_fd_sc_hd__nand2_1 _18917_ (.A(net6876),
    .B(net6801),
    .Y(_10757_));
 sky130_fd_sc_hd__a221o_1 _18918_ (.A1(net6828),
    .A2(_10279_),
    .B1(_10710_),
    .B2(_10757_),
    .C1(net6814),
    .X(_10758_));
 sky130_fd_sc_hd__o211a_1 _18919_ (.A1(_10752_),
    .A2(_10753_),
    .B1(_10756_),
    .C1(_10758_),
    .X(_10759_));
 sky130_fd_sc_hd__nor2_1 _18920_ (.A(_10716_),
    .B(_10738_),
    .Y(_10760_));
 sky130_fd_sc_hd__a21o_1 _18921_ (.A1(_10716_),
    .A2(_10738_),
    .B1(net6777),
    .X(_10761_));
 sky130_fd_sc_hd__a2bb2o_1 _18922_ (.A1_N(_10717_),
    .A2_N(_10760_),
    .B1(_10761_),
    .B2(_10713_),
    .X(_10762_));
 sky130_fd_sc_hd__a2bb2o_1 _18923_ (.A1_N(net3223),
    .A2_N(_10436_),
    .B1(net1427),
    .B2(_10762_),
    .X(_10763_));
 sky130_fd_sc_hd__o21ba_1 _18924_ (.A1(net1427),
    .A2(_10762_),
    .B1_N(_10763_),
    .X(_10764_));
 sky130_fd_sc_hd__a21o_1 _18925_ (.A1(_10742_),
    .A2(_10745_),
    .B1(_10741_),
    .X(_10765_));
 sky130_fd_sc_hd__xor2_1 _18926_ (.A(_10764_),
    .B(_10765_),
    .X(_10766_));
 sky130_fd_sc_hd__o21a_1 _18927_ (.A1(net275),
    .A2(_10747_),
    .B1(net6376),
    .X(_10767_));
 sky130_fd_sc_hd__xnor2_1 _18928_ (.A(net245),
    .B(_10767_),
    .Y(_10768_));
 sky130_fd_sc_hd__nor2_1 _18929_ (.A(net1437),
    .B(_10768_),
    .Y(_10769_));
 sky130_fd_sc_hd__a31o_1 _18930_ (.A1(net9074),
    .A2(net2287),
    .A3(net1450),
    .B1(_10769_),
    .X(_00450_));
 sky130_fd_sc_hd__buf_1 _18931_ (.A(_06500_),
    .X(_10770_));
 sky130_fd_sc_hd__clkbuf_1 _18932_ (.A(net2537),
    .X(_10771_));
 sky130_fd_sc_hd__or3_1 _18933_ (.A(net275),
    .B(_10747_),
    .C(net245),
    .X(_10772_));
 sky130_fd_sc_hd__a21oi_1 _18934_ (.A1(net3982),
    .A2(_10751_),
    .B1(net3224),
    .Y(_10773_));
 sky130_fd_sc_hd__o221a_1 _18935_ (.A1(net6816),
    .A2(net6779),
    .B1(_10773_),
    .B2(net6830),
    .C1(net6794),
    .X(_10774_));
 sky130_fd_sc_hd__a31o_1 _18936_ (.A1(net6863),
    .A2(net6878),
    .A3(net6813),
    .B1(net6779),
    .X(_10775_));
 sky130_fd_sc_hd__a221o_1 _18937_ (.A1(net6813),
    .A2(net6779),
    .B1(_10775_),
    .B2(net6830),
    .C1(net6796),
    .X(_10776_));
 sky130_fd_sc_hd__and2b_1 _18938_ (.A_N(_10774_),
    .B(_10776_),
    .X(_10777_));
 sky130_fd_sc_hd__xnor2_1 _18939_ (.A(_10763_),
    .B(_10777_),
    .Y(_10778_));
 sky130_fd_sc_hd__a21oi_1 _18940_ (.A1(_10764_),
    .A2(_10765_),
    .B1(_10778_),
    .Y(_10779_));
 sky130_fd_sc_hd__a31oi_1 _18941_ (.A1(_10764_),
    .A2(_10765_),
    .A3(_10778_),
    .B1(_10779_),
    .Y(_10780_));
 sky130_fd_sc_hd__a21oi_1 _18942_ (.A1(net6375),
    .A2(_10772_),
    .B1(net207),
    .Y(_10781_));
 sky130_fd_sc_hd__and3_1 _18943_ (.A(net6375),
    .B(net207),
    .C(_10772_),
    .X(_10782_));
 sky130_fd_sc_hd__o21a_1 _18944_ (.A1(_10781_),
    .A2(_10782_),
    .B1(net2133),
    .X(_10783_));
 sky130_fd_sc_hd__a31o_1 _18945_ (.A1(net9101),
    .A2(net2121),
    .A3(net1450),
    .B1(_10783_),
    .X(_00451_));
 sky130_fd_sc_hd__and3_1 _18946_ (.A(net6375),
    .B(net207),
    .C(_10772_),
    .X(_10784_));
 sky130_fd_sc_hd__nor2_1 _18947_ (.A(net6375),
    .B(net207),
    .Y(_10785_));
 sky130_fd_sc_hd__o21a_1 _18948_ (.A1(_10784_),
    .A2(_10785_),
    .B1(net2133),
    .X(_10786_));
 sky130_fd_sc_hd__a31o_1 _18949_ (.A1(net9073),
    .A2(net2121),
    .A3(net1446),
    .B1(_10786_),
    .X(_00452_));
 sky130_fd_sc_hd__inv_2 _18950_ (.A(net6194),
    .Y(_10787_));
 sky130_fd_sc_hd__nand2_1 _18951_ (.A(net6166),
    .B(net6093),
    .Y(_10788_));
 sky130_fd_sc_hd__nor2_1 _18952_ (.A(net3917),
    .B(_10788_),
    .Y(_10789_));
 sky130_fd_sc_hd__inv_2 _18953_ (.A(net6085),
    .Y(_10790_));
 sky130_fd_sc_hd__nand2_1 _18954_ (.A(net6189),
    .B(net6143),
    .Y(_10791_));
 sky130_fd_sc_hd__xnor2_1 _18955_ (.A(net3910),
    .B(_10791_),
    .Y(_10792_));
 sky130_fd_sc_hd__xnor2_1 _18956_ (.A(net3216),
    .B(net3215),
    .Y(_10793_));
 sky130_fd_sc_hd__nand2_1 _18957_ (.A(net6318),
    .B(net6343),
    .Y(_10794_));
 sky130_fd_sc_hd__or2_2 _18958_ (.A(net6298),
    .B(_10794_),
    .X(_10795_));
 sky130_fd_sc_hd__and2b_2 _18959_ (.A_N(net6248),
    .B(net6231),
    .X(_10796_));
 sky130_fd_sc_hd__xnor2_4 _18960_ (.A(net6209),
    .B(_10796_),
    .Y(_10797_));
 sky130_fd_sc_hd__xnor2_1 _18961_ (.A(net6189),
    .B(net6142),
    .Y(_10798_));
 sky130_fd_sc_hd__xnor2_1 _18962_ (.A(_10797_),
    .B(_10798_),
    .Y(_10799_));
 sky130_fd_sc_hd__inv_2 _18963_ (.A(net6268),
    .Y(_10800_));
 sky130_fd_sc_hd__and2_1 _18964_ (.A(net6222),
    .B(net6241),
    .X(_10801_));
 sky130_fd_sc_hd__or2b_1 _18965_ (.A(net6232),
    .B_N(net6264),
    .X(_10802_));
 sky130_fd_sc_hd__xnor2_1 _18966_ (.A(net6203),
    .B(net6162),
    .Y(_10803_));
 sky130_fd_sc_hd__nor2_1 _18967_ (.A(net6232),
    .B(net6249),
    .Y(_10804_));
 sky130_fd_sc_hd__a221o_1 _18968_ (.A1(_10800_),
    .A2(net3906),
    .B1(_10802_),
    .B2(net3905),
    .C1(_10804_),
    .X(_10805_));
 sky130_fd_sc_hd__or2_1 _18969_ (.A(net2530),
    .B(net3214),
    .X(_10806_));
 sky130_fd_sc_hd__nand2_1 _18970_ (.A(net2530),
    .B(net3214),
    .Y(_10807_));
 sky130_fd_sc_hd__a21boi_2 _18971_ (.A1(_10795_),
    .A2(_10806_),
    .B1_N(_10807_),
    .Y(_10808_));
 sky130_fd_sc_hd__xor2_1 _18972_ (.A(_10793_),
    .B(_10808_),
    .X(_10809_));
 sky130_fd_sc_hd__or2b_1 _18973_ (.A(net6339),
    .B_N(net6318),
    .X(_10810_));
 sky130_fd_sc_hd__clkbuf_2 _18974_ (.A(_10810_),
    .X(_10811_));
 sky130_fd_sc_hd__or2_1 _18975_ (.A(net6270),
    .B(net6290),
    .X(_10812_));
 sky130_fd_sc_hd__and2b_1 _18976_ (.A_N(net6314),
    .B(net6339),
    .X(_10813_));
 sky130_fd_sc_hd__xnor2_1 _18977_ (.A(net6313),
    .B(net6340),
    .Y(_10814_));
 sky130_fd_sc_hd__mux2_1 _18978_ (.A0(net3902),
    .A1(_10814_),
    .S(net6260),
    .X(_10815_));
 sky130_fd_sc_hd__a2bb2o_1 _18979_ (.A1_N(net3213),
    .A2_N(net3903),
    .B1(_10815_),
    .B2(net6291),
    .X(_10816_));
 sky130_fd_sc_hd__nand2_1 _18980_ (.A(net6356),
    .B(net2529),
    .Y(_10817_));
 sky130_fd_sc_hd__xnor2_1 _18981_ (.A(_10795_),
    .B(net3214),
    .Y(_10818_));
 sky130_fd_sc_hd__xnor2_2 _18982_ (.A(net2530),
    .B(_10818_),
    .Y(_10819_));
 sky130_fd_sc_hd__or2b_1 _18983_ (.A(net6352),
    .B_N(net6342),
    .X(_10820_));
 sky130_fd_sc_hd__buf_1 _18984_ (.A(_10820_),
    .X(_10821_));
 sky130_fd_sc_hd__nor2b_1 _18985_ (.A(net6320),
    .B_N(net6289),
    .Y(_10822_));
 sky130_fd_sc_hd__or2b_1 _18986_ (.A(net6312),
    .B_N(net6352),
    .X(_10823_));
 sky130_fd_sc_hd__xor2_1 _18987_ (.A(net6312),
    .B(net6352),
    .X(_10824_));
 sky130_fd_sc_hd__mux2_1 _18988_ (.A0(_10823_),
    .A1(_10824_),
    .S(net6296),
    .X(_10825_));
 sky130_fd_sc_hd__o221ai_1 _18989_ (.A1(_10821_),
    .A2(net3899),
    .B1(_10825_),
    .B2(net6339),
    .C1(net6262),
    .Y(_10826_));
 sky130_fd_sc_hd__inv_2 _18990_ (.A(net6295),
    .Y(_10827_));
 sky130_fd_sc_hd__or2b_1 _18991_ (.A(net6343),
    .B_N(net6357),
    .X(_10828_));
 sky130_fd_sc_hd__clkbuf_2 _18992_ (.A(_10828_),
    .X(_10829_));
 sky130_fd_sc_hd__nand3b_1 _18993_ (.A_N(net6314),
    .B(net6343),
    .C(net6293),
    .Y(_10830_));
 sky130_fd_sc_hd__a21oi_1 _18994_ (.A1(_10811_),
    .A2(_10830_),
    .B1(net6356),
    .Y(_10831_));
 sky130_fd_sc_hd__a311o_1 _18995_ (.A1(_10827_),
    .A2(net3212),
    .A3(_10829_),
    .B1(_10831_),
    .C1(net6266),
    .X(_10832_));
 sky130_fd_sc_hd__nand2_1 _18996_ (.A(net2528),
    .B(_10832_),
    .Y(_10833_));
 sky130_fd_sc_hd__or2b_1 _18997_ (.A(_10819_),
    .B_N(_10833_),
    .X(_10834_));
 sky130_fd_sc_hd__nand2_1 _18998_ (.A(_10817_),
    .B(_10834_),
    .Y(_10835_));
 sky130_fd_sc_hd__buf_1 _18999_ (.A(_10800_),
    .X(_10836_));
 sky130_fd_sc_hd__and2b_1 _19000_ (.A_N(net6342),
    .B(net6351),
    .X(_10837_));
 sky130_fd_sc_hd__nand2_1 _19001_ (.A(net6295),
    .B(net3898),
    .Y(_10838_));
 sky130_fd_sc_hd__nand2_1 _19002_ (.A(net6267),
    .B(net6300),
    .Y(_10839_));
 sky130_fd_sc_hd__nand2_1 _19003_ (.A(net3209),
    .B(_10839_),
    .Y(_10840_));
 sky130_fd_sc_hd__a22o_1 _19004_ (.A1(_10836_),
    .A2(net3211),
    .B1(_10838_),
    .B2(_10840_),
    .X(_10841_));
 sky130_fd_sc_hd__and2b_1 _19005_ (.A_N(net6352),
    .B(net6342),
    .X(_10842_));
 sky130_fd_sc_hd__buf_1 _19006_ (.A(_10842_),
    .X(_10843_));
 sky130_fd_sc_hd__mux2_1 _19007_ (.A0(net3202),
    .A1(net3898),
    .S(_10800_),
    .X(_10844_));
 sky130_fd_sc_hd__a21oi_1 _19008_ (.A1(net6268),
    .A2(_10828_),
    .B1(net3202),
    .Y(_10845_));
 sky130_fd_sc_hd__or2_1 _19009_ (.A(net6292),
    .B(net6313),
    .X(_10846_));
 sky130_fd_sc_hd__nor2_1 _19010_ (.A(_10845_),
    .B(_10846_),
    .Y(_10847_));
 sky130_fd_sc_hd__a221o_1 _19011_ (.A1(net6319),
    .A2(_10841_),
    .B1(_10844_),
    .B2(net6303),
    .C1(_10847_),
    .X(_10848_));
 sky130_fd_sc_hd__xnor2_1 _19012_ (.A(net6114),
    .B(net6155),
    .Y(_10849_));
 sky130_fd_sc_hd__nor2b_2 _19013_ (.A(net6226),
    .B_N(net6205),
    .Y(_10850_));
 sky130_fd_sc_hd__xnor2_4 _19014_ (.A(net6181),
    .B(_10850_),
    .Y(_10851_));
 sky130_fd_sc_hd__xnor2_1 _19015_ (.A(_10849_),
    .B(_10851_),
    .Y(_10852_));
 sky130_fd_sc_hd__or2b_1 _19016_ (.A(net6209),
    .B_N(net6248),
    .X(_10853_));
 sky130_fd_sc_hd__nor2_1 _19017_ (.A(net6209),
    .B(net6234),
    .Y(_10854_));
 sky130_fd_sc_hd__a221o_1 _19018_ (.A1(net6208),
    .A2(_10796_),
    .B1(_10798_),
    .B2(_10853_),
    .C1(_10854_),
    .X(_10855_));
 sky130_fd_sc_hd__and3b_1 _19019_ (.A_N(net6265),
    .B(net6298),
    .C(net6317),
    .X(_10856_));
 sky130_fd_sc_hd__xnor2_1 _19020_ (.A(net6248),
    .B(_10856_),
    .Y(_10857_));
 sky130_fd_sc_hd__xnor2_1 _19021_ (.A(_10855_),
    .B(_10857_),
    .Y(_10858_));
 sky130_fd_sc_hd__xnor2_1 _19022_ (.A(net2527),
    .B(_10858_),
    .Y(_10859_));
 sky130_fd_sc_hd__xnor2_1 _19023_ (.A(net1759),
    .B(_10859_),
    .Y(_10860_));
 sky130_fd_sc_hd__a21o_1 _19024_ (.A1(_10809_),
    .A2(_10835_),
    .B1(_10860_),
    .X(_10861_));
 sky130_fd_sc_hd__o21ai_2 _19025_ (.A1(_10809_),
    .A2(_10835_),
    .B1(_10861_),
    .Y(_10862_));
 sky130_fd_sc_hd__a21o_1 _19026_ (.A1(net2528),
    .A2(_10832_),
    .B1(net3214),
    .X(_10863_));
 sky130_fd_sc_hd__a32o_1 _19027_ (.A1(net3214),
    .A2(net2528),
    .A3(_10832_),
    .B1(_10863_),
    .B2(net2530),
    .X(_10864_));
 sky130_fd_sc_hd__a2111o_1 _19028_ (.A1(net2528),
    .A2(_10832_),
    .B1(_10795_),
    .C1(net2530),
    .D1(net3214),
    .X(_10865_));
 sky130_fd_sc_hd__o221ai_1 _19029_ (.A1(_10817_),
    .A2(_10806_),
    .B1(_10807_),
    .B2(_10833_),
    .C1(_10865_),
    .Y(_10866_));
 sky130_fd_sc_hd__a31o_1 _19030_ (.A1(_10795_),
    .A2(_10864_),
    .A3(_10817_),
    .B1(_10866_),
    .X(_10867_));
 sky130_fd_sc_hd__xnor2_1 _19031_ (.A(_10860_),
    .B(_10793_),
    .Y(_10868_));
 sky130_fd_sc_hd__xnor2_2 _19032_ (.A(_10867_),
    .B(_10868_),
    .Y(_10869_));
 sky130_fd_sc_hd__inv_2 _19033_ (.A(net6105),
    .Y(_10870_));
 sky130_fd_sc_hd__buf_1 _19034_ (.A(_10870_),
    .X(_10871_));
 sky130_fd_sc_hd__a21oi_1 _19035_ (.A1(net6204),
    .A2(net6154),
    .B1(_10871_),
    .Y(_10872_));
 sky130_fd_sc_hd__and3_1 _19036_ (.A(net6204),
    .B(net6154),
    .C(_10870_),
    .X(_10873_));
 sky130_fd_sc_hd__o2111a_1 _19037_ (.A1(_10872_),
    .A2(_10873_),
    .B1(net6178),
    .C1(net6220),
    .D1(net6115),
    .X(_10874_));
 sky130_fd_sc_hd__and2b_1 _19038_ (.A_N(net6260),
    .B(net6245),
    .X(_10875_));
 sky130_fd_sc_hd__xnor2_2 _19039_ (.A(net6229),
    .B(_10875_),
    .Y(_10876_));
 sky130_fd_sc_hd__xnor2_1 _19040_ (.A(_10876_),
    .B(net3904),
    .Y(_10877_));
 sky130_fd_sc_hd__nor2b_1 _19041_ (.A(net6298),
    .B_N(net6266),
    .Y(_10878_));
 sky130_fd_sc_hd__inv_2 _19042_ (.A(net6252),
    .Y(_10879_));
 sky130_fd_sc_hd__xor2_2 _19043_ (.A(net6187),
    .B(net6229),
    .X(_10880_));
 sky130_fd_sc_hd__a21oi_1 _19044_ (.A1(net6296),
    .A2(net3891),
    .B1(_10880_),
    .Y(_10881_));
 sky130_fd_sc_hd__nor2_1 _19045_ (.A(net6261),
    .B(net6245),
    .Y(_10882_));
 sky130_fd_sc_hd__a211o_1 _19046_ (.A1(net6245),
    .A2(net3896),
    .B1(_10881_),
    .C1(_10882_),
    .X(_10883_));
 sky130_fd_sc_hd__or2_1 _19047_ (.A(_10877_),
    .B(_10883_),
    .X(_10884_));
 sky130_fd_sc_hd__nand2_1 _19048_ (.A(net6356),
    .B(_10813_),
    .Y(_10885_));
 sky130_fd_sc_hd__a21o_1 _19049_ (.A1(_10877_),
    .A2(_10883_),
    .B1(_10885_),
    .X(_10886_));
 sky130_fd_sc_hd__a311o_1 _19050_ (.A1(net6178),
    .A2(net6220),
    .A3(net6120),
    .B1(_10872_),
    .C1(_10873_),
    .X(_10887_));
 sky130_fd_sc_hd__a21boi_1 _19051_ (.A1(_10884_),
    .A2(_10886_),
    .B1_N(net2113),
    .Y(_10888_));
 sky130_fd_sc_hd__nor2_1 _19052_ (.A(net2117),
    .B(_10888_),
    .Y(_10889_));
 sky130_fd_sc_hd__and2b_1 _19053_ (.A_N(net2117),
    .B(net2113),
    .X(_10890_));
 sky130_fd_sc_hd__a21oi_1 _19054_ (.A1(_10884_),
    .A2(_10886_),
    .B1(_10890_),
    .Y(_10891_));
 sky130_fd_sc_hd__and3_1 _19055_ (.A(_10884_),
    .B(_10886_),
    .C(_10890_),
    .X(_10892_));
 sky130_fd_sc_hd__or2_1 _19056_ (.A(_10891_),
    .B(_10892_),
    .X(_10893_));
 sky130_fd_sc_hd__o21ai_1 _19057_ (.A1(net6314),
    .A2(_10829_),
    .B1(net3211),
    .Y(_10894_));
 sky130_fd_sc_hd__o221a_1 _19058_ (.A1(net6360),
    .A2(_10811_),
    .B1(_10894_),
    .B2(net6293),
    .C1(_10830_),
    .X(_10895_));
 sky130_fd_sc_hd__xnor2_1 _19059_ (.A(net3208),
    .B(_10895_),
    .Y(_10896_));
 sky130_fd_sc_hd__xnor2_2 _19060_ (.A(_10819_),
    .B(_10896_),
    .Y(_10897_));
 sky130_fd_sc_hd__inv_2 _19061_ (.A(net6352),
    .Y(_10898_));
 sky130_fd_sc_hd__xnor2_2 _19062_ (.A(_10827_),
    .B(_10811_),
    .Y(_10899_));
 sky130_fd_sc_hd__nor2_1 _19063_ (.A(_10898_),
    .B(net2525),
    .Y(_10900_));
 sky130_fd_sc_hd__and2_1 _19064_ (.A(_10898_),
    .B(net2525),
    .X(_10901_));
 sky130_fd_sc_hd__nor2_1 _19065_ (.A(_10900_),
    .B(_10901_),
    .Y(_10902_));
 sky130_fd_sc_hd__xor2_1 _19066_ (.A(_10877_),
    .B(_10883_),
    .X(_10903_));
 sky130_fd_sc_hd__xnor2_1 _19067_ (.A(_10885_),
    .B(_10903_),
    .Y(_10904_));
 sky130_fd_sc_hd__o311a_1 _19068_ (.A1(_10891_),
    .A2(_10892_),
    .A3(_10897_),
    .B1(net1758),
    .C1(_10904_),
    .X(_10905_));
 sky130_fd_sc_hd__a21oi_1 _19069_ (.A1(_10893_),
    .A2(_10897_),
    .B1(_10905_),
    .Y(_10906_));
 sky130_fd_sc_hd__a21o_1 _19070_ (.A1(_10869_),
    .A2(_10889_),
    .B1(_10906_),
    .X(_10907_));
 sky130_fd_sc_hd__or2_1 _19071_ (.A(_10869_),
    .B(_10889_),
    .X(_10908_));
 sky130_fd_sc_hd__and3_1 _19072_ (.A(_10862_),
    .B(_10907_),
    .C(_10908_),
    .X(_10909_));
 sky130_fd_sc_hd__or2_1 _19073_ (.A(net2527),
    .B(_10855_),
    .X(_10910_));
 sky130_fd_sc_hd__buf_1 _19074_ (.A(_10827_),
    .X(_10911_));
 sky130_fd_sc_hd__or2_1 _19075_ (.A(net6260),
    .B(net6311),
    .X(_10912_));
 sky130_fd_sc_hd__nor2_1 _19076_ (.A(net3211),
    .B(_10912_),
    .Y(_10913_));
 sky130_fd_sc_hd__a211oi_1 _19077_ (.A1(net6319),
    .A2(_10845_),
    .B1(_10913_),
    .C1(net6249),
    .Y(_10914_));
 sky130_fd_sc_hd__o221a_1 _19078_ (.A1(net6357),
    .A2(net3908),
    .B1(_10829_),
    .B2(_10912_),
    .C1(net6249),
    .X(_10915_));
 sky130_fd_sc_hd__nand2_1 _19079_ (.A(net6268),
    .B(_10911_),
    .Y(_10916_));
 sky130_fd_sc_hd__or2_1 _19080_ (.A(net6247),
    .B(net6328),
    .X(_10917_));
 sky130_fd_sc_hd__nand2_1 _19081_ (.A(net6247),
    .B(net6321),
    .Y(_10918_));
 sky130_fd_sc_hd__nand2_1 _19082_ (.A(_10917_),
    .B(_10918_),
    .Y(_10919_));
 sky130_fd_sc_hd__mux2_1 _19083_ (.A0(net3211),
    .A1(_10829_),
    .S(net3192),
    .X(_10920_));
 sky130_fd_sc_hd__o32a_1 _19084_ (.A1(_10911_),
    .A2(_10914_),
    .A3(_10915_),
    .B1(_10916_),
    .B2(_10920_),
    .X(_10921_));
 sky130_fd_sc_hd__nor2_1 _19085_ (.A(_10910_),
    .B(net1757),
    .Y(_10922_));
 sky130_fd_sc_hd__nand2_1 _19086_ (.A(net3894),
    .B(net6321),
    .Y(_10923_));
 sky130_fd_sc_hd__a21o_1 _19087_ (.A1(net3892),
    .A2(_10829_),
    .B1(net6268),
    .X(_10924_));
 sky130_fd_sc_hd__a21o_1 _19088_ (.A1(net3191),
    .A2(_10924_),
    .B1(_10911_),
    .X(_10925_));
 sky130_fd_sc_hd__o21ai_1 _19089_ (.A1(net3896),
    .A2(net3192),
    .B1(net3202),
    .Y(_10926_));
 sky130_fd_sc_hd__a21o_1 _19090_ (.A1(_10827_),
    .A2(net6318),
    .B1(net3898),
    .X(_10927_));
 sky130_fd_sc_hd__a21oi_1 _19091_ (.A1(net3209),
    .A2(_10917_),
    .B1(net6300),
    .Y(_10928_));
 sky130_fd_sc_hd__a21oi_1 _19092_ (.A1(net6246),
    .A2(_10927_),
    .B1(_10928_),
    .Y(_10929_));
 sky130_fd_sc_hd__nand2_1 _19093_ (.A(net6292),
    .B(net6244),
    .Y(_10930_));
 sky130_fd_sc_hd__o22a_1 _19094_ (.A1(net6268),
    .A2(net3192),
    .B1(net3885),
    .B2(net6319),
    .X(_10931_));
 sky130_fd_sc_hd__o22a_1 _19095_ (.A1(net3208),
    .A2(_10929_),
    .B1(_10931_),
    .B2(net3202),
    .X(_10932_));
 sky130_fd_sc_hd__and2_1 _19096_ (.A(net2527),
    .B(_10855_),
    .X(_10933_));
 sky130_fd_sc_hd__a41oi_2 _19097_ (.A1(_10925_),
    .A2(_10926_),
    .A3(net1756),
    .A4(_10910_),
    .B1(_10933_),
    .Y(_10934_));
 sky130_fd_sc_hd__or2b_1 _19098_ (.A(_10934_),
    .B_N(net1757),
    .X(_10935_));
 sky130_fd_sc_hd__or2b_1 _19099_ (.A(_10922_),
    .B_N(_10935_),
    .X(_10936_));
 sky130_fd_sc_hd__and2b_1 _19100_ (.A_N(net6204),
    .B(net6178),
    .X(_10937_));
 sky130_fd_sc_hd__xnor2_2 _19101_ (.A(net6162),
    .B(_10937_),
    .Y(_10938_));
 sky130_fd_sc_hd__xnor2_2 _19102_ (.A(net6147),
    .B(net6101),
    .Y(_10939_));
 sky130_fd_sc_hd__xnor2_2 _19103_ (.A(net3190),
    .B(_10939_),
    .Y(_10940_));
 sky130_fd_sc_hd__nand2_1 _19104_ (.A(net6340),
    .B(net6353),
    .Y(_10941_));
 sky130_fd_sc_hd__a21o_1 _19105_ (.A1(net6243),
    .A2(_10941_),
    .B1(net3889),
    .X(_10942_));
 sky130_fd_sc_hd__and2_1 _19106_ (.A(net6336),
    .B(net6359),
    .X(_10943_));
 sky130_fd_sc_hd__nand2_1 _19107_ (.A(net6272),
    .B(net6241),
    .Y(_10944_));
 sky130_fd_sc_hd__a21oi_1 _19108_ (.A1(_10943_),
    .A2(_10944_),
    .B1(net6302),
    .Y(_10945_));
 sky130_fd_sc_hd__inv_2 _19109_ (.A(net6226),
    .Y(_10946_));
 sky130_fd_sc_hd__o2bb2a_1 _19110_ (.A1_N(_10946_),
    .A2_N(_10849_),
    .B1(net6181),
    .B2(net6205),
    .X(_10947_));
 sky130_fd_sc_hd__o21ai_1 _19111_ (.A1(_10849_),
    .A2(_10850_),
    .B1(net6182),
    .Y(_10948_));
 sky130_fd_sc_hd__o211ai_1 _19112_ (.A1(net3189),
    .A2(_10945_),
    .B1(_10947_),
    .C1(_10948_),
    .Y(_10949_));
 sky130_fd_sc_hd__a211o_1 _19113_ (.A1(_10947_),
    .A2(_10948_),
    .B1(net3189),
    .C1(_10945_),
    .X(_10950_));
 sky130_fd_sc_hd__nand3_1 _19114_ (.A(_10940_),
    .B(_10949_),
    .C(_10950_),
    .Y(_10951_));
 sky130_fd_sc_hd__a21o_1 _19115_ (.A1(_10949_),
    .A2(_10950_),
    .B1(_10940_),
    .X(_10952_));
 sky130_fd_sc_hd__xnor2_1 _19116_ (.A(_10876_),
    .B(_10899_),
    .Y(_10953_));
 sky130_fd_sc_hd__o21a_1 _19117_ (.A1(net6311),
    .A2(net3212),
    .B1(_10811_),
    .X(_10954_));
 sky130_fd_sc_hd__xnor2_2 _19118_ (.A(net6245),
    .B(net3896),
    .Y(_10955_));
 sky130_fd_sc_hd__mux2_1 _19119_ (.A0(_10954_),
    .A1(_10885_),
    .S(_10955_),
    .X(_10956_));
 sky130_fd_sc_hd__xnor2_1 _19120_ (.A(net2110),
    .B(net2109),
    .Y(_10957_));
 sky130_fd_sc_hd__nand3_1 _19121_ (.A(net2112),
    .B(net2111),
    .C(_10957_),
    .Y(_10958_));
 sky130_fd_sc_hd__a21o_1 _19122_ (.A1(net2112),
    .A2(net2111),
    .B1(_10957_),
    .X(_10959_));
 sky130_fd_sc_hd__nand2_1 _19123_ (.A(_10958_),
    .B(_10959_),
    .Y(_10960_));
 sky130_fd_sc_hd__nand2_1 _19124_ (.A(net6119),
    .B(net6155),
    .Y(_10961_));
 sky130_fd_sc_hd__xnor2_1 _19125_ (.A(net6069),
    .B(_10961_),
    .Y(_10962_));
 sky130_fd_sc_hd__nor2_1 _19126_ (.A(net3910),
    .B(_10791_),
    .Y(_10963_));
 sky130_fd_sc_hd__xor2_1 _19127_ (.A(net3187),
    .B(_10963_),
    .X(_10964_));
 sky130_fd_sc_hd__xnor2_1 _19128_ (.A(_10960_),
    .B(_10964_),
    .Y(_10965_));
 sky130_fd_sc_hd__xnor2_2 _19129_ (.A(_10936_),
    .B(_10965_),
    .Y(_10966_));
 sky130_fd_sc_hd__a21bo_1 _19130_ (.A1(net3216),
    .A2(_10808_),
    .B1_N(net3215),
    .X(_10967_));
 sky130_fd_sc_hd__o21ai_1 _19131_ (.A1(net3216),
    .A2(_10808_),
    .B1(_10967_),
    .Y(_10968_));
 sky130_fd_sc_hd__o211a_1 _19132_ (.A1(_10862_),
    .A2(_10966_),
    .B1(_10908_),
    .C1(_10907_),
    .X(_10969_));
 sky130_fd_sc_hd__a21o_1 _19133_ (.A1(_10862_),
    .A2(_10966_),
    .B1(_10969_),
    .X(_10970_));
 sky130_fd_sc_hd__xor2_2 _19134_ (.A(net6119),
    .B(net6086),
    .X(_10971_));
 sky130_fd_sc_hd__and2b_1 _19135_ (.A_N(net6175),
    .B(net6151),
    .X(_10972_));
 sky130_fd_sc_hd__xnor2_1 _19136_ (.A(net6130),
    .B(_10972_),
    .Y(_10973_));
 sky130_fd_sc_hd__xor2_2 _19137_ (.A(_10971_),
    .B(net3185),
    .X(_10974_));
 sky130_fd_sc_hd__nand2_1 _19138_ (.A(net6184),
    .B(net6153),
    .Y(_10975_));
 sky130_fd_sc_hd__or2b_1 _19139_ (.A(_10939_),
    .B_N(_10975_),
    .X(_10976_));
 sky130_fd_sc_hd__nor2_1 _19140_ (.A(net6180),
    .B(net6158),
    .Y(_10977_));
 sky130_fd_sc_hd__a221oi_1 _19141_ (.A1(net6153),
    .A2(_10939_),
    .B1(_10976_),
    .B2(net3915),
    .C1(_10977_),
    .Y(_10978_));
 sky130_fd_sc_hd__or2_1 _19142_ (.A(net3908),
    .B(net3906),
    .X(_10979_));
 sky130_fd_sc_hd__a221o_1 _19143_ (.A1(net6232),
    .A2(net3908),
    .B1(_10979_),
    .B2(net3206),
    .C1(_10804_),
    .X(_10980_));
 sky130_fd_sc_hd__xnor2_1 _19144_ (.A(net2522),
    .B(net2521),
    .Y(_10981_));
 sky130_fd_sc_hd__xnor2_2 _19145_ (.A(_10974_),
    .B(_10981_),
    .Y(_10982_));
 sky130_fd_sc_hd__nand2_2 _19146_ (.A(net6299),
    .B(net6327),
    .Y(_10983_));
 sky130_fd_sc_hd__xnor2_2 _19147_ (.A(_10983_),
    .B(_10797_),
    .Y(_10984_));
 sky130_fd_sc_hd__and2b_1 _19148_ (.A_N(net6267),
    .B(net6300),
    .X(_10985_));
 sky130_fd_sc_hd__nor2_2 _19149_ (.A(net3895),
    .B(_10985_),
    .Y(_10986_));
 sky130_fd_sc_hd__xnor2_1 _19150_ (.A(net6355),
    .B(_10986_),
    .Y(_10987_));
 sky130_fd_sc_hd__xnor2_1 _19151_ (.A(_10984_),
    .B(_10987_),
    .Y(_10988_));
 sky130_fd_sc_hd__nor2_1 _19152_ (.A(net6290),
    .B(net6334),
    .Y(_10989_));
 sky130_fd_sc_hd__a21o_1 _19153_ (.A1(net6323),
    .A2(_10989_),
    .B1(net3901),
    .X(_10990_));
 sky130_fd_sc_hd__nor2_1 _19154_ (.A(net6295),
    .B(net3909),
    .Y(_10991_));
 sky130_fd_sc_hd__mux2_1 _19155_ (.A0(net3184),
    .A1(_10991_),
    .S(_10876_),
    .X(_10992_));
 sky130_fd_sc_hd__xor2_1 _19156_ (.A(_10988_),
    .B(net2520),
    .X(_10993_));
 sky130_fd_sc_hd__xnor2_2 _19157_ (.A(_10982_),
    .B(_10993_),
    .Y(_10994_));
 sky130_fd_sc_hd__inv_2 _19158_ (.A(net6069),
    .Y(_10995_));
 sky130_fd_sc_hd__inv_2 _19159_ (.A(net6049),
    .Y(_10996_));
 sky130_fd_sc_hd__a21oi_1 _19160_ (.A1(net6138),
    .A2(net6101),
    .B1(net3878),
    .Y(_10997_));
 sky130_fd_sc_hd__and3_1 _19161_ (.A(net6147),
    .B(net6101),
    .C(net3878),
    .X(_10998_));
 sky130_fd_sc_hd__nor2_1 _19162_ (.A(_10997_),
    .B(_10998_),
    .Y(_10999_));
 sky130_fd_sc_hd__or3_1 _19163_ (.A(_10995_),
    .B(_10961_),
    .C(_10999_),
    .X(_11000_));
 sky130_fd_sc_hd__a311o_1 _19164_ (.A1(net6119),
    .A2(net6155),
    .A3(net6069),
    .B1(_10997_),
    .C1(_10998_),
    .X(_11001_));
 sky130_fd_sc_hd__nand2_1 _19165_ (.A(_11000_),
    .B(_11001_),
    .Y(_11002_));
 sky130_fd_sc_hd__or2_1 _19166_ (.A(net3189),
    .B(_10945_),
    .X(_11003_));
 sky130_fd_sc_hd__nand2_1 _19167_ (.A(_10947_),
    .B(_10948_),
    .Y(_11004_));
 sky130_fd_sc_hd__a21o_1 _19168_ (.A1(_10940_),
    .A2(_11003_),
    .B1(_11004_),
    .X(_11005_));
 sky130_fd_sc_hd__o21a_1 _19169_ (.A1(_10940_),
    .A2(_11003_),
    .B1(_11005_),
    .X(_11006_));
 sky130_fd_sc_hd__xnor2_1 _19170_ (.A(_11002_),
    .B(_11006_),
    .Y(_11007_));
 sky130_fd_sc_hd__o2bb2a_1 _19171_ (.A1_N(net2112),
    .A2_N(net2111),
    .B1(net2110),
    .B2(net2109),
    .X(_11008_));
 sky130_fd_sc_hd__a21o_1 _19172_ (.A1(net2110),
    .A2(net2109),
    .B1(_11008_),
    .X(_11009_));
 sky130_fd_sc_hd__xor2_1 _19173_ (.A(net1426),
    .B(_11009_),
    .X(_11010_));
 sky130_fd_sc_hd__xnor2_1 _19174_ (.A(_10994_),
    .B(_11010_),
    .Y(_11011_));
 sky130_fd_sc_hd__inv_2 _19175_ (.A(_10963_),
    .Y(_11012_));
 sky130_fd_sc_hd__nand3_1 _19176_ (.A(_11012_),
    .B(_10958_),
    .C(_10959_),
    .Y(_11013_));
 sky130_fd_sc_hd__inv_2 _19177_ (.A(net3187),
    .Y(_11014_));
 sky130_fd_sc_hd__a21oi_1 _19178_ (.A1(_11014_),
    .A2(_10910_),
    .B1(net1757),
    .Y(_11015_));
 sky130_fd_sc_hd__a21o_1 _19179_ (.A1(net3187),
    .A2(_10934_),
    .B1(_11015_),
    .X(_11016_));
 sky130_fd_sc_hd__a21oi_1 _19180_ (.A1(_10958_),
    .A2(_10959_),
    .B1(_11012_),
    .Y(_11017_));
 sky130_fd_sc_hd__a32o_1 _19181_ (.A1(net3187),
    .A2(_10922_),
    .A3(_11013_),
    .B1(_11016_),
    .B2(_11017_),
    .X(_11018_));
 sky130_fd_sc_hd__or2_1 _19182_ (.A(_11016_),
    .B(_11013_),
    .X(_11019_));
 sky130_fd_sc_hd__or3_1 _19183_ (.A(net3187),
    .B(_11017_),
    .C(_10935_),
    .X(_11020_));
 sky130_fd_sc_hd__and3b_1 _19184_ (.A_N(_11018_),
    .B(_11019_),
    .C(_11020_),
    .X(_11021_));
 sky130_fd_sc_hd__xnor2_1 _19185_ (.A(net1064),
    .B(_11021_),
    .Y(_11022_));
 sky130_fd_sc_hd__a221o_1 _19186_ (.A1(_10909_),
    .A2(_10966_),
    .B1(_10968_),
    .B2(_10970_),
    .C1(net872),
    .X(_11023_));
 sky130_fd_sc_hd__or2b_1 _19187_ (.A(net6259),
    .B_N(net6315),
    .X(_11024_));
 sky130_fd_sc_hd__xnor2_1 _19188_ (.A(net6201),
    .B(net6240),
    .Y(_11025_));
 sky130_fd_sc_hd__nor2_1 _19189_ (.A(net6259),
    .B(net6294),
    .Y(_11026_));
 sky130_fd_sc_hd__a221o_1 _19190_ (.A1(net6259),
    .A2(net3900),
    .B1(_11024_),
    .B2(net3877),
    .C1(_11026_),
    .X(_11027_));
 sky130_fd_sc_hd__xor2_2 _19191_ (.A(_10955_),
    .B(_10880_),
    .X(_11028_));
 sky130_fd_sc_hd__xnor2_1 _19192_ (.A(net6312),
    .B(_10843_),
    .Y(_11029_));
 sky130_fd_sc_hd__a21o_1 _19193_ (.A1(net3183),
    .A2(_11028_),
    .B1(_11029_),
    .X(_11030_));
 sky130_fd_sc_hd__nor2_1 _19194_ (.A(_10898_),
    .B(_10813_),
    .Y(_11031_));
 sky130_fd_sc_hd__xnor2_1 _19195_ (.A(_10899_),
    .B(_11031_),
    .Y(_11032_));
 sky130_fd_sc_hd__xnor2_1 _19196_ (.A(_10903_),
    .B(_11032_),
    .Y(_11033_));
 sky130_fd_sc_hd__or2_1 _19197_ (.A(net3183),
    .B(_11028_),
    .X(_11034_));
 sky130_fd_sc_hd__inv_2 _19198_ (.A(net6115),
    .Y(_11035_));
 sky130_fd_sc_hd__nand2_1 _19199_ (.A(net6179),
    .B(net6227),
    .Y(_11036_));
 sky130_fd_sc_hd__xnor2_1 _19200_ (.A(net3876),
    .B(_11036_),
    .Y(_11037_));
 sky130_fd_sc_hd__and3_1 _19201_ (.A(net6207),
    .B(net6141),
    .C(net6244),
    .X(_11038_));
 sky130_fd_sc_hd__xnor2_1 _19202_ (.A(net3180),
    .B(_11038_),
    .Y(_11039_));
 sky130_fd_sc_hd__nand2_1 _19203_ (.A(_11034_),
    .B(_11039_),
    .Y(_11040_));
 sky130_fd_sc_hd__and2_1 _19204_ (.A(net3183),
    .B(_11029_),
    .X(_11041_));
 sky130_fd_sc_hd__nor2_1 _19205_ (.A(net3183),
    .B(_11029_),
    .Y(_11042_));
 sky130_fd_sc_hd__o21ba_1 _19206_ (.A1(_11028_),
    .A2(_11041_),
    .B1_N(_11042_),
    .X(_11043_));
 sky130_fd_sc_hd__or3_1 _19207_ (.A(_11043_),
    .B(_11033_),
    .C(_11039_),
    .X(_11044_));
 sky130_fd_sc_hd__a22o_1 _19208_ (.A1(_11030_),
    .A2(_11033_),
    .B1(_11040_),
    .B2(_11044_),
    .X(_11045_));
 sky130_fd_sc_hd__inv_2 _19209_ (.A(net6152),
    .Y(_11046_));
 sky130_fd_sc_hd__nand2_1 _19210_ (.A(net6276),
    .B(net6218),
    .Y(_11047_));
 sky130_fd_sc_hd__nor2_2 _19211_ (.A(_11046_),
    .B(_11047_),
    .Y(_11048_));
 sky130_fd_sc_hd__and2_1 _19212_ (.A(net6258),
    .B(net6313),
    .X(_11049_));
 sky130_fd_sc_hd__or2b_1 _19213_ (.A(net6335),
    .B_N(net6287),
    .X(_11050_));
 sky130_fd_sc_hd__and2b_1 _19214_ (.A_N(net6287),
    .B(net6337),
    .X(_11051_));
 sky130_fd_sc_hd__a21o_1 _19215_ (.A1(net3883),
    .A2(_11050_),
    .B1(_11051_),
    .X(_11052_));
 sky130_fd_sc_hd__a32o_1 _19216_ (.A1(net3205),
    .A2(net6225),
    .A3(net3901),
    .B1(_11049_),
    .B2(_11052_),
    .X(_11053_));
 sky130_fd_sc_hd__xor2_2 _19217_ (.A(net6271),
    .B(net6224),
    .X(_11054_));
 sky130_fd_sc_hd__o221a_1 _19218_ (.A1(net6340),
    .A2(net3882),
    .B1(_11051_),
    .B2(net3874),
    .C1(_10846_),
    .X(_11055_));
 sky130_fd_sc_hd__xnor2_2 _19219_ (.A(net6271),
    .B(_10822_),
    .Y(_11056_));
 sky130_fd_sc_hd__a21o_1 _19220_ (.A1(net3178),
    .A2(_11056_),
    .B1(net3890),
    .X(_11057_));
 sky130_fd_sc_hd__o21a_1 _19221_ (.A1(net6240),
    .A2(net2519),
    .B1(_11057_),
    .X(_11058_));
 sky130_fd_sc_hd__a21o_1 _19222_ (.A1(_11048_),
    .A2(_11057_),
    .B1(net6139),
    .X(_11059_));
 sky130_fd_sc_hd__o21a_1 _19223_ (.A1(_11048_),
    .A2(_11058_),
    .B1(_11059_),
    .X(_11060_));
 sky130_fd_sc_hd__clkbuf_1 _19224_ (.A(net3890),
    .X(_11061_));
 sky130_fd_sc_hd__a21o_1 _19225_ (.A1(net2519),
    .A2(_11048_),
    .B1(net3175),
    .X(_11062_));
 sky130_fd_sc_hd__a21o_1 _19226_ (.A1(net3178),
    .A2(_11056_),
    .B1(_11048_),
    .X(_11063_));
 sky130_fd_sc_hd__nor2_1 _19227_ (.A(net6139),
    .B(net3175),
    .Y(_11064_));
 sky130_fd_sc_hd__a311o_1 _19228_ (.A1(net6139),
    .A2(_11062_),
    .A3(_11063_),
    .B1(_11064_),
    .C1(net3918),
    .X(_11065_));
 sky130_fd_sc_hd__a211o_1 _19229_ (.A1(net6240),
    .A2(_11048_),
    .B1(net2519),
    .C1(net6139),
    .X(_11066_));
 sky130_fd_sc_hd__o211a_1 _19230_ (.A1(net6201),
    .A2(_11060_),
    .B1(_11065_),
    .C1(_11066_),
    .X(_11067_));
 sky130_fd_sc_hd__xnor2_1 _19231_ (.A(_11043_),
    .B(_11039_),
    .Y(_11068_));
 sky130_fd_sc_hd__xnor2_1 _19232_ (.A(_11033_),
    .B(_11068_),
    .Y(_11069_));
 sky130_fd_sc_hd__nor2_1 _19233_ (.A(net1422),
    .B(_11069_),
    .Y(_11070_));
 sky130_fd_sc_hd__o21ba_1 _19234_ (.A1(net6230),
    .A2(net6340),
    .B1_N(_11024_),
    .X(_11071_));
 sky130_fd_sc_hd__or2b_1 _19235_ (.A(net6336),
    .B_N(net6225),
    .X(_11072_));
 sky130_fd_sc_hd__a21oi_1 _19236_ (.A1(net6321),
    .A2(_11072_),
    .B1(net3206),
    .Y(_11073_));
 sky130_fd_sc_hd__o21a_1 _19237_ (.A1(_11071_),
    .A2(_11073_),
    .B1(net3198),
    .X(_11074_));
 sky130_fd_sc_hd__or2b_1 _19238_ (.A(net6323),
    .B_N(net6221),
    .X(_11075_));
 sky130_fd_sc_hd__or2b_1 _19239_ (.A(net6222),
    .B_N(net6323),
    .X(_11076_));
 sky130_fd_sc_hd__a21o_1 _19240_ (.A1(_11076_),
    .A2(_11072_),
    .B1(net6273),
    .X(_11077_));
 sky130_fd_sc_hd__and3_1 _19241_ (.A(net6288),
    .B(_11075_),
    .C(_11077_),
    .X(_11078_));
 sky130_fd_sc_hd__o22a_1 _19242_ (.A1(net3908),
    .A2(_10802_),
    .B1(_11074_),
    .B2(_11078_),
    .X(_11079_));
 sky130_fd_sc_hd__xor2_1 _19243_ (.A(net3877),
    .B(_11079_),
    .X(_11080_));
 sky130_fd_sc_hd__a21oi_1 _19244_ (.A1(_10821_),
    .A2(net3210),
    .B1(_11080_),
    .Y(_11081_));
 sky130_fd_sc_hd__mux2_1 _19245_ (.A0(net6240),
    .A1(_11056_),
    .S(net3178),
    .X(_11082_));
 sky130_fd_sc_hd__nor2_1 _19246_ (.A(net6201),
    .B(net6240),
    .Y(_11083_));
 sky130_fd_sc_hd__mux2_1 _19247_ (.A0(_11083_),
    .A1(net6240),
    .S(_11056_),
    .X(_11084_));
 sky130_fd_sc_hd__a22o_1 _19248_ (.A1(net6201),
    .A2(_11082_),
    .B1(_11084_),
    .B2(net3178),
    .X(_11085_));
 sky130_fd_sc_hd__xnor2_1 _19249_ (.A(net6129),
    .B(_11048_),
    .Y(_11086_));
 sky130_fd_sc_hd__xnor2_1 _19250_ (.A(_11085_),
    .B(_11086_),
    .Y(_11087_));
 sky130_fd_sc_hd__nor2_1 _19251_ (.A(_11042_),
    .B(_11041_),
    .Y(_11088_));
 sky130_fd_sc_hd__xnor2_1 _19252_ (.A(_11028_),
    .B(_11088_),
    .Y(_11089_));
 sky130_fd_sc_hd__or2_1 _19253_ (.A(net1753),
    .B(_11089_),
    .X(_11090_));
 sky130_fd_sc_hd__and2_1 _19254_ (.A(net1753),
    .B(_11089_),
    .X(_11091_));
 sky130_fd_sc_hd__a21oi_1 _19255_ (.A1(net1193),
    .A2(_11090_),
    .B1(_11091_),
    .Y(_11092_));
 sky130_fd_sc_hd__nand2_1 _19256_ (.A(net1422),
    .B(_11069_),
    .Y(_11093_));
 sky130_fd_sc_hd__o21a_1 _19257_ (.A1(_11070_),
    .A2(_11092_),
    .B1(_11093_),
    .X(_11094_));
 sky130_fd_sc_hd__xor2_1 _19258_ (.A(_10906_),
    .B(_10889_),
    .X(_11095_));
 sky130_fd_sc_hd__xnor2_2 _19259_ (.A(_10869_),
    .B(_11095_),
    .Y(_11096_));
 sky130_fd_sc_hd__or3b_1 _19260_ (.A(_11045_),
    .B(_11094_),
    .C_N(_11096_),
    .X(_11097_));
 sky130_fd_sc_hd__o21ba_1 _19261_ (.A1(_11034_),
    .A2(net3180),
    .B1_N(_11038_),
    .X(_11098_));
 sky130_fd_sc_hd__a21o_1 _19262_ (.A1(_11034_),
    .A2(net3180),
    .B1(_11098_),
    .X(_11099_));
 sky130_fd_sc_hd__nand2_1 _19263_ (.A(_10904_),
    .B(net1758),
    .Y(_11100_));
 sky130_fd_sc_hd__xnor2_1 _19264_ (.A(_11100_),
    .B(_10893_),
    .Y(_11101_));
 sky130_fd_sc_hd__xnor2_1 _19265_ (.A(_10897_),
    .B(_11101_),
    .Y(_11102_));
 sky130_fd_sc_hd__nor2_1 _19266_ (.A(_11099_),
    .B(_11102_),
    .Y(_11103_));
 sky130_fd_sc_hd__a21oi_1 _19267_ (.A1(_11099_),
    .A2(_11102_),
    .B1(_11045_),
    .Y(_11104_));
 sky130_fd_sc_hd__o21ai_1 _19268_ (.A1(_11103_),
    .A2(_11104_),
    .B1(_11096_),
    .Y(_11105_));
 sky130_fd_sc_hd__nand2_1 _19269_ (.A(_11097_),
    .B(_11105_),
    .Y(_11106_));
 sky130_fd_sc_hd__nand2_1 _19270_ (.A(_11099_),
    .B(_11102_),
    .Y(_11107_));
 sky130_fd_sc_hd__and3b_1 _19271_ (.A_N(_11094_),
    .B(_11096_),
    .C(_11107_),
    .X(_11108_));
 sky130_fd_sc_hd__and2_1 _19272_ (.A(_10966_),
    .B(_10968_),
    .X(_11109_));
 sky130_fd_sc_hd__nor2_1 _19273_ (.A(_10966_),
    .B(_10968_),
    .Y(_11110_));
 sky130_fd_sc_hd__nor2_1 _19274_ (.A(_11109_),
    .B(_11110_),
    .Y(_11111_));
 sky130_fd_sc_hd__a21oi_1 _19275_ (.A1(_10907_),
    .A2(_10908_),
    .B1(_10862_),
    .Y(_11112_));
 sky130_fd_sc_hd__mux2_1 _19276_ (.A0(_10909_),
    .A1(_11112_),
    .S(net872),
    .X(_11113_));
 sky130_fd_sc_hd__nand2_1 _19277_ (.A(_10907_),
    .B(_10908_),
    .Y(_11114_));
 sky130_fd_sc_hd__xnor2_1 _19278_ (.A(_10862_),
    .B(_11114_),
    .Y(_11115_));
 sky130_fd_sc_hd__mux2_1 _19279_ (.A0(_11109_),
    .A1(_11110_),
    .S(net872),
    .X(_11116_));
 sky130_fd_sc_hd__a22o_1 _19280_ (.A1(_11111_),
    .A2(_11113_),
    .B1(_11115_),
    .B2(_11116_),
    .X(_11117_));
 sky130_fd_sc_hd__o21ai_1 _19281_ (.A1(_11106_),
    .A2(_11108_),
    .B1(net763),
    .Y(_11118_));
 sky130_fd_sc_hd__a21o_1 _19282_ (.A1(net6294),
    .A2(net3213),
    .B1(net3902),
    .X(_11119_));
 sky130_fd_sc_hd__or2b_1 _19283_ (.A(net6323),
    .B_N(net6335),
    .X(_11120_));
 sky130_fd_sc_hd__a21o_1 _19284_ (.A1(net6290),
    .A2(_11120_),
    .B1(_11049_),
    .X(_11121_));
 sky130_fd_sc_hd__buf_1 _19285_ (.A(net3886),
    .X(_11122_));
 sky130_fd_sc_hd__a22o_1 _19286_ (.A1(net6258),
    .A2(_11119_),
    .B1(_11121_),
    .B2(net3173),
    .X(_11123_));
 sky130_fd_sc_hd__a211oi_1 _19287_ (.A1(net3197),
    .A2(net2526),
    .B1(_11123_),
    .C1(net3176),
    .Y(_11124_));
 sky130_fd_sc_hd__nand2_1 _19288_ (.A(net3909),
    .B(net3209),
    .Y(_11125_));
 sky130_fd_sc_hd__a221o_1 _19289_ (.A1(net6313),
    .A2(net3898),
    .B1(_11125_),
    .B2(net6261),
    .C1(net6293),
    .X(_11126_));
 sky130_fd_sc_hd__clkbuf_1 _19290_ (.A(net3205),
    .X(_11127_));
 sky130_fd_sc_hd__o211ai_1 _19291_ (.A1(net2515),
    .A2(net3213),
    .B1(_10941_),
    .C1(net6291),
    .Y(_11128_));
 sky130_fd_sc_hd__a21oi_1 _19292_ (.A1(_11126_),
    .A2(_11128_),
    .B1(net6243),
    .Y(_11129_));
 sky130_fd_sc_hd__o2bb2a_1 _19293_ (.A1_N(net3884),
    .A2_N(net3901),
    .B1(_11124_),
    .B2(_11129_),
    .X(_11130_));
 sky130_fd_sc_hd__or3_1 _19294_ (.A(net3173),
    .B(_10986_),
    .C(_10918_),
    .X(_11131_));
 sky130_fd_sc_hd__clkbuf_1 _19295_ (.A(_10946_),
    .X(_11132_));
 sky130_fd_sc_hd__nand2_1 _19296_ (.A(net6290),
    .B(net6334),
    .Y(_11133_));
 sky130_fd_sc_hd__xnor2_2 _19297_ (.A(net3167),
    .B(_11133_),
    .Y(_11134_));
 sky130_fd_sc_hd__nand2_1 _19298_ (.A(net2512),
    .B(_11134_),
    .Y(_11135_));
 sky130_fd_sc_hd__mux2_1 _19299_ (.A0(net6319),
    .A1(net3191),
    .S(_10986_),
    .X(_11136_));
 sky130_fd_sc_hd__xnor2_1 _19300_ (.A(net6258),
    .B(_10814_),
    .Y(_11137_));
 sky130_fd_sc_hd__mux2_1 _19301_ (.A0(_11136_),
    .A1(_11137_),
    .S(net3887),
    .X(_11138_));
 sky130_fd_sc_hd__mux2_1 _19302_ (.A0(_11134_),
    .A1(_11135_),
    .S(_11138_),
    .X(_11139_));
 sky130_fd_sc_hd__xnor2_2 _19303_ (.A(net6292),
    .B(net6244),
    .Y(_11140_));
 sky130_fd_sc_hd__a21o_1 _19304_ (.A1(net6312),
    .A2(net3888),
    .B1(net6342),
    .X(_11141_));
 sky130_fd_sc_hd__a21bo_1 _19305_ (.A1(net6312),
    .A2(net6352),
    .B1_N(net6338),
    .X(_11142_));
 sky130_fd_sc_hd__o211a_1 _19306_ (.A1(net6312),
    .A2(net6352),
    .B1(_11142_),
    .C1(net6262),
    .X(_11143_));
 sky130_fd_sc_hd__a31o_1 _19307_ (.A1(net3207),
    .A2(_10823_),
    .A3(_11141_),
    .B1(_11143_),
    .X(_11144_));
 sky130_fd_sc_hd__xor2_1 _19308_ (.A(_11140_),
    .B(_11144_),
    .X(_11145_));
 sky130_fd_sc_hd__and3_1 _19309_ (.A(net6224),
    .B(net6290),
    .C(net6334),
    .X(_11146_));
 sky130_fd_sc_hd__nor2_1 _19310_ (.A(net6312),
    .B(net6338),
    .Y(_11147_));
 sky130_fd_sc_hd__a22o_1 _19311_ (.A1(_10985_),
    .A2(_11147_),
    .B1(_10912_),
    .B2(_11051_),
    .X(_11148_));
 sky130_fd_sc_hd__a22o_1 _19312_ (.A1(_11049_),
    .A2(_10838_),
    .B1(_11148_),
    .B2(net6354),
    .X(_11149_));
 sky130_fd_sc_hd__xnor2_2 _19313_ (.A(net3918),
    .B(net2511),
    .Y(_11150_));
 sky130_fd_sc_hd__xnor2_2 _19314_ (.A(_11146_),
    .B(_11150_),
    .Y(_11151_));
 sky130_fd_sc_hd__xor2_1 _19315_ (.A(net2108),
    .B(_11151_),
    .X(_11152_));
 sky130_fd_sc_hd__inv_2 _19316_ (.A(_11152_),
    .Y(_11153_));
 sky130_fd_sc_hd__o22a_1 _19317_ (.A1(net2512),
    .A2(_11134_),
    .B1(_11139_),
    .B2(_11153_),
    .X(_11154_));
 sky130_fd_sc_hd__nor2_1 _19318_ (.A(_11130_),
    .B(_11154_),
    .Y(_11155_));
 sky130_fd_sc_hd__xor2_2 _19319_ (.A(net6186),
    .B(_10930_),
    .X(_11156_));
 sky130_fd_sc_hd__xor2_2 _19320_ (.A(net2523),
    .B(_11054_),
    .X(_11157_));
 sky130_fd_sc_hd__a221o_1 _19321_ (.A1(net6312),
    .A2(net3203),
    .B1(_10823_),
    .B2(_11140_),
    .C1(_11147_),
    .X(_11158_));
 sky130_fd_sc_hd__xnor2_2 _19322_ (.A(net3888),
    .B(net2510),
    .Y(_11159_));
 sky130_fd_sc_hd__xnor2_2 _19323_ (.A(net2107),
    .B(_11159_),
    .Y(_11160_));
 sky130_fd_sc_hd__mux2_1 _19324_ (.A0(_10837_),
    .A1(net3203),
    .S(_11140_),
    .X(_11161_));
 sky130_fd_sc_hd__nand2_1 _19325_ (.A(net6263),
    .B(_11161_),
    .Y(_11162_));
 sky130_fd_sc_hd__mux2_1 _19326_ (.A0(_10821_),
    .A1(net3210),
    .S(_11140_),
    .X(_11163_));
 sky130_fd_sc_hd__nand2_1 _19327_ (.A(net6199),
    .B(net6276),
    .Y(_11164_));
 sky130_fd_sc_hd__o21a_1 _19328_ (.A1(net6263),
    .A2(_11163_),
    .B1(net3871),
    .X(_11165_));
 sky130_fd_sc_hd__mux2_1 _19329_ (.A0(_11162_),
    .A1(_11165_),
    .S(net6315),
    .X(_11166_));
 sky130_fd_sc_hd__o21a_1 _19330_ (.A1(_11156_),
    .A2(_11160_),
    .B1(_11166_),
    .X(_11167_));
 sky130_fd_sc_hd__a21o_1 _19331_ (.A1(_11156_),
    .A2(_11160_),
    .B1(_11167_),
    .X(_11168_));
 sky130_fd_sc_hd__nor2_1 _19332_ (.A(net6352),
    .B(net2525),
    .Y(_11169_));
 sky130_fd_sc_hd__and2_1 _19333_ (.A(net6352),
    .B(net2525),
    .X(_11170_));
 sky130_fd_sc_hd__or2_1 _19334_ (.A(net6262),
    .B(net6229),
    .X(_11171_));
 sky130_fd_sc_hd__mux4_1 _19335_ (.A0(_11169_),
    .A1(_10901_),
    .A2(_11170_),
    .A3(_10900_),
    .S0(_11171_),
    .S1(_11158_),
    .X(_11172_));
 sky130_fd_sc_hd__a31o_1 _19336_ (.A1(net6259),
    .A2(net6230),
    .A3(_11159_),
    .B1(net1752),
    .X(_11173_));
 sky130_fd_sc_hd__o211ai_1 _19337_ (.A1(net3204),
    .A2(_10989_),
    .B1(_11133_),
    .C1(net3167),
    .Y(_11174_));
 sky130_fd_sc_hd__a21boi_1 _19338_ (.A1(net6287),
    .A2(net6334),
    .B1_N(net6270),
    .Y(_11175_));
 sky130_fd_sc_hd__o31a_1 _19339_ (.A1(net3883),
    .A2(_10989_),
    .A3(_11175_),
    .B1(net6320),
    .X(_11176_));
 sky130_fd_sc_hd__nand2_1 _19340_ (.A(net6227),
    .B(net6289),
    .Y(_11177_));
 sky130_fd_sc_hd__a21oi_1 _19341_ (.A1(_10812_),
    .A2(_11177_),
    .B1(_11120_),
    .Y(_11178_));
 sky130_fd_sc_hd__and4b_1 _19342_ (.A_N(net6335),
    .B(_11076_),
    .C(_10812_),
    .D(_11177_),
    .X(_11179_));
 sky130_fd_sc_hd__a211o_1 _19343_ (.A1(_11174_),
    .A2(_11176_),
    .B1(_11178_),
    .C1(_11179_),
    .X(_11180_));
 sky130_fd_sc_hd__a21o_1 _19344_ (.A1(net6179),
    .A2(net6289),
    .B1(net3890),
    .X(_11181_));
 sky130_fd_sc_hd__xnor2_1 _19345_ (.A(_10803_),
    .B(_11181_),
    .Y(_11182_));
 sky130_fd_sc_hd__xnor2_1 _19346_ (.A(_11180_),
    .B(_11182_),
    .Y(_11183_));
 sky130_fd_sc_hd__xnor2_2 _19347_ (.A(net1421),
    .B(_11183_),
    .Y(_11184_));
 sky130_fd_sc_hd__xnor2_1 _19348_ (.A(_11168_),
    .B(_11184_),
    .Y(_11185_));
 sky130_fd_sc_hd__nor2_1 _19349_ (.A(net2108),
    .B(_11151_),
    .Y(_11186_));
 sky130_fd_sc_hd__inv_2 _19350_ (.A(_11138_),
    .Y(_11187_));
 sky130_fd_sc_hd__o21ai_1 _19351_ (.A1(_11187_),
    .A2(_11134_),
    .B1(net2512),
    .Y(_11188_));
 sky130_fd_sc_hd__a21o_1 _19352_ (.A1(net6295),
    .A2(_11147_),
    .B1(_10991_),
    .X(_11189_));
 sky130_fd_sc_hd__or2b_1 _19353_ (.A(net6288),
    .B_N(net6203),
    .X(_11190_));
 sky130_fd_sc_hd__or2b_1 _19354_ (.A(net6202),
    .B_N(net6288),
    .X(_11191_));
 sky130_fd_sc_hd__o22a_1 _19355_ (.A1(_11120_),
    .A2(_11190_),
    .B1(_11191_),
    .B2(net3213),
    .X(_11192_));
 sky130_fd_sc_hd__nor2_1 _19356_ (.A(net3204),
    .B(_11192_),
    .Y(_11193_));
 sky130_fd_sc_hd__a31o_1 _19357_ (.A1(net6202),
    .A2(net2515),
    .A3(net2508),
    .B1(_11193_),
    .X(_11194_));
 sky130_fd_sc_hd__a22o_1 _19358_ (.A1(_11146_),
    .A2(_11150_),
    .B1(_11194_),
    .B2(net6362),
    .X(_11195_));
 sky130_fd_sc_hd__a21oi_1 _19359_ (.A1(_11152_),
    .A2(_11188_),
    .B1(_11195_),
    .Y(_11196_));
 sky130_fd_sc_hd__xor2_1 _19360_ (.A(_11156_),
    .B(_11160_),
    .X(_11197_));
 sky130_fd_sc_hd__xnor2_1 _19361_ (.A(_11166_),
    .B(_11197_),
    .Y(_11198_));
 sky130_fd_sc_hd__and3_1 _19362_ (.A(_11195_),
    .B(_11152_),
    .C(_11188_),
    .X(_11199_));
 sky130_fd_sc_hd__or4_1 _19363_ (.A(_11186_),
    .B(_11196_),
    .C(_11198_),
    .D(_11199_),
    .X(_11200_));
 sky130_fd_sc_hd__xor2_1 _19364_ (.A(_11186_),
    .B(_11198_),
    .X(_11201_));
 sky130_fd_sc_hd__mux2_1 _19365_ (.A0(_11196_),
    .A1(_11199_),
    .S(_11185_),
    .X(_11202_));
 sky130_fd_sc_hd__a2bb2o_1 _19366_ (.A1_N(_11185_),
    .A2_N(_11200_),
    .B1(_11201_),
    .B2(_11202_),
    .X(_11203_));
 sky130_fd_sc_hd__xor2_1 _19367_ (.A(net1753),
    .B(_11089_),
    .X(_11204_));
 sky130_fd_sc_hd__xnor2_1 _19368_ (.A(net1193),
    .B(_11204_),
    .Y(_11205_));
 sky130_fd_sc_hd__and3_1 _19369_ (.A(net6176),
    .B(net6308),
    .C(net6257),
    .X(_11206_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _19370_ (.A(_11206_),
    .X(_11207_));
 sky130_fd_sc_hd__nand2_1 _19371_ (.A(net6152),
    .B(_11207_),
    .Y(_11208_));
 sky130_fd_sc_hd__nor2_1 _19372_ (.A(net6152),
    .B(_11207_),
    .Y(_11209_));
 sky130_fd_sc_hd__nand2_1 _19373_ (.A(net3166),
    .B(net2523),
    .Y(_11210_));
 sky130_fd_sc_hd__nor2_1 _19374_ (.A(_11046_),
    .B(_11207_),
    .Y(_11211_));
 sky130_fd_sc_hd__or2_1 _19375_ (.A(net3166),
    .B(net2523),
    .X(_11212_));
 sky130_fd_sc_hd__o22a_1 _19376_ (.A1(_11209_),
    .A2(_11210_),
    .B1(_11211_),
    .B2(_11212_),
    .X(_11213_));
 sky130_fd_sc_hd__or3b_1 _19377_ (.A(net3166),
    .B(net6152),
    .C_N(_11207_),
    .X(_11214_));
 sky130_fd_sc_hd__o211a_1 _19378_ (.A1(net2509),
    .A2(_11213_),
    .B1(_11214_),
    .C1(net6276),
    .X(_11215_));
 sky130_fd_sc_hd__nand2_1 _19379_ (.A(_11210_),
    .B(_11212_),
    .Y(_11216_));
 sky130_fd_sc_hd__o311a_1 _19380_ (.A1(net2509),
    .A2(_11209_),
    .A3(_11216_),
    .B1(_11208_),
    .C1(net2518),
    .X(_11217_));
 sky130_fd_sc_hd__o22a_1 _19381_ (.A1(net6218),
    .A2(_11208_),
    .B1(_11215_),
    .B2(_11217_),
    .X(_11218_));
 sky130_fd_sc_hd__xnor2_1 _19382_ (.A(net6152),
    .B(_11047_),
    .Y(_11219_));
 sky130_fd_sc_hd__xnor2_1 _19383_ (.A(_11207_),
    .B(_11219_),
    .Y(_11220_));
 sky130_fd_sc_hd__nor2_1 _19384_ (.A(net2509),
    .B(_11157_),
    .Y(_11221_));
 sky130_fd_sc_hd__or2_1 _19385_ (.A(_11220_),
    .B(_11221_),
    .X(_11222_));
 sky130_fd_sc_hd__nand2_1 _19386_ (.A(net2509),
    .B(_11157_),
    .Y(_11223_));
 sky130_fd_sc_hd__o211ai_1 _19387_ (.A1(net6358),
    .A2(_11221_),
    .B1(_11223_),
    .C1(_11220_),
    .Y(_11224_));
 sky130_fd_sc_hd__xnor2_1 _19388_ (.A(_11025_),
    .B(_11180_),
    .Y(_11225_));
 sky130_fd_sc_hd__nor2_1 _19389_ (.A(net6358),
    .B(_11225_),
    .Y(_11226_));
 sky130_fd_sc_hd__a21o_1 _19390_ (.A1(net2509),
    .A2(_11157_),
    .B1(_11220_),
    .X(_11227_));
 sky130_fd_sc_hd__and3_1 _19391_ (.A(net6358),
    .B(_11225_),
    .C(_11227_),
    .X(_11228_));
 sky130_fd_sc_hd__a211o_1 _19392_ (.A1(_11222_),
    .A2(_11224_),
    .B1(_11226_),
    .C1(_11228_),
    .X(_11229_));
 sky130_fd_sc_hd__xor2_1 _19393_ (.A(net1192),
    .B(_11229_),
    .X(_11230_));
 sky130_fd_sc_hd__xnor2_1 _19394_ (.A(net1061),
    .B(_11230_),
    .Y(_11231_));
 sky130_fd_sc_hd__nor2_1 _19395_ (.A(_11168_),
    .B(_11184_),
    .Y(_11232_));
 sky130_fd_sc_hd__xor2_1 _19396_ (.A(_11231_),
    .B(_11232_),
    .X(_11233_));
 sky130_fd_sc_hd__or2_1 _19397_ (.A(net2108),
    .B(_11151_),
    .X(_11234_));
 sky130_fd_sc_hd__o2bb2a_1 _19398_ (.A1_N(_11234_),
    .A2_N(_11196_),
    .B1(_11198_),
    .B2(_11199_),
    .X(_11235_));
 sky130_fd_sc_hd__nand2_1 _19399_ (.A(_11168_),
    .B(_11184_),
    .Y(_11236_));
 sky130_fd_sc_hd__o211a_1 _19400_ (.A1(_11235_),
    .A2(_11232_),
    .B1(_11236_),
    .C1(_11231_),
    .X(_11237_));
 sky130_fd_sc_hd__a31o_1 _19401_ (.A1(_11155_),
    .A2(_11203_),
    .A3(_11233_),
    .B1(_11237_),
    .X(_11238_));
 sky130_fd_sc_hd__a21o_1 _19402_ (.A1(net1192),
    .A2(_11229_),
    .B1(net1061),
    .X(_11239_));
 sky130_fd_sc_hd__o21ai_1 _19403_ (.A1(net1192),
    .A2(_11229_),
    .B1(_11239_),
    .Y(_11240_));
 sky130_fd_sc_hd__and2b_1 _19404_ (.A_N(_11070_),
    .B(_11093_),
    .X(_11241_));
 sky130_fd_sc_hd__xnor2_1 _19405_ (.A(_11092_),
    .B(_11241_),
    .Y(_11242_));
 sky130_fd_sc_hd__o21ai_1 _19406_ (.A1(net812),
    .A2(net869),
    .B1(_11242_),
    .Y(_11243_));
 sky130_fd_sc_hd__inv_2 _19407_ (.A(_11107_),
    .Y(_11244_));
 sky130_fd_sc_hd__or2_1 _19408_ (.A(_11094_),
    .B(_11045_),
    .X(_11245_));
 sky130_fd_sc_hd__nand2_1 _19409_ (.A(_11094_),
    .B(_11045_),
    .Y(_11246_));
 sky130_fd_sc_hd__mux2_1 _19410_ (.A0(_11245_),
    .A1(_11246_),
    .S(_11096_),
    .X(_11247_));
 sky130_fd_sc_hd__or2_1 _19411_ (.A(_11099_),
    .B(_11102_),
    .X(_11248_));
 sky130_fd_sc_hd__mux2_1 _19412_ (.A0(_11248_),
    .A1(_11107_),
    .S(_11096_),
    .X(_11249_));
 sky130_fd_sc_hd__nand2_1 _19413_ (.A(_11245_),
    .B(_11246_),
    .Y(_11250_));
 sky130_fd_sc_hd__o32a_1 _19414_ (.A1(_11103_),
    .A2(_11244_),
    .A3(_11247_),
    .B1(_11249_),
    .B2(_11250_),
    .X(_11251_));
 sky130_fd_sc_hd__or3b_1 _19415_ (.A(_11243_),
    .B(_11251_),
    .C_N(net763),
    .X(_11252_));
 sky130_fd_sc_hd__o21a_1 _19416_ (.A1(_11009_),
    .A2(_10994_),
    .B1(net1426),
    .X(_11253_));
 sky130_fd_sc_hd__a21o_1 _19417_ (.A1(_11009_),
    .A2(_10994_),
    .B1(_11253_),
    .X(_11254_));
 sky130_fd_sc_hd__nand2_1 _19418_ (.A(net6265),
    .B(net3886),
    .Y(_11255_));
 sky130_fd_sc_hd__xnor2_1 _19419_ (.A(net6317),
    .B(_10797_),
    .Y(_11256_));
 sky130_fd_sc_hd__nor2_1 _19420_ (.A(net6265),
    .B(net3886),
    .Y(_11257_));
 sky130_fd_sc_hd__a21o_1 _19421_ (.A1(_11255_),
    .A2(_11256_),
    .B1(_11257_),
    .X(_11258_));
 sky130_fd_sc_hd__nor2_1 _19422_ (.A(net6355),
    .B(_10916_),
    .Y(_11259_));
 sky130_fd_sc_hd__mux2_1 _19423_ (.A0(_11257_),
    .A1(_11259_),
    .S(_10797_),
    .X(_11260_));
 sky130_fd_sc_hd__a21o_1 _19424_ (.A1(net6299),
    .A2(_11258_),
    .B1(_11260_),
    .X(_11261_));
 sky130_fd_sc_hd__and2b_1 _19425_ (.A_N(net6333),
    .B(net6241),
    .X(_11262_));
 sky130_fd_sc_hd__and2b_1 _19426_ (.A_N(net6241),
    .B(net6346),
    .X(_11263_));
 sky130_fd_sc_hd__nor2_2 _19427_ (.A(_11262_),
    .B(_11263_),
    .Y(_11264_));
 sky130_fd_sc_hd__xnor2_4 _19428_ (.A(_10851_),
    .B(_11264_),
    .Y(_11265_));
 sky130_fd_sc_hd__inv_2 _19429_ (.A(_11265_),
    .Y(_11266_));
 sky130_fd_sc_hd__xor2_2 _19430_ (.A(net6070),
    .B(net6105),
    .X(_11267_));
 sky130_fd_sc_hd__or2b_1 _19431_ (.A(net6154),
    .B_N(net6140),
    .X(_11268_));
 sky130_fd_sc_hd__xnor2_1 _19432_ (.A(_11035_),
    .B(_11268_),
    .Y(_11269_));
 sky130_fd_sc_hd__xor2_1 _19433_ (.A(_11267_),
    .B(_11269_),
    .X(_11270_));
 sky130_fd_sc_hd__inv_2 _19434_ (.A(net6148),
    .Y(_11271_));
 sky130_fd_sc_hd__or2_1 _19435_ (.A(net6145),
    .B(net6163),
    .X(_11272_));
 sky130_fd_sc_hd__o21a_1 _19436_ (.A1(net3870),
    .A2(_10971_),
    .B1(_11272_),
    .X(_11273_));
 sky130_fd_sc_hd__nand2_1 _19437_ (.A(net6147),
    .B(net6155),
    .Y(_11274_));
 sky130_fd_sc_hd__a21o_1 _19438_ (.A1(_10971_),
    .A2(_11274_),
    .B1(net6183),
    .X(_11275_));
 sky130_fd_sc_hd__a21o_1 _19439_ (.A1(net3893),
    .A2(_10983_),
    .B1(_10854_),
    .X(_11276_));
 sky130_fd_sc_hd__o21a_1 _19440_ (.A1(_10983_),
    .A2(_10796_),
    .B1(net6209),
    .X(_11277_));
 sky130_fd_sc_hd__a211o_1 _19441_ (.A1(net3161),
    .A2(_11275_),
    .B1(_11276_),
    .C1(_11277_),
    .X(_11278_));
 sky130_fd_sc_hd__o211ai_2 _19442_ (.A1(_11276_),
    .A2(_11277_),
    .B1(net3161),
    .C1(_11275_),
    .Y(_11279_));
 sky130_fd_sc_hd__and3_1 _19443_ (.A(net2507),
    .B(_11278_),
    .C(_11279_),
    .X(_11280_));
 sky130_fd_sc_hd__a21oi_2 _19444_ (.A1(_11278_),
    .A2(_11279_),
    .B1(net2507),
    .Y(_11281_));
 sky130_fd_sc_hd__or3_1 _19445_ (.A(_11266_),
    .B(_11280_),
    .C(_11281_),
    .X(_11282_));
 sky130_fd_sc_hd__o21ai_1 _19446_ (.A1(_11280_),
    .A2(_11281_),
    .B1(_11266_),
    .Y(_11283_));
 sky130_fd_sc_hd__and3_1 _19447_ (.A(_11261_),
    .B(_11282_),
    .C(_11283_),
    .X(_11284_));
 sky130_fd_sc_hd__a21oi_1 _19448_ (.A1(_11282_),
    .A2(_11283_),
    .B1(_11261_),
    .Y(_11285_));
 sky130_fd_sc_hd__or2_1 _19449_ (.A(_11284_),
    .B(_11285_),
    .X(_11286_));
 sky130_fd_sc_hd__a21o_1 _19450_ (.A1(_10982_),
    .A2(net2520),
    .B1(_10988_),
    .X(_11287_));
 sky130_fd_sc_hd__o21a_1 _19451_ (.A1(_10982_),
    .A2(net2520),
    .B1(_11287_),
    .X(_11288_));
 sky130_fd_sc_hd__inv_2 _19452_ (.A(net6025),
    .Y(_11289_));
 sky130_fd_sc_hd__nand2_1 _19453_ (.A(net6119),
    .B(net6086),
    .Y(_11290_));
 sky130_fd_sc_hd__xnor2_1 _19454_ (.A(net3866),
    .B(_11290_),
    .Y(_11291_));
 sky130_fd_sc_hd__nand2_1 _19455_ (.A(net6099),
    .B(net6050),
    .Y(_11292_));
 sky130_fd_sc_hd__nor2_1 _19456_ (.A(net3869),
    .B(_11292_),
    .Y(_11293_));
 sky130_fd_sc_hd__xor2_1 _19457_ (.A(_11291_),
    .B(net3158),
    .X(_11294_));
 sky130_fd_sc_hd__nor2_1 _19458_ (.A(_10974_),
    .B(net2521),
    .Y(_11295_));
 sky130_fd_sc_hd__nand2_1 _19459_ (.A(_10974_),
    .B(net2521),
    .Y(_11296_));
 sky130_fd_sc_hd__o21a_1 _19460_ (.A1(net2522),
    .A2(_11295_),
    .B1(_11296_),
    .X(_11297_));
 sky130_fd_sc_hd__xnor2_1 _19461_ (.A(_11294_),
    .B(_11297_),
    .Y(_11298_));
 sky130_fd_sc_hd__xor2_1 _19462_ (.A(_11288_),
    .B(_11298_),
    .X(_11299_));
 sky130_fd_sc_hd__xnor2_1 _19463_ (.A(_11286_),
    .B(_11299_),
    .Y(_11300_));
 sky130_fd_sc_hd__or2_1 _19464_ (.A(_11254_),
    .B(_11300_),
    .X(_11301_));
 sky130_fd_sc_hd__nand2_1 _19465_ (.A(_11254_),
    .B(_11300_),
    .Y(_11302_));
 sky130_fd_sc_hd__nand2_1 _19466_ (.A(_11301_),
    .B(_11302_),
    .Y(_11303_));
 sky130_fd_sc_hd__a31o_1 _19467_ (.A1(net1064),
    .A2(_11019_),
    .A3(_11020_),
    .B1(_11018_),
    .X(_11304_));
 sky130_fd_sc_hd__a21boi_1 _19468_ (.A1(_11000_),
    .A2(_11006_),
    .B1_N(_11001_),
    .Y(_11305_));
 sky130_fd_sc_hd__or2_1 _19469_ (.A(net960),
    .B(net1420),
    .X(_11306_));
 sky130_fd_sc_hd__nand2_1 _19470_ (.A(net960),
    .B(net1420),
    .Y(_11307_));
 sky130_fd_sc_hd__mux2_1 _19471_ (.A0(net3895),
    .A1(net2514),
    .S(_11265_),
    .X(_11308_));
 sky130_fd_sc_hd__a211o_1 _19472_ (.A1(_11122_),
    .A2(_10984_),
    .B1(_11280_),
    .C1(_11281_),
    .X(_11309_));
 sky130_fd_sc_hd__nor2_1 _19473_ (.A(_11280_),
    .B(_11281_),
    .Y(_11310_));
 sky130_fd_sc_hd__nand2_1 _19474_ (.A(_11266_),
    .B(_11310_),
    .Y(_11311_));
 sky130_fd_sc_hd__a22o_1 _19475_ (.A1(_10984_),
    .A2(_11265_),
    .B1(_11311_),
    .B2(_11122_),
    .X(_11312_));
 sky130_fd_sc_hd__a21oi_1 _19476_ (.A1(net6299),
    .A2(_11265_),
    .B1(_10984_),
    .Y(_11313_));
 sky130_fd_sc_hd__mux2_1 _19477_ (.A0(_10985_),
    .A1(net3895),
    .S(_11265_),
    .X(_11314_));
 sky130_fd_sc_hd__a2bb2o_1 _19478_ (.A1_N(_11310_),
    .A2_N(_11313_),
    .B1(_11314_),
    .B2(net6359),
    .X(_11315_));
 sky130_fd_sc_hd__a221o_1 _19479_ (.A1(_11308_),
    .A2(_11309_),
    .B1(_11312_),
    .B2(_10986_),
    .C1(_11315_),
    .X(_11316_));
 sky130_fd_sc_hd__a211o_1 _19480_ (.A1(_10851_),
    .A2(_11264_),
    .B1(net3196),
    .C1(_11122_),
    .X(_11317_));
 sky130_fd_sc_hd__o21a_1 _19481_ (.A1(_10851_),
    .A2(_11264_),
    .B1(_11317_),
    .X(_11318_));
 sky130_fd_sc_hd__or3b_1 _19482_ (.A(net6297),
    .B(net6359),
    .C_N(_10851_),
    .X(_11319_));
 sky130_fd_sc_hd__mux2_1 _19483_ (.A0(net3196),
    .A1(_11264_),
    .S(_10851_),
    .X(_11320_));
 sky130_fd_sc_hd__o2111a_1 _19484_ (.A1(net6359),
    .A2(_11264_),
    .B1(_11319_),
    .C1(_11320_),
    .D1(net6267),
    .X(_11321_));
 sky130_fd_sc_hd__o21ba_1 _19485_ (.A1(net6267),
    .A2(_11318_),
    .B1_N(_11321_),
    .X(_11322_));
 sky130_fd_sc_hd__mux2_1 _19486_ (.A0(_11262_),
    .A1(_11263_),
    .S(net6272),
    .X(_11323_));
 sky130_fd_sc_hd__nand2_1 _19487_ (.A(_11076_),
    .B(_11075_),
    .Y(_11324_));
 sky130_fd_sc_hd__xnor2_1 _19488_ (.A(_11323_),
    .B(_11324_),
    .Y(_11325_));
 sky130_fd_sc_hd__xnor2_1 _19489_ (.A(net3190),
    .B(_11325_),
    .Y(_11326_));
 sky130_fd_sc_hd__inv_2 _19490_ (.A(_11326_),
    .Y(_11327_));
 sky130_fd_sc_hd__xnor2_2 _19491_ (.A(net6085),
    .B(net6048),
    .Y(_11328_));
 sky130_fd_sc_hd__nor2b_2 _19492_ (.A(net6128),
    .B_N(net6116),
    .Y(_11329_));
 sky130_fd_sc_hd__xnor2_1 _19493_ (.A(net6097),
    .B(_11329_),
    .Y(_11330_));
 sky130_fd_sc_hd__xnor2_1 _19494_ (.A(_11328_),
    .B(_11330_),
    .Y(_11331_));
 sky130_fd_sc_hd__inv_2 _19495_ (.A(_11331_),
    .Y(_11332_));
 sky130_fd_sc_hd__nand2_1 _19496_ (.A(net3168),
    .B(net3897),
    .Y(_11333_));
 sky130_fd_sc_hd__o21ai_1 _19497_ (.A1(_10850_),
    .A2(net3897),
    .B1(net6177),
    .Y(_11334_));
 sky130_fd_sc_hd__o211a_1 _19498_ (.A1(net6182),
    .A2(net6205),
    .B1(_11333_),
    .C1(_11334_),
    .X(_11335_));
 sky130_fd_sc_hd__or2_1 _19499_ (.A(net6116),
    .B(net6128),
    .X(_11336_));
 sky130_fd_sc_hd__a21o_1 _19500_ (.A1(_11267_),
    .A2(_11268_),
    .B1(_11035_),
    .X(_11337_));
 sky130_fd_sc_hd__o211a_1 _19501_ (.A1(net6154),
    .A2(_11267_),
    .B1(_11336_),
    .C1(_11337_),
    .X(_11338_));
 sky130_fd_sc_hd__xnor2_1 _19502_ (.A(_11335_),
    .B(_11338_),
    .Y(_11339_));
 sky130_fd_sc_hd__xnor2_1 _19503_ (.A(_11332_),
    .B(_11339_),
    .Y(_11340_));
 sky130_fd_sc_hd__xnor2_1 _19504_ (.A(_11327_),
    .B(net1419),
    .Y(_11341_));
 sky130_fd_sc_hd__xnor2_2 _19505_ (.A(net1751),
    .B(_11341_),
    .Y(_11342_));
 sky130_fd_sc_hd__nor2_1 _19506_ (.A(_11276_),
    .B(_11277_),
    .Y(_11343_));
 sky130_fd_sc_hd__or2b_1 _19507_ (.A(_11343_),
    .B_N(net2507),
    .X(_11344_));
 sky130_fd_sc_hd__and2b_1 _19508_ (.A_N(net2507),
    .B(_11343_),
    .X(_11345_));
 sky130_fd_sc_hd__a31oi_4 _19509_ (.A1(net3161),
    .A2(_11275_),
    .A3(_11344_),
    .B1(_11345_),
    .Y(_11346_));
 sky130_fd_sc_hd__or2_1 _19510_ (.A(net3866),
    .B(_11290_),
    .X(_11347_));
 sky130_fd_sc_hd__nand2_2 _19511_ (.A(net6067),
    .B(net6103),
    .Y(_11348_));
 sky130_fd_sc_hd__xnor2_1 _19512_ (.A(net4045),
    .B(_11348_),
    .Y(_11349_));
 sky130_fd_sc_hd__xnor2_1 _19513_ (.A(_11347_),
    .B(net3155),
    .Y(_11350_));
 sky130_fd_sc_hd__xnor2_1 _19514_ (.A(_11346_),
    .B(_11350_),
    .Y(_11351_));
 sky130_fd_sc_hd__xnor2_1 _19515_ (.A(_11342_),
    .B(_11351_),
    .Y(_11352_));
 sky130_fd_sc_hd__xnor2_2 _19516_ (.A(net1060),
    .B(_11352_),
    .Y(_11353_));
 sky130_fd_sc_hd__o21ai_1 _19517_ (.A1(net2522),
    .A2(_11295_),
    .B1(_11296_),
    .Y(_11354_));
 sky130_fd_sc_hd__or2_1 _19518_ (.A(_11294_),
    .B(_11354_),
    .X(_11355_));
 sky130_fd_sc_hd__nand2_1 _19519_ (.A(_11294_),
    .B(_11354_),
    .Y(_11356_));
 sky130_fd_sc_hd__or3_1 _19520_ (.A(_11284_),
    .B(_11285_),
    .C(_11298_),
    .X(_11357_));
 sky130_fd_sc_hd__a32o_1 _19521_ (.A1(_11286_),
    .A2(_11355_),
    .A3(_11356_),
    .B1(_11357_),
    .B2(_11288_),
    .X(_11358_));
 sky130_fd_sc_hd__inv_2 _19522_ (.A(_11291_),
    .Y(_11359_));
 sky130_fd_sc_hd__a21o_1 _19523_ (.A1(_11359_),
    .A2(net3158),
    .B1(_11297_),
    .X(_11360_));
 sky130_fd_sc_hd__o21ai_2 _19524_ (.A1(_11359_),
    .A2(net3158),
    .B1(_11360_),
    .Y(_11361_));
 sky130_fd_sc_hd__xor2_1 _19525_ (.A(_11358_),
    .B(_11361_),
    .X(_11362_));
 sky130_fd_sc_hd__xnor2_2 _19526_ (.A(_11353_),
    .B(_11362_),
    .Y(_11363_));
 sky130_fd_sc_hd__mux2_1 _19527_ (.A0(_11306_),
    .A1(_11307_),
    .S(_11363_),
    .X(_11364_));
 sky130_fd_sc_hd__nand2_1 _19528_ (.A(_11307_),
    .B(_11306_),
    .Y(_11365_));
 sky130_fd_sc_hd__mux2_1 _19529_ (.A0(_11302_),
    .A1(_11301_),
    .S(_11363_),
    .X(_11366_));
 sky130_fd_sc_hd__o22a_1 _19530_ (.A1(_11303_),
    .A2(_11364_),
    .B1(_11365_),
    .B2(_11366_),
    .X(_11367_));
 sky130_fd_sc_hd__a31o_1 _19531_ (.A1(_11023_),
    .A2(net713),
    .A3(net712),
    .B1(net709),
    .X(_11368_));
 sky130_fd_sc_hd__a21bo_1 _19532_ (.A1(_11300_),
    .A2(_11307_),
    .B1_N(_11306_),
    .X(_11369_));
 sky130_fd_sc_hd__and2_1 _19533_ (.A(_11254_),
    .B(_11369_),
    .X(_11370_));
 sky130_fd_sc_hd__and2b_1 _19534_ (.A_N(_11306_),
    .B(_11300_),
    .X(_11371_));
 sky130_fd_sc_hd__a21o_1 _19535_ (.A1(net1060),
    .A2(_11342_),
    .B1(_11351_),
    .X(_11372_));
 sky130_fd_sc_hd__o21a_1 _19536_ (.A1(net1060),
    .A2(_11342_),
    .B1(_11372_),
    .X(_11373_));
 sky130_fd_sc_hd__o21a_1 _19537_ (.A1(_11346_),
    .A2(net3155),
    .B1(_11347_),
    .X(_11374_));
 sky130_fd_sc_hd__a21oi_2 _19538_ (.A1(_11346_),
    .A2(net3155),
    .B1(_11374_),
    .Y(_11375_));
 sky130_fd_sc_hd__buf_1 _19539_ (.A(_11035_),
    .X(_11376_));
 sky130_fd_sc_hd__nand2_1 _19540_ (.A(net3153),
    .B(net6098),
    .Y(_11377_));
 sky130_fd_sc_hd__xnor2_1 _19541_ (.A(_10790_),
    .B(_11377_),
    .Y(_11378_));
 sky130_fd_sc_hd__xnor2_2 _19542_ (.A(net6073),
    .B(net6029),
    .Y(_11379_));
 sky130_fd_sc_hd__xnor2_2 _19543_ (.A(net2106),
    .B(_11379_),
    .Y(_11380_));
 sky130_fd_sc_hd__a21o_1 _19544_ (.A1(net6116),
    .A2(net6105),
    .B1(_11328_),
    .X(_11381_));
 sky130_fd_sc_hd__buf_1 _19545_ (.A(net3870),
    .X(_11382_));
 sky130_fd_sc_hd__nor2_1 _19546_ (.A(net6116),
    .B(net6097),
    .Y(_11383_));
 sky130_fd_sc_hd__a221o_1 _19547_ (.A1(net6105),
    .A2(_11328_),
    .B1(_11381_),
    .B2(net3151),
    .C1(_11383_),
    .X(_11384_));
 sky130_fd_sc_hd__or2b_1 _19548_ (.A(_10944_),
    .B_N(_10975_),
    .X(_11385_));
 sky130_fd_sc_hd__a221o_1 _19549_ (.A1(net6158),
    .A2(_10944_),
    .B1(_11385_),
    .B2(net3915),
    .C1(_10977_),
    .X(_11386_));
 sky130_fd_sc_hd__nand2_1 _19550_ (.A(_11384_),
    .B(_11386_),
    .Y(_11387_));
 sky130_fd_sc_hd__or2_1 _19551_ (.A(_11384_),
    .B(_11386_),
    .X(_11388_));
 sky130_fd_sc_hd__nand2_1 _19552_ (.A(_11387_),
    .B(_11388_),
    .Y(_11389_));
 sky130_fd_sc_hd__xnor2_1 _19553_ (.A(_11380_),
    .B(_11389_),
    .Y(_11390_));
 sky130_fd_sc_hd__nor2_1 _19554_ (.A(net6252),
    .B(net3190),
    .Y(_11391_));
 sky130_fd_sc_hd__mux2_1 _19555_ (.A0(net3177),
    .A1(_10938_),
    .S(_11324_),
    .X(_11392_));
 sky130_fd_sc_hd__and2_1 _19556_ (.A(_11076_),
    .B(_11075_),
    .X(_11393_));
 sky130_fd_sc_hd__a211o_1 _19557_ (.A1(_10938_),
    .A2(_11393_),
    .B1(net2513),
    .C1(net6252),
    .X(_11394_));
 sky130_fd_sc_hd__o21ai_1 _19558_ (.A1(net6274),
    .A2(_11392_),
    .B1(_11394_),
    .Y(_11395_));
 sky130_fd_sc_hd__or2_1 _19559_ (.A(net2513),
    .B(_10938_),
    .X(_11396_));
 sky130_fd_sc_hd__nand2_1 _19560_ (.A(net2513),
    .B(_10938_),
    .Y(_11397_));
 sky130_fd_sc_hd__and4_1 _19561_ (.A(net6252),
    .B(_11393_),
    .C(_11396_),
    .D(_11397_),
    .X(_11398_));
 sky130_fd_sc_hd__a221o_1 _19562_ (.A1(_11324_),
    .A2(_11391_),
    .B1(_11395_),
    .B2(net6346),
    .C1(_11398_),
    .X(_11399_));
 sky130_fd_sc_hd__mux2_1 _19563_ (.A0(_11076_),
    .A1(_11075_),
    .S(net3177),
    .X(_11400_));
 sky130_fd_sc_hd__and2_1 _19564_ (.A(_11190_),
    .B(_11191_),
    .X(_11401_));
 sky130_fd_sc_hd__xnor2_1 _19565_ (.A(_11400_),
    .B(_11401_),
    .Y(_11402_));
 sky130_fd_sc_hd__xnor2_2 _19566_ (.A(net3185),
    .B(net2103),
    .Y(_11403_));
 sky130_fd_sc_hd__xnor2_1 _19567_ (.A(net1417),
    .B(_11403_),
    .Y(_11404_));
 sky130_fd_sc_hd__xnor2_2 _19568_ (.A(net1418),
    .B(_11404_),
    .Y(_11405_));
 sky130_fd_sc_hd__a21o_1 _19569_ (.A1(_11332_),
    .A2(_11338_),
    .B1(_11335_),
    .X(_11406_));
 sky130_fd_sc_hd__o21ai_1 _19570_ (.A1(_11332_),
    .A2(_11338_),
    .B1(_11406_),
    .Y(_11407_));
 sky130_fd_sc_hd__nand2_1 _19571_ (.A(net6012),
    .B(_11348_),
    .Y(_11408_));
 sky130_fd_sc_hd__buf_1 _19572_ (.A(_10790_),
    .X(_11409_));
 sky130_fd_sc_hd__buf_1 _19573_ (.A(_10996_),
    .X(_11410_));
 sky130_fd_sc_hd__nor2_1 _19574_ (.A(net3146),
    .B(net3142),
    .Y(_11411_));
 sky130_fd_sc_hd__xnor2_1 _19575_ (.A(_11408_),
    .B(_11411_),
    .Y(_11412_));
 sky130_fd_sc_hd__xnor2_2 _19576_ (.A(net1416),
    .B(_11412_),
    .Y(_11413_));
 sky130_fd_sc_hd__a21bo_1 _19577_ (.A1(_11327_),
    .A2(net1419),
    .B1_N(net1751),
    .X(_11414_));
 sky130_fd_sc_hd__o21a_1 _19578_ (.A1(_11327_),
    .A2(net1419),
    .B1(_11414_),
    .X(_11415_));
 sky130_fd_sc_hd__xnor2_1 _19579_ (.A(_11413_),
    .B(_11415_),
    .Y(_11416_));
 sky130_fd_sc_hd__xnor2_2 _19580_ (.A(_11405_),
    .B(_11416_),
    .Y(_11417_));
 sky130_fd_sc_hd__xor2_1 _19581_ (.A(_11375_),
    .B(_11417_),
    .X(_11418_));
 sky130_fd_sc_hd__xnor2_1 _19582_ (.A(_11373_),
    .B(_11418_),
    .Y(_11419_));
 sky130_fd_sc_hd__nand2_1 _19583_ (.A(_11353_),
    .B(_11361_),
    .Y(_11420_));
 sky130_fd_sc_hd__nor2_1 _19584_ (.A(_11353_),
    .B(_11361_),
    .Y(_11421_));
 sky130_fd_sc_hd__a21o_1 _19585_ (.A1(_11358_),
    .A2(_11420_),
    .B1(_11421_),
    .X(_11422_));
 sky130_fd_sc_hd__nand2_1 _19586_ (.A(_11419_),
    .B(_11422_),
    .Y(_11423_));
 sky130_fd_sc_hd__o31a_1 _19587_ (.A1(_11363_),
    .A2(_11370_),
    .A3(_11371_),
    .B1(_11423_),
    .X(_11424_));
 sky130_fd_sc_hd__nor2_1 _19588_ (.A(_11419_),
    .B(_11422_),
    .Y(_11425_));
 sky130_fd_sc_hd__a21o_1 _19589_ (.A1(net653),
    .A2(_11424_),
    .B1(_11425_),
    .X(_11426_));
 sky130_fd_sc_hd__nor2_1 _19590_ (.A(_11375_),
    .B(_11417_),
    .Y(_11427_));
 sky130_fd_sc_hd__nand2_1 _19591_ (.A(_11375_),
    .B(_11417_),
    .Y(_11428_));
 sky130_fd_sc_hd__o21ai_1 _19592_ (.A1(_11373_),
    .A2(_11427_),
    .B1(_11428_),
    .Y(_11429_));
 sky130_fd_sc_hd__or2_1 _19593_ (.A(_11289_),
    .B(net2106),
    .X(_11430_));
 sky130_fd_sc_hd__buf_1 _19594_ (.A(_11289_),
    .X(_11431_));
 sky130_fd_sc_hd__nand2_1 _19595_ (.A(_11431_),
    .B(net2106),
    .Y(_11432_));
 sky130_fd_sc_hd__inv_2 _19596_ (.A(_11388_),
    .Y(_11433_));
 sky130_fd_sc_hd__a311o_1 _19597_ (.A1(_11387_),
    .A2(_11430_),
    .A3(_11432_),
    .B1(_11433_),
    .C1(net6071),
    .X(_11434_));
 sky130_fd_sc_hd__or3_1 _19598_ (.A(_10995_),
    .B(net2106),
    .C(_11389_),
    .X(_11435_));
 sky130_fd_sc_hd__nand2_1 _19599_ (.A(net6063),
    .B(net6027),
    .Y(_11436_));
 sky130_fd_sc_hd__o22a_1 _19600_ (.A1(net6029),
    .A2(_11387_),
    .B1(_11388_),
    .B2(net3864),
    .X(_11437_));
 sky130_fd_sc_hd__and3_1 _19601_ (.A(_11434_),
    .B(_11435_),
    .C(_11437_),
    .X(_11438_));
 sky130_fd_sc_hd__nand2_1 _19602_ (.A(net6087),
    .B(net6045),
    .Y(_11439_));
 sky130_fd_sc_hd__nand2_1 _19603_ (.A(net6012),
    .B(_11439_),
    .Y(_11440_));
 sky130_fd_sc_hd__xor2_2 _19604_ (.A(_11438_),
    .B(_11440_),
    .X(_11441_));
 sky130_fd_sc_hd__a21bo_1 _19605_ (.A1(net1418),
    .A2(_11403_),
    .B1_N(net1417),
    .X(_11442_));
 sky130_fd_sc_hd__o21a_1 _19606_ (.A1(net1418),
    .A2(_11403_),
    .B1(_11442_),
    .X(_11443_));
 sky130_fd_sc_hd__and2b_1 _19607_ (.A_N(net6097),
    .B(net6085),
    .X(_11444_));
 sky130_fd_sc_hd__xnor2_1 _19608_ (.A(net6065),
    .B(_11444_),
    .Y(_11445_));
 sky130_fd_sc_hd__buf_1 _19609_ (.A(_11445_),
    .X(_11446_));
 sky130_fd_sc_hd__nor2_1 _19610_ (.A(net6050),
    .B(net4046),
    .Y(_11447_));
 sky130_fd_sc_hd__nor2_1 _19611_ (.A(_10996_),
    .B(net6013),
    .Y(_11448_));
 sky130_fd_sc_hd__nor2_2 _19612_ (.A(net3136),
    .B(_11448_),
    .Y(_11449_));
 sky130_fd_sc_hd__xnor2_2 _19613_ (.A(net2505),
    .B(_11449_),
    .Y(_11450_));
 sky130_fd_sc_hd__nand2_1 _19614_ (.A(net6088),
    .B(net6103),
    .Y(_11451_));
 sky130_fd_sc_hd__or2b_1 _19615_ (.A(_11379_),
    .B_N(_11451_),
    .X(_11452_));
 sky130_fd_sc_hd__nor2_1 _19616_ (.A(net6087),
    .B(net6102),
    .Y(_11453_));
 sky130_fd_sc_hd__a221o_1 _19617_ (.A1(net6087),
    .A2(_11379_),
    .B1(_11452_),
    .B2(_11376_),
    .C1(_11453_),
    .X(_11454_));
 sky130_fd_sc_hd__a21o_1 _19618_ (.A1(net3907),
    .A2(net3868),
    .B1(net6183),
    .X(_11455_));
 sky130_fd_sc_hd__o211ai_4 _19619_ (.A1(_11382_),
    .A2(net3907),
    .B1(_11272_),
    .C1(_11455_),
    .Y(_11456_));
 sky130_fd_sc_hd__xnor2_1 _19620_ (.A(_11454_),
    .B(_11456_),
    .Y(_11457_));
 sky130_fd_sc_hd__xnor2_2 _19621_ (.A(_11450_),
    .B(_11457_),
    .Y(_11458_));
 sky130_fd_sc_hd__a21o_1 _19622_ (.A1(net3186),
    .A2(_10918_),
    .B1(_11401_),
    .X(_11459_));
 sky130_fd_sc_hd__or2_1 _19623_ (.A(net3186),
    .B(_10918_),
    .X(_11460_));
 sky130_fd_sc_hd__a21o_1 _19624_ (.A1(_11459_),
    .A2(_11460_),
    .B1(net6221),
    .X(_11461_));
 sky130_fd_sc_hd__mux2_1 _19625_ (.A0(net3176),
    .A1(_10917_),
    .S(net3186),
    .X(_11462_));
 sky130_fd_sc_hd__nand3_1 _19626_ (.A(net6225),
    .B(_11401_),
    .C(_11462_),
    .Y(_11463_));
 sky130_fd_sc_hd__o311a_1 _19627_ (.A1(net3186),
    .A2(_10923_),
    .A3(_11401_),
    .B1(_11461_),
    .C1(_11463_),
    .X(_11464_));
 sky130_fd_sc_hd__mux2_1 _19628_ (.A0(_11190_),
    .A1(_11191_),
    .S(net6222),
    .X(_11465_));
 sky130_fd_sc_hd__xnor2_2 _19629_ (.A(net6178),
    .B(net6269),
    .Y(_11466_));
 sky130_fd_sc_hd__xnor2_1 _19630_ (.A(_11465_),
    .B(_11466_),
    .Y(_11467_));
 sky130_fd_sc_hd__xnor2_1 _19631_ (.A(net3162),
    .B(_11467_),
    .Y(_11468_));
 sky130_fd_sc_hd__xnor2_1 _19632_ (.A(net1749),
    .B(net2101),
    .Y(_11469_));
 sky130_fd_sc_hd__xnor2_2 _19633_ (.A(_11458_),
    .B(_11469_),
    .Y(_11470_));
 sky130_fd_sc_hd__xor2_1 _19634_ (.A(_11443_),
    .B(_11470_),
    .X(_11471_));
 sky130_fd_sc_hd__xnor2_2 _19635_ (.A(_11441_),
    .B(_11471_),
    .Y(_11472_));
 sky130_fd_sc_hd__or2_1 _19636_ (.A(_11348_),
    .B(_11411_),
    .X(_11473_));
 sky130_fd_sc_hd__and3_1 _19637_ (.A(net6012),
    .B(_11348_),
    .C(_11411_),
    .X(_11474_));
 sky130_fd_sc_hd__a221oi_1 _19638_ (.A1(net3291),
    .A2(_11439_),
    .B1(_11473_),
    .B2(net1416),
    .C1(_11474_),
    .Y(_11475_));
 sky130_fd_sc_hd__and2_1 _19639_ (.A(_11413_),
    .B(_11415_),
    .X(_11476_));
 sky130_fd_sc_hd__or2_1 _19640_ (.A(_11413_),
    .B(_11415_),
    .X(_11477_));
 sky130_fd_sc_hd__o21ai_1 _19641_ (.A1(_11405_),
    .A2(_11476_),
    .B1(_11477_),
    .Y(_11478_));
 sky130_fd_sc_hd__xor2_1 _19642_ (.A(net1191),
    .B(_11478_),
    .X(_11479_));
 sky130_fd_sc_hd__xnor2_1 _19643_ (.A(_11472_),
    .B(_11479_),
    .Y(_11480_));
 sky130_fd_sc_hd__nand2_1 _19644_ (.A(_11429_),
    .B(_11480_),
    .Y(_11481_));
 sky130_fd_sc_hd__nor2_1 _19645_ (.A(_11429_),
    .B(_11480_),
    .Y(_11482_));
 sky130_fd_sc_hd__inv_2 _19646_ (.A(_11482_),
    .Y(_11483_));
 sky130_fd_sc_hd__nand2_1 _19647_ (.A(_11481_),
    .B(_11483_),
    .Y(_11484_));
 sky130_fd_sc_hd__xnor2_1 _19648_ (.A(_11426_),
    .B(_11484_),
    .Y(_11485_));
 sky130_fd_sc_hd__nor2_1 _19649_ (.A(_10344_),
    .B(net568),
    .Y(_11486_));
 sky130_fd_sc_hd__a31o_1 _19650_ (.A1(net9049),
    .A2(net2122),
    .A3(net1444),
    .B1(_11486_),
    .X(_00453_));
 sky130_fd_sc_hd__a21bo_1 _19651_ (.A1(net1191),
    .A2(_11472_),
    .B1_N(_11478_),
    .X(_11487_));
 sky130_fd_sc_hd__o21ai_2 _19652_ (.A1(net1191),
    .A2(_11472_),
    .B1(_11487_),
    .Y(_11488_));
 sky130_fd_sc_hd__buf_1 _19653_ (.A(net3880),
    .X(_11489_));
 sky130_fd_sc_hd__nand2_2 _19654_ (.A(net6002),
    .B(net6022),
    .Y(_11490_));
 sky130_fd_sc_hd__nor2_1 _19655_ (.A(net3133),
    .B(net3863),
    .Y(_11491_));
 sky130_fd_sc_hd__nor2_1 _19656_ (.A(_11454_),
    .B(_11456_),
    .Y(_11492_));
 sky130_fd_sc_hd__nand2_1 _19657_ (.A(_11454_),
    .B(_11456_),
    .Y(_11493_));
 sky130_fd_sc_hd__o211a_1 _19658_ (.A1(net2504),
    .A2(_11492_),
    .B1(_11493_),
    .C1(net3135),
    .X(_11494_));
 sky130_fd_sc_hd__xnor2_1 _19659_ (.A(net6012),
    .B(net2504),
    .Y(_11495_));
 sky130_fd_sc_hd__and3_1 _19660_ (.A(net3142),
    .B(net3291),
    .C(net2504),
    .X(_11496_));
 sky130_fd_sc_hd__a21oi_1 _19661_ (.A1(net6045),
    .A2(_11495_),
    .B1(_11496_),
    .Y(_11497_));
 sky130_fd_sc_hd__o22a_1 _19662_ (.A1(_11492_),
    .A2(_11497_),
    .B1(_11493_),
    .B2(net3135),
    .X(_11498_));
 sky130_fd_sc_hd__and2b_1 _19663_ (.A_N(_11494_),
    .B(_11498_),
    .X(_11499_));
 sky130_fd_sc_hd__xnor2_2 _19664_ (.A(net2502),
    .B(_11499_),
    .Y(_11500_));
 sky130_fd_sc_hd__or2_2 _19665_ (.A(net3136),
    .B(_11448_),
    .X(_11501_));
 sky130_fd_sc_hd__a21o_1 _19666_ (.A1(net3201),
    .A2(_11501_),
    .B1(_11409_),
    .X(_11502_));
 sky130_fd_sc_hd__nand2_1 _19667_ (.A(net3881),
    .B(net6102),
    .Y(_11503_));
 sky130_fd_sc_hd__nor3_1 _19668_ (.A(_11409_),
    .B(_11503_),
    .C(_11501_),
    .Y(_11504_));
 sky130_fd_sc_hd__a221o_1 _19669_ (.A1(_11409_),
    .A2(_11501_),
    .B1(_11502_),
    .B2(net6066),
    .C1(_11504_),
    .X(_11505_));
 sky130_fd_sc_hd__nand2_1 _19670_ (.A(net6113),
    .B(net6136),
    .Y(_11506_));
 sky130_fd_sc_hd__a22o_1 _19671_ (.A1(net6198),
    .A2(net6238),
    .B1(net3154),
    .B2(net6156),
    .X(_11507_));
 sky130_fd_sc_hd__o211ai_4 _19672_ (.A1(net6156),
    .A2(_11506_),
    .B1(_11507_),
    .C1(_11336_),
    .Y(_11508_));
 sky130_fd_sc_hd__xnor2_1 _19673_ (.A(net6030),
    .B(_11508_),
    .Y(_11509_));
 sky130_fd_sc_hd__xnor2_1 _19674_ (.A(_11505_),
    .B(_11509_),
    .Y(_11510_));
 sky130_fd_sc_hd__a21o_1 _19675_ (.A1(net3162),
    .A2(_11177_),
    .B1(_11466_),
    .X(_11511_));
 sky130_fd_sc_hd__o21a_1 _19676_ (.A1(net3162),
    .A2(_11177_),
    .B1(_11511_),
    .X(_11512_));
 sky130_fd_sc_hd__nor2_1 _19677_ (.A(net6220),
    .B(net6286),
    .Y(_11513_));
 sky130_fd_sc_hd__mux2_1 _19678_ (.A0(net6220),
    .A1(_11513_),
    .S(net3162),
    .X(_11514_));
 sky130_fd_sc_hd__nand2_1 _19679_ (.A(net6200),
    .B(_11466_),
    .Y(_11515_));
 sky130_fd_sc_hd__or4_1 _19680_ (.A(net6220),
    .B(net3195),
    .C(net3162),
    .D(_11466_),
    .X(_11516_));
 sky130_fd_sc_hd__o221a_1 _19681_ (.A1(net6200),
    .A2(_11512_),
    .B1(_11514_),
    .B2(_11515_),
    .C1(_11516_),
    .X(_11517_));
 sky130_fd_sc_hd__or2_1 _19682_ (.A(net6199),
    .B(net6275),
    .X(_11518_));
 sky130_fd_sc_hd__mux2_1 _19683_ (.A0(_11164_),
    .A1(_11518_),
    .S(net6176),
    .X(_11519_));
 sky130_fd_sc_hd__nor2_1 _19684_ (.A(_11046_),
    .B(net6257),
    .Y(_11520_));
 sky130_fd_sc_hd__nor2_1 _19685_ (.A(net6151),
    .B(net3175),
    .Y(_11521_));
 sky130_fd_sc_hd__nor2_2 _19686_ (.A(_11520_),
    .B(_11521_),
    .Y(_11522_));
 sky130_fd_sc_hd__xnor2_1 _19687_ (.A(_11519_),
    .B(_11522_),
    .Y(_11523_));
 sky130_fd_sc_hd__xnor2_2 _19688_ (.A(net3157),
    .B(_11523_),
    .Y(_11524_));
 sky130_fd_sc_hd__xor2_1 _19689_ (.A(_11517_),
    .B(_11524_),
    .X(_11525_));
 sky130_fd_sc_hd__xnor2_1 _19690_ (.A(net1415),
    .B(_11525_),
    .Y(_11526_));
 sky130_fd_sc_hd__o21a_1 _19691_ (.A1(_11458_),
    .A2(net2101),
    .B1(net1749),
    .X(_11527_));
 sky130_fd_sc_hd__a21oi_1 _19692_ (.A1(_11458_),
    .A2(net2101),
    .B1(_11527_),
    .Y(_11528_));
 sky130_fd_sc_hd__nor2_1 _19693_ (.A(net1058),
    .B(_11528_),
    .Y(_11529_));
 sky130_fd_sc_hd__nand2_1 _19694_ (.A(net1058),
    .B(_11528_),
    .Y(_11530_));
 sky130_fd_sc_hd__and2b_1 _19695_ (.A_N(_11529_),
    .B(_11530_),
    .X(_11531_));
 sky130_fd_sc_hd__xnor2_2 _19696_ (.A(_11500_),
    .B(_11531_),
    .Y(_11532_));
 sky130_fd_sc_hd__a21o_1 _19697_ (.A1(_11443_),
    .A2(_11470_),
    .B1(_11441_),
    .X(_11533_));
 sky130_fd_sc_hd__o21ai_2 _19698_ (.A1(_11443_),
    .A2(_11470_),
    .B1(_11533_),
    .Y(_11534_));
 sky130_fd_sc_hd__nor2_1 _19699_ (.A(net3131),
    .B(net3138),
    .Y(_11535_));
 sky130_fd_sc_hd__nor2_1 _19700_ (.A(_11439_),
    .B(_11535_),
    .Y(_11536_));
 sky130_fd_sc_hd__o21a_1 _19701_ (.A1(_11380_),
    .A2(_11384_),
    .B1(_11386_),
    .X(_11537_));
 sky130_fd_sc_hd__a21oi_1 _19702_ (.A1(_11380_),
    .A2(_11384_),
    .B1(_11537_),
    .Y(_11538_));
 sky130_fd_sc_hd__or3_1 _19703_ (.A(net3291),
    .B(_11411_),
    .C(net3864),
    .X(_11539_));
 sky130_fd_sc_hd__o221a_1 _19704_ (.A1(net6012),
    .A2(_11535_),
    .B1(_11536_),
    .B2(_11538_),
    .C1(_11539_),
    .X(_11540_));
 sky130_fd_sc_hd__xor2_1 _19705_ (.A(_11534_),
    .B(net1057),
    .X(_11541_));
 sky130_fd_sc_hd__xnor2_2 _19706_ (.A(_11532_),
    .B(_11541_),
    .Y(_11542_));
 sky130_fd_sc_hd__nand2_1 _19707_ (.A(_11488_),
    .B(_11542_),
    .Y(_11543_));
 sky130_fd_sc_hd__inv_2 _19708_ (.A(_11543_),
    .Y(_11544_));
 sky130_fd_sc_hd__nor2_1 _19709_ (.A(_11488_),
    .B(_11542_),
    .Y(_11545_));
 sky130_fd_sc_hd__nor2_1 _19710_ (.A(_11544_),
    .B(_11545_),
    .Y(_11546_));
 sky130_fd_sc_hd__a21o_1 _19711_ (.A1(_11425_),
    .A2(_11481_),
    .B1(_11482_),
    .X(_11547_));
 sky130_fd_sc_hd__a31o_1 _19712_ (.A1(net653),
    .A2(_11424_),
    .A3(_11481_),
    .B1(_11547_),
    .X(_11548_));
 sky130_fd_sc_hd__xnor2_1 _19713_ (.A(net6382),
    .B(net6386),
    .Y(_11549_));
 sky130_fd_sc_hd__or2_1 _19714_ (.A(net570),
    .B(net3857),
    .X(_11550_));
 sky130_fd_sc_hd__xnor2_1 _19715_ (.A(_11548_),
    .B(_11550_),
    .Y(_11551_));
 sky130_fd_sc_hd__xnor2_1 _19716_ (.A(_11546_),
    .B(_11551_),
    .Y(_11552_));
 sky130_fd_sc_hd__a22o_1 _19717_ (.A1(net9029),
    .A2(net1199),
    .B1(_11552_),
    .B2(net1767),
    .X(_00454_));
 sky130_fd_sc_hd__or2_1 _19718_ (.A(_11488_),
    .B(_11542_),
    .X(_11553_));
 sky130_fd_sc_hd__a22o_1 _19719_ (.A1(net569),
    .A2(_11544_),
    .B1(_11553_),
    .B2(net3857),
    .X(_11554_));
 sky130_fd_sc_hd__nand2_1 _19720_ (.A(net604),
    .B(_11554_),
    .Y(_11555_));
 sky130_fd_sc_hd__o21a_1 _19721_ (.A1(_11544_),
    .A2(net604),
    .B1(_11553_),
    .X(_11556_));
 sky130_fd_sc_hd__o22a_1 _19722_ (.A1(_11553_),
    .A2(net604),
    .B1(_11556_),
    .B2(net569),
    .X(_11557_));
 sky130_fd_sc_hd__mux2_1 _19723_ (.A0(_11557_),
    .A1(_11543_),
    .S(net3857),
    .X(_11558_));
 sky130_fd_sc_hd__nor2b_1 _19724_ (.A(net6080),
    .B_N(net6062),
    .Y(_11559_));
 sky130_fd_sc_hd__inv_2 _19725_ (.A(net3856),
    .Y(_11560_));
 sky130_fd_sc_hd__mux2_1 _19726_ (.A0(_11449_),
    .A1(_11508_),
    .S(_11431_),
    .X(_11561_));
 sky130_fd_sc_hd__nand2_1 _19727_ (.A(net6030),
    .B(_11449_),
    .Y(_11562_));
 sky130_fd_sc_hd__nand2_1 _19728_ (.A(_11431_),
    .B(_11501_),
    .Y(_11563_));
 sky130_fd_sc_hd__o21a_1 _19729_ (.A1(net6066),
    .A2(_11562_),
    .B1(_11563_),
    .X(_11564_));
 sky130_fd_sc_hd__a21oi_1 _19730_ (.A1(_11508_),
    .A2(_11562_),
    .B1(_11503_),
    .Y(_11565_));
 sky130_fd_sc_hd__nand2_1 _19731_ (.A(net6030),
    .B(_11508_),
    .Y(_11566_));
 sky130_fd_sc_hd__or3_1 _19732_ (.A(net3881),
    .B(net6099),
    .C(_11449_),
    .X(_11567_));
 sky130_fd_sc_hd__o211a_1 _19733_ (.A1(net6030),
    .A2(_11501_),
    .B1(_11566_),
    .C1(_11567_),
    .X(_11568_));
 sky130_fd_sc_hd__o21ai_1 _19734_ (.A1(_11565_),
    .A2(_11568_),
    .B1(net6084),
    .Y(_11569_));
 sky130_fd_sc_hd__o221a_1 _19735_ (.A1(_11560_),
    .A2(_11561_),
    .B1(_11564_),
    .B2(_11508_),
    .C1(_11569_),
    .X(_11570_));
 sky130_fd_sc_hd__nand2_1 _19736_ (.A(net6045),
    .B(net3138),
    .Y(_11571_));
 sky130_fd_sc_hd__nand2_1 _19737_ (.A(net3879),
    .B(net6026),
    .Y(_11572_));
 sky130_fd_sc_hd__and3_1 _19738_ (.A(net6008),
    .B(_11571_),
    .C(net3129),
    .X(_11573_));
 sky130_fd_sc_hd__xor2_2 _19739_ (.A(net1056),
    .B(_11573_),
    .X(_11574_));
 sky130_fd_sc_hd__a21o_1 _19740_ (.A1(net3157),
    .A2(_11522_),
    .B1(_11164_),
    .X(_11575_));
 sky130_fd_sc_hd__o21a_1 _19741_ (.A1(net3157),
    .A2(_11522_),
    .B1(_11575_),
    .X(_11576_));
 sky130_fd_sc_hd__a21bo_1 _19742_ (.A1(_11518_),
    .A2(_11522_),
    .B1_N(net3157),
    .X(_11577_));
 sky130_fd_sc_hd__o22a_1 _19743_ (.A1(net3919),
    .A2(net3157),
    .B1(_11522_),
    .B2(net6275),
    .X(_11578_));
 sky130_fd_sc_hd__nand2_1 _19744_ (.A(_11577_),
    .B(_11578_),
    .Y(_11579_));
 sky130_fd_sc_hd__mux2_1 _19745_ (.A0(_11576_),
    .A1(_11579_),
    .S(net6176),
    .X(_11580_));
 sky130_fd_sc_hd__a22o_1 _19746_ (.A1(net3175),
    .A2(_10972_),
    .B1(_11521_),
    .B2(net6175),
    .X(_11581_));
 sky130_fd_sc_hd__xnor2_2 _19747_ (.A(net6219),
    .B(net6131),
    .Y(_11582_));
 sky130_fd_sc_hd__xor2_1 _19748_ (.A(net2104),
    .B(_11582_),
    .X(_11583_));
 sky130_fd_sc_hd__xnor2_2 _19749_ (.A(_11581_),
    .B(_11583_),
    .Y(_11584_));
 sky130_fd_sc_hd__o2bb2a_1 _19750_ (.A1_N(net6171),
    .A2_N(net6198),
    .B1(net3150),
    .B2(net6097),
    .X(_11585_));
 sky130_fd_sc_hd__a211oi_2 _19751_ (.A1(net6097),
    .A2(_11329_),
    .B1(_11383_),
    .C1(_11585_),
    .Y(_11586_));
 sky130_fd_sc_hd__a211o_1 _19752_ (.A1(net6050),
    .A2(net6030),
    .B1(net3136),
    .C1(net6088),
    .X(_11587_));
 sky130_fd_sc_hd__nand2_2 _19753_ (.A(net6046),
    .B(net4045),
    .Y(_11588_));
 sky130_fd_sc_hd__a21o_1 _19754_ (.A1(_11588_),
    .A2(net3129),
    .B1(net3146),
    .X(_11589_));
 sky130_fd_sc_hd__a21oi_1 _19755_ (.A1(_11588_),
    .A2(net3129),
    .B1(net6067),
    .Y(_11590_));
 sky130_fd_sc_hd__a31o_1 _19756_ (.A1(net6072),
    .A2(_11587_),
    .A3(_11589_),
    .B1(_11590_),
    .X(_11591_));
 sky130_fd_sc_hd__xnor2_2 _19757_ (.A(_11586_),
    .B(net2099),
    .Y(_11592_));
 sky130_fd_sc_hd__xor2_1 _19758_ (.A(_11584_),
    .B(_11592_),
    .X(_11593_));
 sky130_fd_sc_hd__xnor2_1 _19759_ (.A(_11580_),
    .B(_11593_),
    .Y(_11594_));
 sky130_fd_sc_hd__a21o_1 _19760_ (.A1(_11517_),
    .A2(_11524_),
    .B1(net1415),
    .X(_11595_));
 sky130_fd_sc_hd__o21ai_1 _19761_ (.A1(_11517_),
    .A2(_11524_),
    .B1(_11595_),
    .Y(_11596_));
 sky130_fd_sc_hd__nor2_1 _19762_ (.A(_11594_),
    .B(_11596_),
    .Y(_11597_));
 sky130_fd_sc_hd__nand2_1 _19763_ (.A(_11594_),
    .B(_11596_),
    .Y(_11598_));
 sky130_fd_sc_hd__or2b_1 _19764_ (.A(net958),
    .B_N(net956),
    .X(_11599_));
 sky130_fd_sc_hd__xnor2_2 _19765_ (.A(_11574_),
    .B(_11599_),
    .Y(_11600_));
 sky130_fd_sc_hd__a21o_1 _19766_ (.A1(_11500_),
    .A2(_11530_),
    .B1(_11529_),
    .X(_11601_));
 sky130_fd_sc_hd__inv_2 _19767_ (.A(net2504),
    .Y(_11602_));
 sky130_fd_sc_hd__a21o_1 _19768_ (.A1(_11602_),
    .A2(_11493_),
    .B1(net3135),
    .X(_11603_));
 sky130_fd_sc_hd__o21ai_2 _19769_ (.A1(net2502),
    .A2(_11494_),
    .B1(_11603_),
    .Y(_11604_));
 sky130_fd_sc_hd__xnor2_1 _19770_ (.A(_11601_),
    .B(_11604_),
    .Y(_11605_));
 sky130_fd_sc_hd__xnor2_2 _19771_ (.A(_11600_),
    .B(_11605_),
    .Y(_11606_));
 sky130_fd_sc_hd__a21o_1 _19772_ (.A1(_11534_),
    .A2(net1057),
    .B1(_11532_),
    .X(_11607_));
 sky130_fd_sc_hd__o21a_1 _19773_ (.A1(_11534_),
    .A2(net1057),
    .B1(_11607_),
    .X(_11608_));
 sky130_fd_sc_hd__xnor2_2 _19774_ (.A(_11606_),
    .B(_11608_),
    .Y(_11609_));
 sky130_fd_sc_hd__a21o_1 _19775_ (.A1(_11555_),
    .A2(_11558_),
    .B1(_11609_),
    .X(_11610_));
 sky130_fd_sc_hd__nand3_1 _19776_ (.A(_11609_),
    .B(_11555_),
    .C(_11558_),
    .Y(_11611_));
 sky130_fd_sc_hd__and3_1 _19777_ (.A(\cordic0.cos[2] ),
    .B(net2942),
    .C(net1782),
    .X(_11612_));
 sky130_fd_sc_hd__a31o_1 _19778_ (.A1(net1767),
    .A2(_11610_),
    .A3(_11611_),
    .B1(_11612_),
    .X(_00455_));
 sky130_fd_sc_hd__nand2_1 _19779_ (.A(_11542_),
    .B(net604),
    .Y(_11613_));
 sky130_fd_sc_hd__or2_1 _19780_ (.A(_11542_),
    .B(net604),
    .X(_11614_));
 sky130_fd_sc_hd__and2b_1 _19781_ (.A_N(_11488_),
    .B(_11609_),
    .X(_11615_));
 sky130_fd_sc_hd__or3b_1 _19782_ (.A(_11542_),
    .B(net604),
    .C_N(_11609_),
    .X(_11616_));
 sky130_fd_sc_hd__nand3b_1 _19783_ (.A_N(_11609_),
    .B(net604),
    .C(_11542_),
    .Y(_11617_));
 sky130_fd_sc_hd__nand2_1 _19784_ (.A(_11616_),
    .B(_11617_),
    .Y(_11618_));
 sky130_fd_sc_hd__a32o_1 _19785_ (.A1(_11613_),
    .A2(_11614_),
    .A3(_11615_),
    .B1(_11618_),
    .B2(_11488_),
    .X(_11619_));
 sky130_fd_sc_hd__buf_1 _19786_ (.A(net3859),
    .X(_11620_));
 sky130_fd_sc_hd__a21oi_1 _19787_ (.A1(net568),
    .A2(net488),
    .B1(_11620_),
    .Y(_11621_));
 sky130_fd_sc_hd__o21a_1 _19788_ (.A1(_11584_),
    .A2(_11592_),
    .B1(_11580_),
    .X(_11622_));
 sky130_fd_sc_hd__a21oi_1 _19789_ (.A1(_11584_),
    .A2(_11592_),
    .B1(_11622_),
    .Y(_11623_));
 sky130_fd_sc_hd__o211a_1 _19790_ (.A1(net6088),
    .A2(net3136),
    .B1(_11588_),
    .C1(net2100),
    .X(_11624_));
 sky130_fd_sc_hd__a21o_1 _19791_ (.A1(net6088),
    .A2(net3141),
    .B1(net2100),
    .X(_11625_));
 sky130_fd_sc_hd__or2b_1 _19792_ (.A(net3862),
    .B_N(_11625_),
    .X(_11626_));
 sky130_fd_sc_hd__o211a_1 _19793_ (.A1(net6032),
    .A2(_11624_),
    .B1(_11626_),
    .C1(net6067),
    .X(_11627_));
 sky130_fd_sc_hd__a21oi_1 _19794_ (.A1(net6008),
    .A2(net2100),
    .B1(net3138),
    .Y(_11628_));
 sky130_fd_sc_hd__o221a_1 _19795_ (.A1(net6008),
    .A2(net2100),
    .B1(_11628_),
    .B2(net6043),
    .C1(net3130),
    .X(_11629_));
 sky130_fd_sc_hd__or4_1 _19796_ (.A(net6088),
    .B(net3141),
    .C(net6016),
    .D(net2100),
    .X(_11630_));
 sky130_fd_sc_hd__o21ai_4 _19797_ (.A1(_11627_),
    .A2(_11629_),
    .B1(_11630_),
    .Y(_11631_));
 sky130_fd_sc_hd__mux2_1 _19798_ (.A0(net2104),
    .A1(_11046_),
    .S(_11582_),
    .X(_11632_));
 sky130_fd_sc_hd__a21o_1 _19799_ (.A1(net2104),
    .A2(_11582_),
    .B1(net6151),
    .X(_11633_));
 sky130_fd_sc_hd__mux2_1 _19800_ (.A0(_11632_),
    .A1(_11633_),
    .S(net6170),
    .X(_11634_));
 sky130_fd_sc_hd__or3_1 _19801_ (.A(net6151),
    .B(net2104),
    .C(_11582_),
    .X(_11635_));
 sky130_fd_sc_hd__xnor2_1 _19802_ (.A(net6170),
    .B(net2104),
    .Y(_11636_));
 sky130_fd_sc_hd__nand3_1 _19803_ (.A(net6151),
    .B(_11582_),
    .C(_11636_),
    .Y(_11637_));
 sky130_fd_sc_hd__o211a_1 _19804_ (.A1(net3174),
    .A2(_11634_),
    .B1(_11635_),
    .C1(_11637_),
    .X(_11638_));
 sky130_fd_sc_hd__or2_1 _19805_ (.A(net6215),
    .B(net6157),
    .X(_11639_));
 sky130_fd_sc_hd__nand2_1 _19806_ (.A(net6215),
    .B(net6157),
    .Y(_11640_));
 sky130_fd_sc_hd__mux2_1 _19807_ (.A0(_11639_),
    .A1(_11640_),
    .S(net3150),
    .X(_11641_));
 sky130_fd_sc_hd__xnor2_2 _19808_ (.A(net6214),
    .B(net6117),
    .Y(_11642_));
 sky130_fd_sc_hd__xnor2_1 _19809_ (.A(_11641_),
    .B(_11642_),
    .Y(_11643_));
 sky130_fd_sc_hd__xnor2_1 _19810_ (.A(net2506),
    .B(_11643_),
    .Y(_11644_));
 sky130_fd_sc_hd__nand2_1 _19811_ (.A(net6121),
    .B(net3913),
    .Y(_11645_));
 sky130_fd_sc_hd__nor2_1 _19812_ (.A(net6121),
    .B(_11451_),
    .Y(_11646_));
 sky130_fd_sc_hd__a211o_1 _19813_ (.A1(_11645_),
    .A2(_10975_),
    .B1(_11453_),
    .C1(_11646_),
    .X(_11647_));
 sky130_fd_sc_hd__nand2_1 _19814_ (.A(net6068),
    .B(net6041),
    .Y(_11648_));
 sky130_fd_sc_hd__o21a_1 _19815_ (.A1(net6034),
    .A2(_11648_),
    .B1(net3128),
    .X(_11649_));
 sky130_fd_sc_hd__xnor2_1 _19816_ (.A(net6010),
    .B(_11649_),
    .Y(_11650_));
 sky130_fd_sc_hd__xnor2_1 _19817_ (.A(net2500),
    .B(_11650_),
    .Y(_11651_));
 sky130_fd_sc_hd__xor2_1 _19818_ (.A(net1747),
    .B(_11651_),
    .X(_11652_));
 sky130_fd_sc_hd__xnor2_2 _19819_ (.A(net1188),
    .B(_11652_),
    .Y(_11653_));
 sky130_fd_sc_hd__xor2_2 _19820_ (.A(_11631_),
    .B(_11653_),
    .X(_11654_));
 sky130_fd_sc_hd__xnor2_4 _19821_ (.A(net953),
    .B(_11654_),
    .Y(_11655_));
 sky130_fd_sc_hd__o21ai_2 _19822_ (.A1(_11574_),
    .A2(net958),
    .B1(net956),
    .Y(_11656_));
 sky130_fd_sc_hd__a21o_1 _19823_ (.A1(net6037),
    .A2(net1056),
    .B1(net3141),
    .X(_11657_));
 sky130_fd_sc_hd__or2_1 _19824_ (.A(net6032),
    .B(net1056),
    .X(_11658_));
 sky130_fd_sc_hd__a21o_1 _19825_ (.A1(_11657_),
    .A2(_11658_),
    .B1(net3291),
    .X(_11659_));
 sky130_fd_sc_hd__xnor2_2 _19826_ (.A(_11656_),
    .B(_11659_),
    .Y(_11660_));
 sky130_fd_sc_hd__xnor2_4 _19827_ (.A(_11655_),
    .B(_11660_),
    .Y(_11661_));
 sky130_fd_sc_hd__and2b_1 _19828_ (.A_N(_11606_),
    .B(_11608_),
    .X(_11662_));
 sky130_fd_sc_hd__nor2_1 _19829_ (.A(_11545_),
    .B(_11662_),
    .Y(_11663_));
 sky130_fd_sc_hd__or2b_1 _19830_ (.A(_11608_),
    .B_N(_11606_),
    .X(_11664_));
 sky130_fd_sc_hd__o21ai_1 _19831_ (.A1(_11543_),
    .A2(_11662_),
    .B1(_11664_),
    .Y(_11665_));
 sky130_fd_sc_hd__a21oi_1 _19832_ (.A1(net604),
    .A2(_11663_),
    .B1(_11665_),
    .Y(_11666_));
 sky130_fd_sc_hd__buf_2 _19833_ (.A(net567),
    .X(_11667_));
 sky130_fd_sc_hd__o21a_1 _19834_ (.A1(_11601_),
    .A2(_11604_),
    .B1(_11600_),
    .X(_11668_));
 sky130_fd_sc_hd__a21oi_1 _19835_ (.A1(_11601_),
    .A2(_11604_),
    .B1(_11668_),
    .Y(_11669_));
 sky130_fd_sc_hd__xnor2_1 _19836_ (.A(_11667_),
    .B(net708),
    .Y(_11670_));
 sky130_fd_sc_hd__xor2_1 _19837_ (.A(_11661_),
    .B(_11670_),
    .X(_11671_));
 sky130_fd_sc_hd__xnor2_1 _19838_ (.A(_11621_),
    .B(_11671_),
    .Y(_11672_));
 sky130_fd_sc_hd__a22o_1 _19839_ (.A1(net8968),
    .A2(net1200),
    .B1(_11672_),
    .B2(net1768),
    .X(_00456_));
 sky130_fd_sc_hd__o21ba_1 _19840_ (.A1(_11631_),
    .A2(_11653_),
    .B1_N(net953),
    .X(_11673_));
 sky130_fd_sc_hd__a21oi_2 _19841_ (.A1(_11631_),
    .A2(_11653_),
    .B1(_11673_),
    .Y(_11674_));
 sky130_fd_sc_hd__or2b_1 _19842_ (.A(net1747),
    .B_N(_11651_),
    .X(_11675_));
 sky130_fd_sc_hd__and2b_1 _19843_ (.A_N(_11651_),
    .B(net1747),
    .X(_11676_));
 sky130_fd_sc_hd__a21oi_1 _19844_ (.A1(net1188),
    .A2(_11675_),
    .B1(_11676_),
    .Y(_11677_));
 sky130_fd_sc_hd__mux2_1 _19845_ (.A0(net2506),
    .A1(net6130),
    .S(net6157),
    .X(_11678_));
 sky130_fd_sc_hd__or3b_1 _19846_ (.A(net6128),
    .B(_11445_),
    .C_N(net6157),
    .X(_11679_));
 sky130_fd_sc_hd__o21a_1 _19847_ (.A1(_11642_),
    .A2(_11678_),
    .B1(_11679_),
    .X(_11680_));
 sky130_fd_sc_hd__nor2_1 _19848_ (.A(net6157),
    .B(net2506),
    .Y(_11681_));
 sky130_fd_sc_hd__a21oi_1 _19849_ (.A1(net2506),
    .A2(_11639_),
    .B1(_11681_),
    .Y(_11682_));
 sky130_fd_sc_hd__nand2_1 _19850_ (.A(net6127),
    .B(_11642_),
    .Y(_11683_));
 sky130_fd_sc_hd__or3_1 _19851_ (.A(net6127),
    .B(net2506),
    .C(_11642_),
    .X(_11684_));
 sky130_fd_sc_hd__o221a_1 _19852_ (.A1(net3165),
    .A2(_11680_),
    .B1(_11682_),
    .B2(_11683_),
    .C1(_11684_),
    .X(_11685_));
 sky130_fd_sc_hd__xnor2_4 _19853_ (.A(net6049),
    .B(net3856),
    .Y(_11686_));
 sky130_fd_sc_hd__nand3b_1 _19854_ (.A_N(net6110),
    .B(net6127),
    .C(net6212),
    .Y(_11687_));
 sky130_fd_sc_hd__or3b_1 _19855_ (.A(net6212),
    .B(net6135),
    .C_N(net6110),
    .X(_11688_));
 sky130_fd_sc_hd__nand2_1 _19856_ (.A(_11687_),
    .B(_11688_),
    .Y(_11689_));
 sky130_fd_sc_hd__xnor2_2 _19857_ (.A(net6169),
    .B(net6098),
    .Y(_11690_));
 sky130_fd_sc_hd__xor2_1 _19858_ (.A(_11689_),
    .B(_11690_),
    .X(_11691_));
 sky130_fd_sc_hd__xnor2_1 _19859_ (.A(_11686_),
    .B(_11691_),
    .Y(_11692_));
 sky130_fd_sc_hd__a21o_1 _19860_ (.A1(net6066),
    .A2(net3201),
    .B1(_10790_),
    .X(_11693_));
 sky130_fd_sc_hd__a22o_1 _19861_ (.A1(_11503_),
    .A2(net3867),
    .B1(_11560_),
    .B2(_11693_),
    .X(_11694_));
 sky130_fd_sc_hd__o21ai_1 _19862_ (.A1(net6041),
    .A2(net6010),
    .B1(net6031),
    .Y(_11695_));
 sky130_fd_sc_hd__xnor2_1 _19863_ (.A(net2095),
    .B(_11695_),
    .Y(_11696_));
 sky130_fd_sc_hd__xnor2_1 _19864_ (.A(net2097),
    .B(_11696_),
    .Y(_11697_));
 sky130_fd_sc_hd__xnor2_2 _19865_ (.A(net1412),
    .B(_11697_),
    .Y(_11698_));
 sky130_fd_sc_hd__o21ai_1 _19866_ (.A1(net3130),
    .A2(net6033),
    .B1(net2501),
    .Y(_11699_));
 sky130_fd_sc_hd__mux2_1 _19867_ (.A0(net6033),
    .A1(net6009),
    .S(net2501),
    .X(_11700_));
 sky130_fd_sc_hd__inv_2 _19868_ (.A(_11700_),
    .Y(_11701_));
 sky130_fd_sc_hd__or4_1 _19869_ (.A(net6009),
    .B(net6033),
    .C(net2500),
    .D(_11648_),
    .X(_11702_));
 sky130_fd_sc_hd__o221a_1 _19870_ (.A1(net3292),
    .A2(_11699_),
    .B1(_11701_),
    .B2(net6043),
    .C1(_11702_),
    .X(_11703_));
 sky130_fd_sc_hd__xnor2_1 _19871_ (.A(_11698_),
    .B(_11703_),
    .Y(_11704_));
 sky130_fd_sc_hd__xnor2_1 _19872_ (.A(_11677_),
    .B(_11704_),
    .Y(_11705_));
 sky130_fd_sc_hd__a22o_1 _19873_ (.A1(net3141),
    .A2(net2100),
    .B1(_11625_),
    .B2(net6064),
    .X(_11706_));
 sky130_fd_sc_hd__and3_1 _19874_ (.A(net6016),
    .B(net6033),
    .C(_11706_),
    .X(_11707_));
 sky130_fd_sc_hd__nand2_1 _19875_ (.A(_11705_),
    .B(_11707_),
    .Y(_11708_));
 sky130_fd_sc_hd__nor2_1 _19876_ (.A(_11705_),
    .B(_11707_),
    .Y(_11709_));
 sky130_fd_sc_hd__inv_2 _19877_ (.A(_11709_),
    .Y(_11710_));
 sky130_fd_sc_hd__nand2_1 _19878_ (.A(_11708_),
    .B(_11710_),
    .Y(_11711_));
 sky130_fd_sc_hd__xnor2_2 _19879_ (.A(_11674_),
    .B(_11711_),
    .Y(_11712_));
 sky130_fd_sc_hd__a21bo_1 _19880_ (.A1(_11655_),
    .A2(_11659_),
    .B1_N(_11656_),
    .X(_11713_));
 sky130_fd_sc_hd__o21ai_2 _19881_ (.A1(_11655_),
    .A2(_11659_),
    .B1(_11713_),
    .Y(_11714_));
 sky130_fd_sc_hd__xor2_2 _19882_ (.A(_11712_),
    .B(_11714_),
    .X(_11715_));
 sky130_fd_sc_hd__or2_1 _19883_ (.A(_11661_),
    .B(net708),
    .X(_11716_));
 sky130_fd_sc_hd__and3_1 _19884_ (.A(_11543_),
    .B(_11553_),
    .C(_11609_),
    .X(_11717_));
 sky130_fd_sc_hd__mux2_1 _19885_ (.A0(_11544_),
    .A1(_11545_),
    .S(_11609_),
    .X(_11718_));
 sky130_fd_sc_hd__mux2_1 _19886_ (.A0(_11717_),
    .A1(_11718_),
    .S(net604),
    .X(_11719_));
 sky130_fd_sc_hd__nand2_2 _19887_ (.A(net569),
    .B(_11719_),
    .Y(_11720_));
 sky130_fd_sc_hd__and2_1 _19888_ (.A(_11667_),
    .B(net708),
    .X(_11721_));
 sky130_fd_sc_hd__or2_1 _19889_ (.A(_11667_),
    .B(net708),
    .X(_11722_));
 sky130_fd_sc_hd__o211a_1 _19890_ (.A1(_11661_),
    .A2(_11721_),
    .B1(_11722_),
    .C1(net3858),
    .X(_11723_));
 sky130_fd_sc_hd__o21ai_1 _19891_ (.A1(_11667_),
    .A2(_11720_),
    .B1(net708),
    .Y(_11724_));
 sky130_fd_sc_hd__a21bo_1 _19892_ (.A1(_11667_),
    .A2(_11720_),
    .B1_N(_11724_),
    .X(_11725_));
 sky130_fd_sc_hd__a221oi_1 _19893_ (.A1(_11720_),
    .A2(_11721_),
    .B1(_11725_),
    .B2(_11661_),
    .C1(net3858),
    .Y(_11726_));
 sky130_fd_sc_hd__o32a_1 _19894_ (.A1(_11667_),
    .A2(_11716_),
    .A3(_11720_),
    .B1(_11723_),
    .B2(_11726_),
    .X(_11727_));
 sky130_fd_sc_hd__or2_1 _19895_ (.A(_11715_),
    .B(_11727_),
    .X(_11728_));
 sky130_fd_sc_hd__nand2_1 _19896_ (.A(_11715_),
    .B(_11727_),
    .Y(_11729_));
 sky130_fd_sc_hd__and3_1 _19897_ (.A(\cordic0.cos[4] ),
    .B(net2942),
    .C(net1782),
    .X(_11730_));
 sky130_fd_sc_hd__a31o_1 _19898_ (.A1(net1768),
    .A2(_11728_),
    .A3(_11729_),
    .B1(_11730_),
    .X(_00457_));
 sky130_fd_sc_hd__nand3_1 _19899_ (.A(_11667_),
    .B(net708),
    .C(_11715_),
    .Y(_11731_));
 sky130_fd_sc_hd__o31a_1 _19900_ (.A1(_11667_),
    .A2(net708),
    .A3(_11715_),
    .B1(_11731_),
    .X(_11732_));
 sky130_fd_sc_hd__nand2_1 _19901_ (.A(_11661_),
    .B(_11715_),
    .Y(_11733_));
 sky130_fd_sc_hd__o22a_1 _19902_ (.A1(_11661_),
    .A2(_11732_),
    .B1(_11733_),
    .B2(_11670_),
    .X(_11734_));
 sky130_fd_sc_hd__nor2_1 _19903_ (.A(_11720_),
    .B(_11734_),
    .Y(_11735_));
 sky130_fd_sc_hd__nor2_1 _19904_ (.A(net3127),
    .B(net351),
    .Y(_11736_));
 sky130_fd_sc_hd__and2_1 _19905_ (.A(_11712_),
    .B(_11714_),
    .X(_11737_));
 sky130_fd_sc_hd__a21oi_1 _19906_ (.A1(_11661_),
    .A2(net708),
    .B1(_11737_),
    .Y(_11738_));
 sky130_fd_sc_hd__inv_2 _19907_ (.A(_11738_),
    .Y(_11739_));
 sky130_fd_sc_hd__nor2_1 _19908_ (.A(_11712_),
    .B(_11714_),
    .Y(_11740_));
 sky130_fd_sc_hd__o21ba_1 _19909_ (.A1(_11716_),
    .A2(_11737_),
    .B1_N(_11740_),
    .X(_11741_));
 sky130_fd_sc_hd__o21ai_1 _19910_ (.A1(_11667_),
    .A2(_11739_),
    .B1(_11741_),
    .Y(_11742_));
 sky130_fd_sc_hd__a21o_1 _19911_ (.A1(net2097),
    .A2(_11696_),
    .B1(net1412),
    .X(_11743_));
 sky130_fd_sc_hd__o21ai_1 _19912_ (.A1(net2097),
    .A2(_11696_),
    .B1(_11743_),
    .Y(_11744_));
 sky130_fd_sc_hd__mux2_1 _19913_ (.A0(net6117),
    .A1(_11686_),
    .S(net3869),
    .X(_11745_));
 sky130_fd_sc_hd__inv_2 _19914_ (.A(_11329_),
    .Y(_11746_));
 sky130_fd_sc_hd__mux2_1 _19915_ (.A0(_11745_),
    .A1(_11746_),
    .S(_11690_),
    .X(_11747_));
 sky130_fd_sc_hd__o31a_1 _19916_ (.A1(net6110),
    .A2(net3149),
    .A3(_11686_),
    .B1(_11747_),
    .X(_11748_));
 sky130_fd_sc_hd__nor2_1 _19917_ (.A(net3149),
    .B(_11686_),
    .Y(_11749_));
 sky130_fd_sc_hd__and2_1 _19918_ (.A(net3149),
    .B(_11686_),
    .X(_11750_));
 sky130_fd_sc_hd__or4b_1 _19919_ (.A(net3154),
    .B(_11749_),
    .C(_11750_),
    .D_N(_11690_),
    .X(_11751_));
 sky130_fd_sc_hd__or3_1 _19920_ (.A(net6110),
    .B(_11686_),
    .C(_11690_),
    .X(_11752_));
 sky130_fd_sc_hd__o211a_1 _19921_ (.A1(net3916),
    .A2(_11748_),
    .B1(_11751_),
    .C1(_11752_),
    .X(_11753_));
 sky130_fd_sc_hd__nor2_1 _19922_ (.A(net6072),
    .B(_10996_),
    .Y(_11754_));
 sky130_fd_sc_hd__xnor2_2 _19923_ (.A(net6027),
    .B(net3125),
    .Y(_11755_));
 sky130_fd_sc_hd__nand2_1 _19924_ (.A(net6111),
    .B(net3200),
    .Y(_11756_));
 sky130_fd_sc_hd__mux2_1 _19925_ (.A0(_11377_),
    .A1(_11756_),
    .S(net6174),
    .X(_11757_));
 sky130_fd_sc_hd__xnor2_2 _19926_ (.A(net6168),
    .B(net6081),
    .Y(_11758_));
 sky130_fd_sc_hd__xnor2_1 _19927_ (.A(_11757_),
    .B(_11758_),
    .Y(_11759_));
 sky130_fd_sc_hd__xnor2_1 _19928_ (.A(_11755_),
    .B(_11759_),
    .Y(_11760_));
 sky130_fd_sc_hd__nand2_1 _19929_ (.A(net6084),
    .B(net3879),
    .Y(_11761_));
 sky130_fd_sc_hd__nor2_1 _19930_ (.A(net6065),
    .B(net6049),
    .Y(_11762_));
 sky130_fd_sc_hd__a221o_1 _19931_ (.A1(_11761_),
    .A2(_11506_),
    .B1(net3856),
    .B2(net6049),
    .C1(_11762_),
    .X(_11763_));
 sky130_fd_sc_hd__nand2_1 _19932_ (.A(net6007),
    .B(net2498),
    .Y(_11764_));
 sky130_fd_sc_hd__or2_1 _19933_ (.A(net6007),
    .B(net2498),
    .X(_11765_));
 sky130_fd_sc_hd__and2_1 _19934_ (.A(_11764_),
    .B(_11765_),
    .X(_11766_));
 sky130_fd_sc_hd__xor2_1 _19935_ (.A(net1409),
    .B(_11766_),
    .X(_11767_));
 sky130_fd_sc_hd__xnor2_1 _19936_ (.A(net1410),
    .B(_11767_),
    .Y(_11768_));
 sky130_fd_sc_hd__nor2_1 _19937_ (.A(net3137),
    .B(net2096),
    .Y(_11769_));
 sky130_fd_sc_hd__mux2_1 _19938_ (.A0(net6013),
    .A1(_11448_),
    .S(_11769_),
    .X(_11770_));
 sky130_fd_sc_hd__xnor2_1 _19939_ (.A(_11768_),
    .B(net1408),
    .Y(_11771_));
 sky130_fd_sc_hd__xnor2_1 _19940_ (.A(_11744_),
    .B(_11771_),
    .Y(_11772_));
 sky130_fd_sc_hd__a2bb2o_1 _19941_ (.A1_N(net6033),
    .A2_N(net2501),
    .B1(_11699_),
    .B2(net6044),
    .X(_11773_));
 sky130_fd_sc_hd__nand2_1 _19942_ (.A(net6009),
    .B(_11773_),
    .Y(_11774_));
 sky130_fd_sc_hd__a21bo_1 _19943_ (.A1(_11698_),
    .A2(_11703_),
    .B1_N(_11677_),
    .X(_11775_));
 sky130_fd_sc_hd__o21a_1 _19944_ (.A1(_11698_),
    .A2(_11703_),
    .B1(_11775_),
    .X(_11776_));
 sky130_fd_sc_hd__nand2_1 _19945_ (.A(_11774_),
    .B(_11776_),
    .Y(_11777_));
 sky130_fd_sc_hd__or2_1 _19946_ (.A(_11774_),
    .B(_11776_),
    .X(_11778_));
 sky130_fd_sc_hd__nand2_1 _19947_ (.A(_11777_),
    .B(_11778_),
    .Y(_11779_));
 sky130_fd_sc_hd__xnor2_1 _19948_ (.A(_11772_),
    .B(_11779_),
    .Y(_11780_));
 sky130_fd_sc_hd__a21bo_1 _19949_ (.A1(_11674_),
    .A2(_11710_),
    .B1_N(_11708_),
    .X(_11781_));
 sky130_fd_sc_hd__nand2_2 _19950_ (.A(_11780_),
    .B(_11781_),
    .Y(_11782_));
 sky130_fd_sc_hd__or2_1 _19951_ (.A(_11780_),
    .B(_11781_),
    .X(_11783_));
 sky130_fd_sc_hd__nand2_1 _19952_ (.A(_11782_),
    .B(_11783_),
    .Y(_11784_));
 sky130_fd_sc_hd__xnor2_1 _19953_ (.A(net487),
    .B(_11784_),
    .Y(_11785_));
 sky130_fd_sc_hd__xnor2_1 _19954_ (.A(_11736_),
    .B(_11785_),
    .Y(_11786_));
 sky130_fd_sc_hd__a22o_1 _19955_ (.A1(net8997),
    .A2(net1202),
    .B1(_11786_),
    .B2(net1770),
    .X(_00458_));
 sky130_fd_sc_hd__o21a_1 _19956_ (.A1(net1409),
    .A2(_11766_),
    .B1(net1410),
    .X(_11787_));
 sky130_fd_sc_hd__a21oi_4 _19957_ (.A1(net1409),
    .A2(_11766_),
    .B1(_11787_),
    .Y(_11788_));
 sky130_fd_sc_hd__mux2_1 _19958_ (.A0(_11755_),
    .A1(net3199),
    .S(_11758_),
    .X(_11789_));
 sky130_fd_sc_hd__a211o_1 _19959_ (.A1(_11755_),
    .A2(_11758_),
    .B1(net3153),
    .C1(net6107),
    .X(_11790_));
 sky130_fd_sc_hd__o21ai_1 _19960_ (.A1(net6111),
    .A2(_11789_),
    .B1(_11790_),
    .Y(_11791_));
 sky130_fd_sc_hd__or2_1 _19961_ (.A(net3153),
    .B(_11755_),
    .X(_11792_));
 sky130_fd_sc_hd__nand2_1 _19962_ (.A(net3153),
    .B(_11755_),
    .Y(_11793_));
 sky130_fd_sc_hd__nor3_1 _19963_ (.A(net6094),
    .B(_11755_),
    .C(_11758_),
    .Y(_11794_));
 sky130_fd_sc_hd__a41o_1 _19964_ (.A1(net6107),
    .A2(_11758_),
    .A3(_11792_),
    .A4(_11793_),
    .B1(_11794_),
    .X(_11795_));
 sky130_fd_sc_hd__a21oi_1 _19965_ (.A1(net6174),
    .A2(_11791_),
    .B1(_11795_),
    .Y(_11796_));
 sky130_fd_sc_hd__xnor2_2 _19966_ (.A(net4046),
    .B(_11572_),
    .Y(_11797_));
 sky130_fd_sc_hd__or2_1 _19967_ (.A(net6166),
    .B(net6093),
    .X(_11798_));
 sky130_fd_sc_hd__mux2_1 _19968_ (.A0(_10788_),
    .A1(_11798_),
    .S(net6081),
    .X(_11799_));
 sky130_fd_sc_hd__xnor2_2 _19969_ (.A(net6137),
    .B(net6060),
    .Y(_11800_));
 sky130_fd_sc_hd__xnor2_1 _19970_ (.A(_11799_),
    .B(_11800_),
    .Y(_11801_));
 sky130_fd_sc_hd__xnor2_1 _19971_ (.A(_11797_),
    .B(_11801_),
    .Y(_11802_));
 sky130_fd_sc_hd__o22a_1 _19972_ (.A1(net3153),
    .A2(net3199),
    .B1(net6027),
    .B2(net3880),
    .X(_11803_));
 sky130_fd_sc_hd__nor2_1 _19973_ (.A(net6052),
    .B(net6021),
    .Y(_11804_));
 sky130_fd_sc_hd__a211o_1 _19974_ (.A1(net6021),
    .A2(net3125),
    .B1(_11803_),
    .C1(_11804_),
    .X(_11805_));
 sky130_fd_sc_hd__nand2_1 _19975_ (.A(net5999),
    .B(net2092),
    .Y(_11806_));
 sky130_fd_sc_hd__or2_1 _19976_ (.A(net5999),
    .B(net2092),
    .X(_11807_));
 sky130_fd_sc_hd__and2_1 _19977_ (.A(_11806_),
    .B(_11807_),
    .X(_11808_));
 sky130_fd_sc_hd__xor2_1 _19978_ (.A(net2093),
    .B(_11808_),
    .X(_11809_));
 sky130_fd_sc_hd__xnor2_2 _19979_ (.A(net1406),
    .B(_11809_),
    .Y(_11810_));
 sky130_fd_sc_hd__xnor2_1 _19980_ (.A(_11764_),
    .B(_11810_),
    .Y(_11811_));
 sky130_fd_sc_hd__xnor2_2 _19981_ (.A(_11788_),
    .B(_11811_),
    .Y(_11812_));
 sky130_fd_sc_hd__o21a_1 _19982_ (.A1(_11768_),
    .A2(net1408),
    .B1(_11744_),
    .X(_11813_));
 sky130_fd_sc_hd__a21o_1 _19983_ (.A1(_11768_),
    .A2(net1408),
    .B1(_11813_),
    .X(_11814_));
 sky130_fd_sc_hd__nor2_1 _19984_ (.A(net3862),
    .B(net2095),
    .Y(_11815_));
 sky130_fd_sc_hd__nand2_1 _19985_ (.A(_11814_),
    .B(_11815_),
    .Y(_11816_));
 sky130_fd_sc_hd__or2_1 _19986_ (.A(_11814_),
    .B(_11815_),
    .X(_11817_));
 sky130_fd_sc_hd__and2_1 _19987_ (.A(_11816_),
    .B(_11817_),
    .X(_11818_));
 sky130_fd_sc_hd__xnor2_1 _19988_ (.A(_11812_),
    .B(_11818_),
    .Y(_11819_));
 sky130_fd_sc_hd__nor2_1 _19989_ (.A(_11774_),
    .B(_11776_),
    .Y(_11820_));
 sky130_fd_sc_hd__a21o_1 _19990_ (.A1(_11772_),
    .A2(_11777_),
    .B1(_11820_),
    .X(_11821_));
 sky130_fd_sc_hd__nor2_1 _19991_ (.A(_11819_),
    .B(_11821_),
    .Y(_11822_));
 sky130_fd_sc_hd__and2_1 _19992_ (.A(_11819_),
    .B(_11821_),
    .X(_11823_));
 sky130_fd_sc_hd__or2_1 _19993_ (.A(_11822_),
    .B(_11823_),
    .X(_11824_));
 sky130_fd_sc_hd__inv_2 _19994_ (.A(_11783_),
    .Y(_11825_));
 sky130_fd_sc_hd__o21a_1 _19995_ (.A1(_11667_),
    .A2(_11739_),
    .B1(_11741_),
    .X(_11826_));
 sky130_fd_sc_hd__inv_2 _19996_ (.A(_11782_),
    .Y(_11827_));
 sky130_fd_sc_hd__o211ai_1 _19997_ (.A1(_11826_),
    .A2(_11827_),
    .B1(_11783_),
    .C1(net3127),
    .Y(_11828_));
 sky130_fd_sc_hd__o21ai_1 _19998_ (.A1(net350),
    .A2(_11825_),
    .B1(_11782_),
    .Y(_11829_));
 sky130_fd_sc_hd__nor2_1 _19999_ (.A(net351),
    .B(_11782_),
    .Y(_11830_));
 sky130_fd_sc_hd__a211o_1 _20000_ (.A1(_11826_),
    .A2(_11829_),
    .B1(_11830_),
    .C1(net3860),
    .X(_11831_));
 sky130_fd_sc_hd__a32o_1 _20001_ (.A1(net351),
    .A2(net487),
    .A3(_11825_),
    .B1(_11828_),
    .B2(_11831_),
    .X(_11832_));
 sky130_fd_sc_hd__xnor2_1 _20002_ (.A(_11824_),
    .B(_11832_),
    .Y(_11833_));
 sky130_fd_sc_hd__nor2_1 _20003_ (.A(_10344_),
    .B(_11833_),
    .Y(_11834_));
 sky130_fd_sc_hd__a31o_1 _20004_ (.A1(net8975),
    .A2(net2122),
    .A3(net1444),
    .B1(_11834_),
    .X(_00459_));
 sky130_fd_sc_hd__or2_1 _20005_ (.A(_11784_),
    .B(_11824_),
    .X(_11835_));
 sky130_fd_sc_hd__nor2_1 _20006_ (.A(_11782_),
    .B(_11822_),
    .Y(_11836_));
 sky130_fd_sc_hd__a21oi_1 _20007_ (.A1(_11825_),
    .A2(_11824_),
    .B1(_11836_),
    .Y(_11837_));
 sky130_fd_sc_hd__mux2_1 _20008_ (.A0(_11835_),
    .A1(_11837_),
    .S(net487),
    .X(_11838_));
 sky130_fd_sc_hd__inv_2 _20009_ (.A(_11838_),
    .Y(_11839_));
 sky130_fd_sc_hd__a21o_1 _20010_ (.A1(net350),
    .A2(_11839_),
    .B1(net3126),
    .X(_11840_));
 sky130_fd_sc_hd__a2111o_1 _20011_ (.A1(net567),
    .A2(_11716_),
    .B1(_11739_),
    .C1(_11823_),
    .D1(_11836_),
    .X(_11841_));
 sky130_fd_sc_hd__nor2_1 _20012_ (.A(_11823_),
    .B(_11836_),
    .Y(_11842_));
 sky130_fd_sc_hd__o21ai_1 _20013_ (.A1(_11740_),
    .A2(_11835_),
    .B1(_11842_),
    .Y(_11843_));
 sky130_fd_sc_hd__nand2_1 _20014_ (.A(_11841_),
    .B(_11843_),
    .Y(_11844_));
 sky130_fd_sc_hd__nor2_1 _20015_ (.A(_11814_),
    .B(_11815_),
    .Y(_11845_));
 sky130_fd_sc_hd__o21ai_4 _20016_ (.A1(_11812_),
    .A2(_11845_),
    .B1(_11816_),
    .Y(_11846_));
 sky130_fd_sc_hd__a21bo_1 _20017_ (.A1(_11788_),
    .A2(_11810_),
    .B1_N(_11764_),
    .X(_11847_));
 sky130_fd_sc_hd__o21ai_4 _20018_ (.A1(_11788_),
    .A2(_11810_),
    .B1(_11847_),
    .Y(_11848_));
 sky130_fd_sc_hd__o21a_1 _20019_ (.A1(net1406),
    .A2(net2093),
    .B1(_11808_),
    .X(_11849_));
 sky130_fd_sc_hd__a21oi_2 _20020_ (.A1(net1406),
    .A2(net2093),
    .B1(_11849_),
    .Y(_11850_));
 sky130_fd_sc_hd__mux2_1 _20021_ (.A0(net6081),
    .A1(_11797_),
    .S(net3199),
    .X(_11851_));
 sky130_fd_sc_hd__or3_1 _20022_ (.A(net6081),
    .B(net3199),
    .C(_11797_),
    .X(_11852_));
 sky130_fd_sc_hd__o21ai_1 _20023_ (.A1(_11800_),
    .A2(_11851_),
    .B1(_11852_),
    .Y(_11853_));
 sky130_fd_sc_hd__mux2_1 _20024_ (.A0(net3199),
    .A1(_11798_),
    .S(_11797_),
    .X(_11854_));
 sky130_fd_sc_hd__nor3_1 _20025_ (.A(net6081),
    .B(_11797_),
    .C(_11800_),
    .Y(_11855_));
 sky130_fd_sc_hd__a31o_1 _20026_ (.A1(net6081),
    .A2(_11800_),
    .A3(_11854_),
    .B1(_11855_),
    .X(_11856_));
 sky130_fd_sc_hd__a21o_1 _20027_ (.A1(net6168),
    .A2(_11853_),
    .B1(_11856_),
    .X(_11857_));
 sky130_fd_sc_hd__or3_1 _20028_ (.A(net3147),
    .B(net6062),
    .C(net3144),
    .X(_11858_));
 sky130_fd_sc_hd__or3_1 _20029_ (.A(net6134),
    .B(net3132),
    .C(net6077),
    .X(_11859_));
 sky130_fd_sc_hd__nand2_1 _20030_ (.A(net2497),
    .B(_11859_),
    .Y(_11860_));
 sky130_fd_sc_hd__xnor2_2 _20031_ (.A(net6112),
    .B(net6057),
    .Y(_11861_));
 sky130_fd_sc_hd__xor2_1 _20032_ (.A(_11490_),
    .B(_11861_),
    .X(_11862_));
 sky130_fd_sc_hd__xnor2_2 _20033_ (.A(_11860_),
    .B(_11862_),
    .Y(_11863_));
 sky130_fd_sc_hd__nor2_1 _20034_ (.A(net6013),
    .B(net6028),
    .Y(_11864_));
 sky130_fd_sc_hd__a221o_1 _20035_ (.A1(net6028),
    .A2(net3136),
    .B1(_11588_),
    .B2(_11451_),
    .C1(_11864_),
    .X(_11865_));
 sky130_fd_sc_hd__xnor2_1 _20036_ (.A(net3290),
    .B(net2494),
    .Y(_11866_));
 sky130_fd_sc_hd__xnor2_1 _20037_ (.A(_11863_),
    .B(_11866_),
    .Y(_11867_));
 sky130_fd_sc_hd__xnor2_2 _20038_ (.A(net1404),
    .B(_11867_),
    .Y(_11868_));
 sky130_fd_sc_hd__xnor2_1 _20039_ (.A(_11806_),
    .B(_11868_),
    .Y(_11869_));
 sky130_fd_sc_hd__xnor2_2 _20040_ (.A(_11850_),
    .B(_11869_),
    .Y(_11870_));
 sky130_fd_sc_hd__nor2_1 _20041_ (.A(net2581),
    .B(net2498),
    .Y(_11871_));
 sky130_fd_sc_hd__xor2_2 _20042_ (.A(_11870_),
    .B(_11871_),
    .X(_11872_));
 sky130_fd_sc_hd__xnor2_4 _20043_ (.A(_11848_),
    .B(_11872_),
    .Y(_11873_));
 sky130_fd_sc_hd__xnor2_1 _20044_ (.A(_11846_),
    .B(_11873_),
    .Y(_11874_));
 sky130_fd_sc_hd__xnor2_1 _20045_ (.A(_11844_),
    .B(_11874_),
    .Y(_11875_));
 sky130_fd_sc_hd__xnor2_1 _20046_ (.A(_11840_),
    .B(_11875_),
    .Y(_11876_));
 sky130_fd_sc_hd__a22o_1 _20047_ (.A1(net9038),
    .A2(net1202),
    .B1(_11876_),
    .B2(net1771),
    .X(_00460_));
 sky130_fd_sc_hd__o21ba_1 _20048_ (.A1(_11848_),
    .A2(_11870_),
    .B1_N(_11871_),
    .X(_11877_));
 sky130_fd_sc_hd__a21o_1 _20049_ (.A1(_11848_),
    .A2(_11870_),
    .B1(_11877_),
    .X(_11878_));
 sky130_fd_sc_hd__nor2_1 _20050_ (.A(net6058),
    .B(_11490_),
    .Y(_11879_));
 sky130_fd_sc_hd__nor2_1 _20051_ (.A(net6077),
    .B(_11490_),
    .Y(_11880_));
 sky130_fd_sc_hd__a21oi_1 _20052_ (.A1(net3132),
    .A2(net6077),
    .B1(_11880_),
    .Y(_11881_));
 sky130_fd_sc_hd__nor2_1 _20053_ (.A(_11861_),
    .B(_11881_),
    .Y(_11882_));
 sky130_fd_sc_hd__a221o_1 _20054_ (.A1(net3855),
    .A2(_11861_),
    .B1(_11879_),
    .B2(net6077),
    .C1(_11882_),
    .X(_11883_));
 sky130_fd_sc_hd__and2_1 _20055_ (.A(net6077),
    .B(_11490_),
    .X(_11884_));
 sky130_fd_sc_hd__o21a_1 _20056_ (.A1(_11880_),
    .A2(_11884_),
    .B1(net6058),
    .X(_11885_));
 sky130_fd_sc_hd__mux2_1 _20057_ (.A0(_11879_),
    .A1(_11885_),
    .S(_11861_),
    .X(_11886_));
 sky130_fd_sc_hd__a21oi_2 _20058_ (.A1(net6134),
    .A2(_11883_),
    .B1(_11886_),
    .Y(_11887_));
 sky130_fd_sc_hd__and3_1 _20059_ (.A(net6126),
    .B(net6063),
    .C(net3140),
    .X(_11888_));
 sky130_fd_sc_hd__a21o_1 _20060_ (.A1(net3152),
    .A2(net3125),
    .B1(_11888_),
    .X(_11889_));
 sky130_fd_sc_hd__xor2_2 _20061_ (.A(net6095),
    .B(net6021),
    .X(_11890_));
 sky130_fd_sc_hd__xnor2_1 _20062_ (.A(net3294),
    .B(_11890_),
    .Y(_11891_));
 sky130_fd_sc_hd__xor2_1 _20063_ (.A(_11889_),
    .B(_11891_),
    .X(_11892_));
 sky130_fd_sc_hd__o21ai_1 _20064_ (.A1(net3144),
    .A2(_11436_),
    .B1(net6005),
    .Y(_11893_));
 sky130_fd_sc_hd__or2_1 _20065_ (.A(_11892_),
    .B(net2493),
    .X(_11894_));
 sky130_fd_sc_hd__nand2_1 _20066_ (.A(_11892_),
    .B(net2493),
    .Y(_11895_));
 sky130_fd_sc_hd__nand2_1 _20067_ (.A(_11894_),
    .B(_11895_),
    .Y(_11896_));
 sky130_fd_sc_hd__xor2_2 _20068_ (.A(_11887_),
    .B(_11896_),
    .X(_11897_));
 sky130_fd_sc_hd__nor2_1 _20069_ (.A(_11863_),
    .B(net2494),
    .Y(_11898_));
 sky130_fd_sc_hd__nand2_1 _20070_ (.A(_11863_),
    .B(net2494),
    .Y(_11899_));
 sky130_fd_sc_hd__o21a_1 _20071_ (.A1(net1404),
    .A2(_11898_),
    .B1(_11899_),
    .X(_11900_));
 sky130_fd_sc_hd__nor2_1 _20072_ (.A(net1404),
    .B(_11899_),
    .Y(_11901_));
 sky130_fd_sc_hd__a22o_1 _20073_ (.A1(net1404),
    .A2(_11898_),
    .B1(_11901_),
    .B2(net6002),
    .X(_11902_));
 sky130_fd_sc_hd__a21o_1 _20074_ (.A1(net2582),
    .A2(_11900_),
    .B1(_11902_),
    .X(_11903_));
 sky130_fd_sc_hd__xnor2_2 _20075_ (.A(_11897_),
    .B(_11903_),
    .Y(_11904_));
 sky130_fd_sc_hd__a21bo_1 _20076_ (.A1(_11850_),
    .A2(_11868_),
    .B1_N(_11806_),
    .X(_11905_));
 sky130_fd_sc_hd__o21a_1 _20077_ (.A1(_11850_),
    .A2(_11868_),
    .B1(_11905_),
    .X(_11906_));
 sky130_fd_sc_hd__nor2_1 _20078_ (.A(net2581),
    .B(net2092),
    .Y(_11907_));
 sky130_fd_sc_hd__xnor2_1 _20079_ (.A(_11906_),
    .B(_11907_),
    .Y(_11908_));
 sky130_fd_sc_hd__xor2_2 _20080_ (.A(_11904_),
    .B(_11908_),
    .X(_11909_));
 sky130_fd_sc_hd__nand2_1 _20081_ (.A(_11878_),
    .B(_11909_),
    .Y(_11910_));
 sky130_fd_sc_hd__nor2_1 _20082_ (.A(_11878_),
    .B(_11909_),
    .Y(_11911_));
 sky130_fd_sc_hd__inv_2 _20083_ (.A(_11911_),
    .Y(_11912_));
 sky130_fd_sc_hd__nand2_1 _20084_ (.A(_11910_),
    .B(_11912_),
    .Y(_11913_));
 sky130_fd_sc_hd__nand2_1 _20085_ (.A(net350),
    .B(_11839_),
    .Y(_11914_));
 sky130_fd_sc_hd__nand2_1 _20086_ (.A(_11844_),
    .B(_11873_),
    .Y(_11915_));
 sky130_fd_sc_hd__nor2_1 _20087_ (.A(_11844_),
    .B(_11873_),
    .Y(_11916_));
 sky130_fd_sc_hd__a21o_1 _20088_ (.A1(_11914_),
    .A2(_11915_),
    .B1(_11916_),
    .X(_11917_));
 sky130_fd_sc_hd__a221oi_1 _20089_ (.A1(_11914_),
    .A2(_11916_),
    .B1(_11917_),
    .B2(_11846_),
    .C1(net3861),
    .Y(_11918_));
 sky130_fd_sc_hd__inv_2 _20090_ (.A(_11873_),
    .Y(_11919_));
 sky130_fd_sc_hd__a31o_1 _20091_ (.A1(_11841_),
    .A2(_11843_),
    .A3(_11919_),
    .B1(_11846_),
    .X(_11920_));
 sky130_fd_sc_hd__and3_1 _20092_ (.A(net3861),
    .B(_11915_),
    .C(_11920_),
    .X(_11921_));
 sky130_fd_sc_hd__o32a_1 _20093_ (.A1(_11914_),
    .A2(_11846_),
    .A3(_11915_),
    .B1(_11918_),
    .B2(_11921_),
    .X(_11922_));
 sky130_fd_sc_hd__or2_1 _20094_ (.A(_11913_),
    .B(_11922_),
    .X(_11923_));
 sky130_fd_sc_hd__nand2_1 _20095_ (.A(_11913_),
    .B(_11922_),
    .Y(_11924_));
 sky130_fd_sc_hd__a21oi_1 _20096_ (.A1(_11923_),
    .A2(_11924_),
    .B1(net1438),
    .Y(_11925_));
 sky130_fd_sc_hd__a31o_1 _20097_ (.A1(net9025),
    .A2(net2124),
    .A3(net1446),
    .B1(_11925_),
    .X(_00461_));
 sky130_fd_sc_hd__o21ai_1 _20098_ (.A1(net487),
    .A2(_11835_),
    .B1(_11873_),
    .Y(_11926_));
 sky130_fd_sc_hd__a31oi_2 _20099_ (.A1(_11910_),
    .A2(_11920_),
    .A3(net420),
    .B1(_11911_),
    .Y(_11927_));
 sky130_fd_sc_hd__inv_2 _20100_ (.A(_11909_),
    .Y(_11928_));
 sky130_fd_sc_hd__nand2_1 _20101_ (.A(_11928_),
    .B(_11920_),
    .Y(_11929_));
 sky130_fd_sc_hd__or2_1 _20102_ (.A(_11911_),
    .B(net420),
    .X(_11930_));
 sky130_fd_sc_hd__o21ai_1 _20103_ (.A1(_11928_),
    .A2(_11920_),
    .B1(_11930_),
    .Y(_11931_));
 sky130_fd_sc_hd__a21oi_1 _20104_ (.A1(_11878_),
    .A2(_11929_),
    .B1(_11931_),
    .Y(_11932_));
 sky130_fd_sc_hd__a21o_1 _20105_ (.A1(_11906_),
    .A2(_11904_),
    .B1(_11907_),
    .X(_11933_));
 sky130_fd_sc_hd__o21a_2 _20106_ (.A1(_11906_),
    .A2(_11904_),
    .B1(_11933_),
    .X(_11934_));
 sky130_fd_sc_hd__mux2_1 _20107_ (.A0(net6052),
    .A1(net6000),
    .S(_11890_),
    .X(_11935_));
 sky130_fd_sc_hd__o211a_1 _20108_ (.A1(net6001),
    .A2(_11890_),
    .B1(net6063),
    .C1(net3140),
    .X(_11936_));
 sky130_fd_sc_hd__a21o_1 _20109_ (.A1(net3134),
    .A2(_11935_),
    .B1(_11936_),
    .X(_11937_));
 sky130_fd_sc_hd__xor2_1 _20110_ (.A(net6063),
    .B(net6005),
    .X(_11938_));
 sky130_fd_sc_hd__and2_1 _20111_ (.A(net6052),
    .B(_11938_),
    .X(_11939_));
 sky130_fd_sc_hd__mux2_1 _20112_ (.A0(_11939_),
    .A1(_11447_),
    .S(_11890_),
    .X(_11940_));
 sky130_fd_sc_hd__a21oi_2 _20113_ (.A1(net6112),
    .A2(_11937_),
    .B1(_11940_),
    .Y(_11941_));
 sky130_fd_sc_hd__or2_1 _20114_ (.A(net6107),
    .B(net6042),
    .X(_11942_));
 sky130_fd_sc_hd__mux2_1 _20115_ (.A0(_11292_),
    .A1(_11942_),
    .S(net6027),
    .X(_11943_));
 sky130_fd_sc_hd__xnor2_1 _20116_ (.A(net6079),
    .B(_11943_),
    .Y(_11944_));
 sky130_fd_sc_hd__nand2_1 _20117_ (.A(net6006),
    .B(_11648_),
    .Y(_11945_));
 sky130_fd_sc_hd__or2_1 _20118_ (.A(_11944_),
    .B(_11945_),
    .X(_11946_));
 sky130_fd_sc_hd__nand2_1 _20119_ (.A(_11944_),
    .B(_11945_),
    .Y(_11947_));
 sky130_fd_sc_hd__and2_1 _20120_ (.A(_11946_),
    .B(_11947_),
    .X(_11948_));
 sky130_fd_sc_hd__xnor2_2 _20121_ (.A(_11941_),
    .B(_11948_),
    .Y(_11949_));
 sky130_fd_sc_hd__mux2_1 _20122_ (.A0(_11895_),
    .A1(_11894_),
    .S(_11887_),
    .X(_11950_));
 sky130_fd_sc_hd__xnor2_1 _20123_ (.A(_11949_),
    .B(_11950_),
    .Y(_11951_));
 sky130_fd_sc_hd__or2_1 _20124_ (.A(net2582),
    .B(_11901_),
    .X(_11952_));
 sky130_fd_sc_hd__a2bb2o_1 _20125_ (.A1_N(net5999),
    .A2_N(_11900_),
    .B1(_11952_),
    .B2(_11897_),
    .X(_11953_));
 sky130_fd_sc_hd__nor2_1 _20126_ (.A(net1055),
    .B(_11953_),
    .Y(_11954_));
 sky130_fd_sc_hd__and2_1 _20127_ (.A(net1055),
    .B(_11953_),
    .X(_11955_));
 sky130_fd_sc_hd__nor2_1 _20128_ (.A(_11954_),
    .B(_11955_),
    .Y(_11956_));
 sky130_fd_sc_hd__xnor2_1 _20129_ (.A(_11934_),
    .B(_11956_),
    .Y(_11957_));
 sky130_fd_sc_hd__mux2_1 _20130_ (.A0(_11927_),
    .A1(_11932_),
    .S(_11957_),
    .X(_11958_));
 sky130_fd_sc_hd__or2_1 _20131_ (.A(_11844_),
    .B(_11873_),
    .X(_11959_));
 sky130_fd_sc_hd__mux2_1 _20132_ (.A0(_11959_),
    .A1(_11915_),
    .S(_11913_),
    .X(_11960_));
 sky130_fd_sc_hd__or3b_1 _20133_ (.A(_11873_),
    .B(_11913_),
    .C_N(_11846_),
    .X(_11961_));
 sky130_fd_sc_hd__o21a_1 _20134_ (.A1(_11846_),
    .A2(_11960_),
    .B1(_11961_),
    .X(_11962_));
 sky130_fd_sc_hd__or2_1 _20135_ (.A(_11914_),
    .B(_11962_),
    .X(_11963_));
 sky130_fd_sc_hd__and2b_1 _20136_ (.A_N(net3126),
    .B(_11963_),
    .X(_11964_));
 sky130_fd_sc_hd__xnor2_1 _20137_ (.A(net274),
    .B(_11964_),
    .Y(_11965_));
 sky130_fd_sc_hd__nor2_1 _20138_ (.A(net1439),
    .B(_11965_),
    .Y(_11966_));
 sky130_fd_sc_hd__a31o_1 _20139_ (.A1(net8972),
    .A2(net2124),
    .A3(net1445),
    .B1(_11966_),
    .X(_00462_));
 sky130_fd_sc_hd__nor2_1 _20140_ (.A(net274),
    .B(_11963_),
    .Y(_11967_));
 sky130_fd_sc_hd__xnor2_1 _20141_ (.A(_11889_),
    .B(_11891_),
    .Y(_11968_));
 sky130_fd_sc_hd__a21o_1 _20142_ (.A1(_11968_),
    .A2(_11949_),
    .B1(net2493),
    .X(_11969_));
 sky130_fd_sc_hd__o21a_1 _20143_ (.A1(_11968_),
    .A2(_11949_),
    .B1(net2493),
    .X(_11970_));
 sky130_fd_sc_hd__a21oi_1 _20144_ (.A1(_11887_),
    .A2(_11969_),
    .B1(_11970_),
    .Y(_11971_));
 sky130_fd_sc_hd__nand2_1 _20145_ (.A(net3137),
    .B(_11292_),
    .Y(_11972_));
 sky130_fd_sc_hd__a22o_1 _20146_ (.A1(net6027),
    .A2(_11942_),
    .B1(_11972_),
    .B2(net6078),
    .X(_11973_));
 sky130_fd_sc_hd__xnor2_1 _20147_ (.A(_11938_),
    .B(_11973_),
    .Y(_11974_));
 sky130_fd_sc_hd__mux2_1 _20148_ (.A0(_11947_),
    .A1(_11946_),
    .S(_11941_),
    .X(_11975_));
 sky130_fd_sc_hd__xor2_1 _20149_ (.A(_11974_),
    .B(_11975_),
    .X(_11976_));
 sky130_fd_sc_hd__a22oi_2 _20150_ (.A1(net6079),
    .A2(_11491_),
    .B1(_11971_),
    .B2(_11976_),
    .Y(_11977_));
 sky130_fd_sc_hd__o21a_1 _20151_ (.A1(_11971_),
    .A2(_11976_),
    .B1(_11977_),
    .X(_11978_));
 sky130_fd_sc_hd__nand2_1 _20152_ (.A(net1055),
    .B(_11953_),
    .Y(_11979_));
 sky130_fd_sc_hd__a21o_1 _20153_ (.A1(_11934_),
    .A2(_11979_),
    .B1(_11954_),
    .X(_11980_));
 sky130_fd_sc_hd__or2_1 _20154_ (.A(_11911_),
    .B(_11920_),
    .X(_11981_));
 sky130_fd_sc_hd__or3_1 _20155_ (.A(_11927_),
    .B(net1055),
    .C(_11953_),
    .X(_11982_));
 sky130_fd_sc_hd__mux2_1 _20156_ (.A0(_11979_),
    .A1(_11982_),
    .S(_11934_),
    .X(_11983_));
 sky130_fd_sc_hd__and2_1 _20157_ (.A(_11910_),
    .B(_11930_),
    .X(_11984_));
 sky130_fd_sc_hd__or2_1 _20158_ (.A(_11984_),
    .B(_11980_),
    .X(_11985_));
 sky130_fd_sc_hd__o211a_1 _20159_ (.A1(_11980_),
    .A2(_11981_),
    .B1(_11983_),
    .C1(_11985_),
    .X(_11986_));
 sky130_fd_sc_hd__xnor2_1 _20160_ (.A(net868),
    .B(_11986_),
    .Y(_11987_));
 sky130_fd_sc_hd__or3b_1 _20161_ (.A(net3126),
    .B(_11967_),
    .C_N(net244),
    .X(_11988_));
 sky130_fd_sc_hd__o21bai_1 _20162_ (.A1(net3126),
    .A2(_11967_),
    .B1_N(net244),
    .Y(_11989_));
 sky130_fd_sc_hd__a21oi_1 _20163_ (.A1(_11988_),
    .A2(_11989_),
    .B1(net1439),
    .Y(_11990_));
 sky130_fd_sc_hd__a31o_1 _20164_ (.A1(net9006),
    .A2(net2122),
    .A3(net1444),
    .B1(_11990_),
    .X(_00463_));
 sky130_fd_sc_hd__inv_2 _20165_ (.A(_11934_),
    .Y(_11991_));
 sky130_fd_sc_hd__a2bb2o_1 _20166_ (.A1_N(_11927_),
    .A2_N(_11991_),
    .B1(_11979_),
    .B2(net868),
    .X(_11992_));
 sky130_fd_sc_hd__a21o_1 _20167_ (.A1(_11927_),
    .A2(_11955_),
    .B1(_11991_),
    .X(_11993_));
 sky130_fd_sc_hd__o21ai_1 _20168_ (.A1(_11927_),
    .A2(_11955_),
    .B1(_11993_),
    .Y(_11994_));
 sky130_fd_sc_hd__a22oi_2 _20169_ (.A1(_11954_),
    .A2(_11992_),
    .B1(_11994_),
    .B2(net868),
    .Y(_11995_));
 sky130_fd_sc_hd__nor2_1 _20170_ (.A(net6100),
    .B(net6042),
    .Y(_11996_));
 sky130_fd_sc_hd__a32o_1 _20171_ (.A1(net6004),
    .A2(net3137),
    .A3(_11754_),
    .B1(_11996_),
    .B2(net6072),
    .X(_11997_));
 sky130_fd_sc_hd__nor2_1 _20172_ (.A(net6078),
    .B(_11997_),
    .Y(_11998_));
 sky130_fd_sc_hd__o221a_1 _20173_ (.A1(_11348_),
    .A2(_11588_),
    .B1(net3128),
    .B2(net6067),
    .C1(net6088),
    .X(_11999_));
 sky130_fd_sc_hd__and3_1 _20174_ (.A(net6059),
    .B(net2580),
    .C(net6024),
    .X(_12000_));
 sky130_fd_sc_hd__or4_1 _20175_ (.A(net6059),
    .B(net6100),
    .C(net2580),
    .D(net6024),
    .X(_12001_));
 sky130_fd_sc_hd__and3b_1 _20176_ (.A_N(_12000_),
    .B(_12001_),
    .C(net6042),
    .X(_12002_));
 sky130_fd_sc_hd__o211a_1 _20177_ (.A1(net3200),
    .A2(net3137),
    .B1(net6013),
    .C1(_11489_),
    .X(_12003_));
 sky130_fd_sc_hd__o21a_1 _20178_ (.A1(_12000_),
    .A2(_12003_),
    .B1(_11410_),
    .X(_12004_));
 sky130_fd_sc_hd__o22a_1 _20179_ (.A1(_11998_),
    .A2(_11999_),
    .B1(_12002_),
    .B2(_12004_),
    .X(_12005_));
 sky130_fd_sc_hd__or2b_1 _20180_ (.A(_11944_),
    .B_N(_11974_),
    .X(_12006_));
 sky130_fd_sc_hd__or2b_1 _20181_ (.A(_11974_),
    .B_N(_11944_),
    .X(_12007_));
 sky130_fd_sc_hd__a21oi_1 _20182_ (.A1(net2580),
    .A2(_12007_),
    .B1(_11941_),
    .Y(_12008_));
 sky130_fd_sc_hd__a21o_1 _20183_ (.A1(net6004),
    .A2(_12006_),
    .B1(_12008_),
    .X(_12009_));
 sky130_fd_sc_hd__a2bb2o_1 _20184_ (.A1_N(net2580),
    .A2_N(_11648_),
    .B1(_12005_),
    .B2(_12009_),
    .X(_12010_));
 sky130_fd_sc_hd__a311o_1 _20185_ (.A1(net6004),
    .A2(_11648_),
    .A3(_12006_),
    .B1(_12008_),
    .C1(_12005_),
    .X(_12011_));
 sky130_fd_sc_hd__or2b_1 _20186_ (.A(_12010_),
    .B_N(_12011_),
    .X(_12012_));
 sky130_fd_sc_hd__xor2_1 _20187_ (.A(net952),
    .B(net867),
    .X(_12013_));
 sky130_fd_sc_hd__xnor2_1 _20188_ (.A(_11995_),
    .B(_12013_),
    .Y(_12014_));
 sky130_fd_sc_hd__a21o_1 _20189_ (.A1(net244),
    .A2(_11967_),
    .B1(net3126),
    .X(_12015_));
 sky130_fd_sc_hd__xnor2_1 _20190_ (.A(net243),
    .B(_12015_),
    .Y(_12016_));
 sky130_fd_sc_hd__and3_1 _20191_ (.A(\cordic0.cos[11] ),
    .B(net2122),
    .C(net1784),
    .X(_12017_));
 sky130_fd_sc_hd__a21o_1 _20192_ (.A1(net1770),
    .A2(_12016_),
    .B1(_12017_),
    .X(_00464_));
 sky130_fd_sc_hd__and3b_1 _20193_ (.A_N(net952),
    .B(_11954_),
    .C(_11934_),
    .X(_12018_));
 sky130_fd_sc_hd__a21oi_1 _20194_ (.A1(net952),
    .A2(_11995_),
    .B1(net867),
    .Y(_12019_));
 sky130_fd_sc_hd__a31o_1 _20195_ (.A1(_11984_),
    .A2(_11981_),
    .A3(_12018_),
    .B1(_12019_),
    .X(_12020_));
 sky130_fd_sc_hd__a21oi_1 _20196_ (.A1(net3145),
    .A2(_11996_),
    .B1(net2580),
    .Y(_12021_));
 sky130_fd_sc_hd__o221a_1 _20197_ (.A1(net6042),
    .A2(net6000),
    .B1(_12021_),
    .B2(net6063),
    .C1(net6024),
    .X(_12022_));
 sky130_fd_sc_hd__a31o_1 _20198_ (.A1(net6090),
    .A2(net6096),
    .A3(net6042),
    .B1(net6000),
    .X(_12023_));
 sky130_fd_sc_hd__a221o_1 _20199_ (.A1(net6042),
    .A2(net6000),
    .B1(_12023_),
    .B2(net6063),
    .C1(net6034),
    .X(_12024_));
 sky130_fd_sc_hd__and2b_1 _20200_ (.A_N(_12022_),
    .B(_12024_),
    .X(_12025_));
 sky130_fd_sc_hd__xnor2_1 _20201_ (.A(_12010_),
    .B(_12025_),
    .Y(_12026_));
 sky130_fd_sc_hd__xnor2_1 _20202_ (.A(_12020_),
    .B(net866),
    .Y(_12027_));
 sky130_fd_sc_hd__nand2_1 _20203_ (.A(net244),
    .B(_11967_),
    .Y(_12028_));
 sky130_fd_sc_hd__o21ba_1 _20204_ (.A1(net243),
    .A2(_12028_),
    .B1_N(net3126),
    .X(_12029_));
 sky130_fd_sc_hd__xnor2_1 _20205_ (.A(net179),
    .B(_12029_),
    .Y(_12030_));
 sky130_fd_sc_hd__nor2_1 _20206_ (.A(net1785),
    .B(_12030_),
    .Y(_12031_));
 sky130_fd_sc_hd__a31o_1 _20207_ (.A1(net9046),
    .A2(net2123),
    .A3(net1445),
    .B1(_12031_),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _20208_ (.A0(_12029_),
    .A1(net3126),
    .S(net179),
    .X(_12032_));
 sky130_fd_sc_hd__and3_1 _20209_ (.A(\cordic0.cos[13] ),
    .B(net2123),
    .C(net1784),
    .X(_12033_));
 sky130_fd_sc_hd__a21o_1 _20210_ (.A1(net1770),
    .A2(_12032_),
    .B1(_12033_),
    .X(_00466_));
 sky130_fd_sc_hd__nor2_1 _20211_ (.A(net8120),
    .B(net8119),
    .Y(_12034_));
 sky130_fd_sc_hd__xnor2_1 _20212_ (.A(net8953),
    .B(_12034_),
    .Y(_12035_));
 sky130_fd_sc_hd__mux2_1 _20213_ (.A0(_12035_),
    .A1(\cordic0.slte0.opB[2] ),
    .S(net2937),
    .X(_12036_));
 sky130_fd_sc_hd__clkbuf_1 _20214_ (.A(_12036_),
    .X(_00467_));
 sky130_fd_sc_hd__a21oi_1 _20215_ (.A1(net8953),
    .A2(net8119),
    .B1(net8120),
    .Y(_12037_));
 sky130_fd_sc_hd__xnor2_1 _20216_ (.A(net8),
    .B(_12037_),
    .Y(_12038_));
 sky130_fd_sc_hd__mux2_1 _20217_ (.A0(_12038_),
    .A1(\cordic0.slte0.opB[3] ),
    .S(net2937),
    .X(_12039_));
 sky130_fd_sc_hd__clkbuf_1 _20218_ (.A(_12039_),
    .X(_00468_));
 sky130_fd_sc_hd__a31o_1 _20219_ (.A1(net8953),
    .A2(net8119),
    .A3(net8),
    .B1(net8120),
    .X(_12040_));
 sky130_fd_sc_hd__xor2_1 _20220_ (.A(net8100),
    .B(_12040_),
    .X(_12041_));
 sky130_fd_sc_hd__mux2_1 _20221_ (.A0(_12041_),
    .A1(\cordic0.slte0.opB[4] ),
    .S(net2937),
    .X(_12042_));
 sky130_fd_sc_hd__clkbuf_1 _20222_ (.A(_12042_),
    .X(_00469_));
 sky130_fd_sc_hd__and4_1 _20223_ (.A(net8953),
    .B(net8119),
    .C(net8),
    .D(net8100),
    .X(_12043_));
 sky130_fd_sc_hd__nor2_1 _20224_ (.A(net8120),
    .B(_12043_),
    .Y(_12044_));
 sky130_fd_sc_hd__xnor2_1 _20225_ (.A(net10),
    .B(_12044_),
    .Y(_12045_));
 sky130_fd_sc_hd__mux2_1 _20226_ (.A0(_12045_),
    .A1(\cordic0.slte0.opB[5] ),
    .S(net2936),
    .X(_12046_));
 sky130_fd_sc_hd__clkbuf_1 _20227_ (.A(_12046_),
    .X(_00470_));
 sky130_fd_sc_hd__a21oi_1 _20228_ (.A1(net10),
    .A2(_12043_),
    .B1(net8122),
    .Y(_12047_));
 sky130_fd_sc_hd__xnor2_1 _20229_ (.A(net11),
    .B(_12047_),
    .Y(_12048_));
 sky130_fd_sc_hd__mux2_1 _20230_ (.A0(_12048_),
    .A1(net6415),
    .S(net2936),
    .X(_12049_));
 sky130_fd_sc_hd__clkbuf_1 _20231_ (.A(_12049_),
    .X(_00471_));
 sky130_fd_sc_hd__and3_1 _20232_ (.A(net10),
    .B(net11),
    .C(_12043_),
    .X(_12050_));
 sky130_fd_sc_hd__nor2_1 _20233_ (.A(net8122),
    .B(_12050_),
    .Y(_12051_));
 sky130_fd_sc_hd__xnor2_1 _20234_ (.A(net12),
    .B(_12051_),
    .Y(_12052_));
 sky130_fd_sc_hd__mux2_1 _20235_ (.A0(_12052_),
    .A1(net6412),
    .S(net2936),
    .X(_12053_));
 sky130_fd_sc_hd__clkbuf_1 _20236_ (.A(_12053_),
    .X(_00472_));
 sky130_fd_sc_hd__and2_1 _20237_ (.A(net12),
    .B(_12050_),
    .X(_12054_));
 sky130_fd_sc_hd__nor2_1 _20238_ (.A(net8122),
    .B(_12054_),
    .Y(_12055_));
 sky130_fd_sc_hd__xnor2_1 _20239_ (.A(net13),
    .B(_12055_),
    .Y(_12056_));
 sky130_fd_sc_hd__mux2_1 _20240_ (.A0(_12056_),
    .A1(\cordic0.slte0.opB[8] ),
    .S(net2936),
    .X(_12057_));
 sky130_fd_sc_hd__clkbuf_1 _20241_ (.A(_12057_),
    .X(_00473_));
 sky130_fd_sc_hd__a31o_1 _20242_ (.A1(net12),
    .A2(net13),
    .A3(_12050_),
    .B1(net8122),
    .X(_12058_));
 sky130_fd_sc_hd__xor2_1 _20243_ (.A(net14),
    .B(_12058_),
    .X(_12059_));
 sky130_fd_sc_hd__mux2_1 _20244_ (.A0(_12059_),
    .A1(\cordic0.slte0.opB[9] ),
    .S(net2532),
    .X(_12060_));
 sky130_fd_sc_hd__clkbuf_1 _20245_ (.A(_12060_),
    .X(_00474_));
 sky130_fd_sc_hd__and3_1 _20246_ (.A(net13),
    .B(net14),
    .C(_12054_),
    .X(_12061_));
 sky130_fd_sc_hd__nor2_1 _20247_ (.A(net8121),
    .B(_12061_),
    .Y(_12062_));
 sky130_fd_sc_hd__xnor2_1 _20248_ (.A(net15),
    .B(_12062_),
    .Y(_12063_));
 sky130_fd_sc_hd__mux2_1 _20249_ (.A0(_12063_),
    .A1(\cordic0.slte0.opB[10] ),
    .S(net2532),
    .X(_12064_));
 sky130_fd_sc_hd__clkbuf_1 _20250_ (.A(_12064_),
    .X(_00475_));
 sky130_fd_sc_hd__and2_1 _20251_ (.A(net15),
    .B(_12061_),
    .X(_12065_));
 sky130_fd_sc_hd__nor2_1 _20252_ (.A(net8121),
    .B(_12065_),
    .Y(_12066_));
 sky130_fd_sc_hd__xnor2_1 _20253_ (.A(net16),
    .B(_12066_),
    .Y(_12067_));
 sky130_fd_sc_hd__mux2_1 _20254_ (.A0(_12067_),
    .A1(\cordic0.slte0.opB[11] ),
    .S(net2531),
    .X(_12068_));
 sky130_fd_sc_hd__clkbuf_1 _20255_ (.A(_12068_),
    .X(_00476_));
 sky130_fd_sc_hd__a31o_1 _20256_ (.A1(net15),
    .A2(net16),
    .A3(_12061_),
    .B1(net8121),
    .X(_12069_));
 sky130_fd_sc_hd__xor2_1 _20257_ (.A(net2),
    .B(_12069_),
    .X(_12070_));
 sky130_fd_sc_hd__mux2_1 _20258_ (.A0(_12070_),
    .A1(\cordic0.slte0.opB[12] ),
    .S(net2531),
    .X(_12071_));
 sky130_fd_sc_hd__clkbuf_1 _20259_ (.A(_12071_),
    .X(_00477_));
 sky130_fd_sc_hd__and3_1 _20260_ (.A(net16),
    .B(net2),
    .C(_12065_),
    .X(_12072_));
 sky130_fd_sc_hd__nor2_1 _20261_ (.A(net8121),
    .B(_12072_),
    .Y(_12073_));
 sky130_fd_sc_hd__xnor2_1 _20262_ (.A(net3),
    .B(_12073_),
    .Y(_12074_));
 sky130_fd_sc_hd__mux2_1 _20263_ (.A0(_12074_),
    .A1(\cordic0.slte0.opB[13] ),
    .S(net2531),
    .X(_12075_));
 sky130_fd_sc_hd__clkbuf_1 _20264_ (.A(_12075_),
    .X(_00478_));
 sky130_fd_sc_hd__a21oi_1 _20265_ (.A1(net3),
    .A2(_12072_),
    .B1(net8121),
    .Y(_12076_));
 sky130_fd_sc_hd__xnor2_1 _20266_ (.A(net4),
    .B(_12076_),
    .Y(_12077_));
 sky130_fd_sc_hd__mux2_1 _20267_ (.A0(_12077_),
    .A1(\cordic0.slte0.opB[14] ),
    .S(net2531),
    .X(_12078_));
 sky130_fd_sc_hd__clkbuf_1 _20268_ (.A(_12078_),
    .X(_00479_));
 sky130_fd_sc_hd__a31o_1 _20269_ (.A1(net3),
    .A2(net4),
    .A3(_12072_),
    .B1(net8121),
    .X(_12079_));
 sky130_fd_sc_hd__xor2_1 _20270_ (.A(net5),
    .B(_12079_),
    .X(_12080_));
 sky130_fd_sc_hd__mux2_1 _20271_ (.A0(_12080_),
    .A1(\cordic0.slte0.opB[15] ),
    .S(net2531),
    .X(_12081_));
 sky130_fd_sc_hd__clkbuf_1 _20272_ (.A(_12081_),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _20273_ (.A0(net8122),
    .A1(\cordic0.domain[0] ),
    .S(net2533),
    .X(_12082_));
 sky130_fd_sc_hd__clkbuf_1 _20274_ (.A(_12082_),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _20275_ (.A0(net7),
    .A1(\cordic0.domain[1] ),
    .S(net2533),
    .X(_12083_));
 sky130_fd_sc_hd__clkbuf_1 _20276_ (.A(_12083_),
    .X(_00482_));
 sky130_fd_sc_hd__nor2_1 _20277_ (.A(net4041),
    .B(net6472),
    .Y(_12084_));
 sky130_fd_sc_hd__or2_1 _20278_ (.A(net6516),
    .B(_12084_),
    .X(_12085_));
 sky130_fd_sc_hd__o311a_1 _20279_ (.A1(net3314),
    .A2(net6476),
    .A3(net2604),
    .B1(_12085_),
    .C1(net2608),
    .X(_12086_));
 sky130_fd_sc_hd__o21ai_1 _20280_ (.A1(net1835),
    .A2(net2091),
    .B1(net8055),
    .Y(_12087_));
 sky130_fd_sc_hd__nor2_1 _20281_ (.A(\cordic0.slte0.opA[0] ),
    .B(net1556),
    .Y(_12088_));
 sky130_fd_sc_hd__a22o_1 _20282_ (.A1(net9208),
    .A2(_12087_),
    .B1(_12088_),
    .B2(net2091),
    .X(_00483_));
 sky130_fd_sc_hd__nand2_1 _20283_ (.A(\cordic0.slte0.opA[0] ),
    .B(net2091),
    .Y(_12089_));
 sky130_fd_sc_hd__nor2_1 _20284_ (.A(net6499),
    .B(net6468),
    .Y(_12090_));
 sky130_fd_sc_hd__mux2_1 _20285_ (.A0(net6499),
    .A1(_12090_),
    .S(net1824),
    .X(_12091_));
 sky130_fd_sc_hd__nor2_1 _20286_ (.A(_09032_),
    .B(net1485),
    .Y(_12092_));
 sky130_fd_sc_hd__or2_1 _20287_ (.A(net6516),
    .B(net6468),
    .X(_12093_));
 sky130_fd_sc_hd__o221a_1 _20288_ (.A1(net3314),
    .A2(_12091_),
    .B1(_12092_),
    .B2(_12093_),
    .C1(net6479),
    .X(_12094_));
 sky130_fd_sc_hd__or2_1 _20289_ (.A(net4041),
    .B(_06504_),
    .X(_12095_));
 sky130_fd_sc_hd__inv_2 _20290_ (.A(_12095_),
    .Y(_12096_));
 sky130_fd_sc_hd__a21oi_1 _20291_ (.A1(net1482),
    .A2(_12096_),
    .B1(net2604),
    .Y(_12097_));
 sky130_fd_sc_hd__nand2_2 _20292_ (.A(net6468),
    .B(net1486),
    .Y(_12098_));
 sky130_fd_sc_hd__o22ai_1 _20293_ (.A1(net6516),
    .A2(_12097_),
    .B1(_12098_),
    .B2(net6494),
    .Y(_12099_));
 sky130_fd_sc_hd__o21ai_1 _20294_ (.A1(_12094_),
    .A2(_12099_),
    .B1(net2608),
    .Y(_12100_));
 sky130_fd_sc_hd__nor2_1 _20295_ (.A(_12089_),
    .B(_12100_),
    .Y(_12101_));
 sky130_fd_sc_hd__nand2_1 _20296_ (.A(_12089_),
    .B(_12100_),
    .Y(_12102_));
 sky130_fd_sc_hd__or2b_1 _20297_ (.A(_12101_),
    .B_N(_12102_),
    .X(_12103_));
 sky130_fd_sc_hd__a21o_1 _20298_ (.A1(net1471),
    .A2(_12103_),
    .B1(net3317),
    .X(_12104_));
 sky130_fd_sc_hd__or3_1 _20299_ (.A(\cordic0.slte0.opA[1] ),
    .B(net2281),
    .C(_12103_),
    .X(_12105_));
 sky130_fd_sc_hd__a21bo_1 _20300_ (.A1(net9160),
    .A2(_12104_),
    .B1_N(_12105_),
    .X(_00484_));
 sky130_fd_sc_hd__nand2_1 _20301_ (.A(net6499),
    .B(net6471),
    .Y(_12106_));
 sky130_fd_sc_hd__nand2_1 _20302_ (.A(net6516),
    .B(net2600),
    .Y(_12107_));
 sky130_fd_sc_hd__a32o_1 _20303_ (.A1(net6516),
    .A2(net1481),
    .A3(_12106_),
    .B1(_12107_),
    .B2(_12092_),
    .X(_12108_));
 sky130_fd_sc_hd__nor2_1 _20304_ (.A(net4040),
    .B(net6478),
    .Y(_12109_));
 sky130_fd_sc_hd__mux2_1 _20305_ (.A0(net6467),
    .A1(_12109_),
    .S(net1808),
    .X(_12110_));
 sky130_fd_sc_hd__a221o_1 _20306_ (.A1(_09054_),
    .A2(_12098_),
    .B1(_12110_),
    .B2(net3313),
    .C1(net6459),
    .X(_12111_));
 sky130_fd_sc_hd__a21oi_1 _20307_ (.A1(net6479),
    .A2(_12108_),
    .B1(_12111_),
    .Y(_12112_));
 sky130_fd_sc_hd__o21bai_1 _20308_ (.A1(_12089_),
    .A2(_12100_),
    .B1_N(\cordic0.slte0.opA[1] ),
    .Y(_12113_));
 sky130_fd_sc_hd__nand2_1 _20309_ (.A(_12102_),
    .B(_12113_),
    .Y(_12114_));
 sky130_fd_sc_hd__xor2_1 _20310_ (.A(_12112_),
    .B(_12114_),
    .X(_12115_));
 sky130_fd_sc_hd__a21o_1 _20311_ (.A1(net1491),
    .A2(_12115_),
    .B1(net3317),
    .X(_12116_));
 sky130_fd_sc_hd__or3_1 _20312_ (.A(\cordic0.slte0.opA[2] ),
    .B(net2281),
    .C(_12115_),
    .X(_12117_));
 sky130_fd_sc_hd__a21bo_1 _20313_ (.A1(net9187),
    .A2(_12116_),
    .B1_N(_12117_),
    .X(_00485_));
 sky130_fd_sc_hd__nand2_1 _20314_ (.A(net4041),
    .B(net6477),
    .Y(_12118_));
 sky130_fd_sc_hd__a21o_1 _20315_ (.A1(net6467),
    .A2(_12118_),
    .B1(net6509),
    .X(_12119_));
 sky130_fd_sc_hd__nand2_1 _20316_ (.A(net1223),
    .B(_12119_),
    .Y(_12120_));
 sky130_fd_sc_hd__or3_1 _20317_ (.A(net6515),
    .B(net1482),
    .C(_08943_),
    .X(_12121_));
 sky130_fd_sc_hd__a221oi_1 _20318_ (.A1(net4037),
    .A2(_12098_),
    .B1(_12120_),
    .B2(_12121_),
    .C1(net6459),
    .Y(_12122_));
 sky130_fd_sc_hd__or2_1 _20319_ (.A(\cordic0.slte0.opA[2] ),
    .B(_12112_),
    .X(_12123_));
 sky130_fd_sc_hd__and2_1 _20320_ (.A(\cordic0.slte0.opA[2] ),
    .B(_12112_),
    .X(_12124_));
 sky130_fd_sc_hd__a31o_1 _20321_ (.A1(_12102_),
    .A2(_12113_),
    .A3(_12123_),
    .B1(_12124_),
    .X(_12125_));
 sky130_fd_sc_hd__or2_1 _20322_ (.A(net951),
    .B(_12125_),
    .X(_12126_));
 sky130_fd_sc_hd__nand2_1 _20323_ (.A(net951),
    .B(_12125_),
    .Y(_12127_));
 sky130_fd_sc_hd__nand2_1 _20324_ (.A(_12126_),
    .B(_12127_),
    .Y(_12128_));
 sky130_fd_sc_hd__a21o_1 _20325_ (.A1(net2182),
    .A2(_12128_),
    .B1(net4241),
    .X(_12129_));
 sky130_fd_sc_hd__nor2_1 _20326_ (.A(net1911),
    .B(_12128_),
    .Y(_12130_));
 sky130_fd_sc_hd__mux2_1 _20327_ (.A0(_12129_),
    .A1(_12130_),
    .S(_08885_),
    .X(_12131_));
 sky130_fd_sc_hd__clkbuf_1 _20328_ (.A(_12131_),
    .X(_00486_));
 sky130_fd_sc_hd__a2111o_1 _20329_ (.A1(net6479),
    .A2(net6472),
    .B1(net6466),
    .C1(_12084_),
    .D1(net3314),
    .X(_12132_));
 sky130_fd_sc_hd__nand2_2 _20330_ (.A(net2607),
    .B(_08990_),
    .Y(_12133_));
 sky130_fd_sc_hd__or2_1 _20331_ (.A(net3667),
    .B(_12133_),
    .X(_12134_));
 sky130_fd_sc_hd__clkbuf_1 _20332_ (.A(_12134_),
    .X(_12135_));
 sky130_fd_sc_hd__a21oi_1 _20333_ (.A1(net6515),
    .A2(net2586),
    .B1(net949),
    .Y(_12136_));
 sky130_fd_sc_hd__xnor2_1 _20334_ (.A(_12132_),
    .B(_12136_),
    .Y(_12137_));
 sky130_fd_sc_hd__a21o_1 _20335_ (.A1(net951),
    .A2(_12125_),
    .B1(\cordic0.slte0.opA[3] ),
    .X(_12138_));
 sky130_fd_sc_hd__and3_1 _20336_ (.A(_12126_),
    .B(_12137_),
    .C(_12138_),
    .X(_12139_));
 sky130_fd_sc_hd__a21o_1 _20337_ (.A1(_12126_),
    .A2(_12138_),
    .B1(_12137_),
    .X(_12140_));
 sky130_fd_sc_hd__and2b_1 _20338_ (.A_N(_12139_),
    .B(_12140_),
    .X(_12141_));
 sky130_fd_sc_hd__buf_1 _20339_ (.A(net1817),
    .X(_12142_));
 sky130_fd_sc_hd__nor2_1 _20340_ (.A(\cordic0.slte0.opA[4] ),
    .B(net1400),
    .Y(_12143_));
 sky130_fd_sc_hd__o21ai_1 _20341_ (.A1(net1400),
    .A2(_12141_),
    .B1(net8055),
    .Y(_12144_));
 sky130_fd_sc_hd__a22o_1 _20342_ (.A1(_12141_),
    .A2(_12143_),
    .B1(_12144_),
    .B2(net9218),
    .X(_00487_));
 sky130_fd_sc_hd__nor2_2 _20343_ (.A(net3668),
    .B(_12133_),
    .Y(_12145_));
 sky130_fd_sc_hd__nor2_1 _20344_ (.A(net2591),
    .B(_12090_),
    .Y(_12146_));
 sky130_fd_sc_hd__or4_1 _20345_ (.A(net6516),
    .B(net6466),
    .C(_08836_),
    .D(_12146_),
    .X(_12147_));
 sky130_fd_sc_hd__mux2_1 _20346_ (.A0(net1500),
    .A1(net1054),
    .S(_12147_),
    .X(_12148_));
 sky130_fd_sc_hd__a31o_1 _20347_ (.A1(_12126_),
    .A2(_12137_),
    .A3(_12138_),
    .B1(\cordic0.slte0.opA[4] ),
    .X(_12149_));
 sky130_fd_sc_hd__and3_1 _20348_ (.A(_12140_),
    .B(_12148_),
    .C(_12149_),
    .X(_12150_));
 sky130_fd_sc_hd__a21o_1 _20349_ (.A1(_12140_),
    .A2(_12149_),
    .B1(_12148_),
    .X(_12151_));
 sky130_fd_sc_hd__or2b_1 _20350_ (.A(_12150_),
    .B_N(_12151_),
    .X(_12152_));
 sky130_fd_sc_hd__a21o_1 _20351_ (.A1(net1490),
    .A2(_12152_),
    .B1(net3316),
    .X(_12153_));
 sky130_fd_sc_hd__or3_1 _20352_ (.A(\cordic0.slte0.opA[5] ),
    .B(net2280),
    .C(_12152_),
    .X(_12154_));
 sky130_fd_sc_hd__a21bo_1 _20353_ (.A1(net9168),
    .A2(_12153_),
    .B1_N(_12154_),
    .X(_00488_));
 sky130_fd_sc_hd__a31o_1 _20354_ (.A1(_12140_),
    .A2(_12148_),
    .A3(_12149_),
    .B1(\cordic0.slte0.opA[5] ),
    .X(_12155_));
 sky130_fd_sc_hd__nand2_1 _20355_ (.A(_12151_),
    .B(_12155_),
    .Y(_12156_));
 sky130_fd_sc_hd__a21o_1 _20356_ (.A1(net6472),
    .A2(net4037),
    .B1(_12084_),
    .X(_12157_));
 sky130_fd_sc_hd__a21oi_1 _20357_ (.A1(net6515),
    .A2(_12157_),
    .B1(_12096_),
    .Y(_12158_));
 sky130_fd_sc_hd__nor2_2 _20358_ (.A(net6458),
    .B(_12158_),
    .Y(_12159_));
 sky130_fd_sc_hd__xnor2_1 _20359_ (.A(net949),
    .B(_12159_),
    .Y(_12160_));
 sky130_fd_sc_hd__xnor2_1 _20360_ (.A(_12156_),
    .B(_12160_),
    .Y(_12161_));
 sky130_fd_sc_hd__o21ai_1 _20361_ (.A1(net1399),
    .A2(_12161_),
    .B1(net8041),
    .Y(_12162_));
 sky130_fd_sc_hd__nor2_1 _20362_ (.A(net6374),
    .B(net1558),
    .Y(_12163_));
 sky130_fd_sc_hd__a22o_1 _20363_ (.A1(net6374),
    .A2(_12162_),
    .B1(_12163_),
    .B2(_12161_),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _20364_ (.A0(net949),
    .A1(_12159_),
    .S(_12156_),
    .X(_12164_));
 sky130_fd_sc_hd__mux2_1 _20365_ (.A0(_12159_),
    .A1(net1054),
    .S(_12156_),
    .X(_12165_));
 sky130_fd_sc_hd__mux2_1 _20366_ (.A0(_12164_),
    .A1(_12165_),
    .S(net4055),
    .X(_12166_));
 sky130_fd_sc_hd__mux2_1 _20367_ (.A0(_08836_),
    .A1(_12157_),
    .S(net3314),
    .X(_12167_));
 sky130_fd_sc_hd__and2_1 _20368_ (.A(net2608),
    .B(_12167_),
    .X(_12168_));
 sky130_fd_sc_hd__xnor2_2 _20369_ (.A(\cordic0.slte0.opA[7] ),
    .B(_12168_),
    .Y(_12169_));
 sky130_fd_sc_hd__xnor2_1 _20370_ (.A(_12166_),
    .B(_12169_),
    .Y(_12170_));
 sky130_fd_sc_hd__a22o_1 _20371_ (.A1(net3355),
    .A2(\cordic0.slte0.opA[7] ),
    .B1(net1228),
    .B2(_12170_),
    .X(_00490_));
 sky130_fd_sc_hd__xnor2_1 _20372_ (.A(net6508),
    .B(_12109_),
    .Y(_12171_));
 sky130_fd_sc_hd__nor2_1 _20373_ (.A(_09006_),
    .B(_12171_),
    .Y(_12172_));
 sky130_fd_sc_hd__xnor2_1 _20374_ (.A(net950),
    .B(_12172_),
    .Y(_12173_));
 sky130_fd_sc_hd__nand2_1 _20375_ (.A(net6477),
    .B(net1223),
    .Y(_12174_));
 sky130_fd_sc_hd__nand2_1 _20376_ (.A(net3313),
    .B(net1501),
    .Y(_12175_));
 sky130_fd_sc_hd__o21a_1 _20377_ (.A1(_06504_),
    .A2(_12175_),
    .B1(_12098_),
    .X(_12176_));
 sky130_fd_sc_hd__mux2_1 _20378_ (.A0(_12174_),
    .A1(_12176_),
    .S(net6495),
    .X(_12177_));
 sky130_fd_sc_hd__o21ai_1 _20379_ (.A1(net4055),
    .A2(_12159_),
    .B1(_12168_),
    .Y(_12178_));
 sky130_fd_sc_hd__a211o_1 _20380_ (.A1(net6374),
    .A2(_12159_),
    .B1(_12168_),
    .C1(net1054),
    .X(_12179_));
 sky130_fd_sc_hd__o21ai_1 _20381_ (.A1(net949),
    .A2(_12178_),
    .B1(_12179_),
    .Y(_12180_));
 sky130_fd_sc_hd__inv_2 _20382_ (.A(\cordic0.slte0.opA[7] ),
    .Y(_12181_));
 sky130_fd_sc_hd__o32a_1 _20383_ (.A1(net6458),
    .A2(net4055),
    .A3(_12177_),
    .B1(_12180_),
    .B2(_12181_),
    .X(_12182_));
 sky130_fd_sc_hd__xnor2_1 _20384_ (.A(net6374),
    .B(_12159_),
    .Y(_12183_));
 sky130_fd_sc_hd__nor3_1 _20385_ (.A(net1054),
    .B(_12169_),
    .C(_12183_),
    .Y(_12184_));
 sky130_fd_sc_hd__and3_1 _20386_ (.A(net1054),
    .B(_12169_),
    .C(_12183_),
    .X(_12185_));
 sky130_fd_sc_hd__o211ai_1 _20387_ (.A1(_12184_),
    .A2(_12185_),
    .B1(_12151_),
    .C1(_12155_),
    .Y(_12186_));
 sky130_fd_sc_hd__and2_1 _20388_ (.A(_12182_),
    .B(net603),
    .X(_12187_));
 sky130_fd_sc_hd__xnor2_1 _20389_ (.A(net865),
    .B(_12187_),
    .Y(_12188_));
 sky130_fd_sc_hd__nor2_1 _20390_ (.A(\cordic0.slte0.opA[8] ),
    .B(net1399),
    .Y(_12189_));
 sky130_fd_sc_hd__o21ai_1 _20391_ (.A1(net1399),
    .A2(_12188_),
    .B1(net8053),
    .Y(_12190_));
 sky130_fd_sc_hd__a22o_1 _20392_ (.A1(_12188_),
    .A2(_12189_),
    .B1(_12190_),
    .B2(net9188),
    .X(_00491_));
 sky130_fd_sc_hd__inv_2 _20393_ (.A(\cordic0.slte0.opA[9] ),
    .Y(_12191_));
 sky130_fd_sc_hd__nand2_1 _20394_ (.A(_08836_),
    .B(net1501),
    .Y(_12192_));
 sky130_fd_sc_hd__nand2_1 _20395_ (.A(_08835_),
    .B(net1223),
    .Y(_12193_));
 sky130_fd_sc_hd__a21o_1 _20396_ (.A1(_12192_),
    .A2(_12193_),
    .B1(net3313),
    .X(_12194_));
 sky130_fd_sc_hd__o311a_1 _20397_ (.A1(net6467),
    .A2(net4037),
    .A3(_12175_),
    .B1(_12194_),
    .C1(_12098_),
    .X(_12195_));
 sky130_fd_sc_hd__nor2_1 _20398_ (.A(net6458),
    .B(_12195_),
    .Y(_12196_));
 sky130_fd_sc_hd__nand2_1 _20399_ (.A(\cordic0.slte0.opA[8] ),
    .B(net865),
    .Y(_12197_));
 sky130_fd_sc_hd__or2_1 _20400_ (.A(\cordic0.slte0.opA[8] ),
    .B(net865),
    .X(_12198_));
 sky130_fd_sc_hd__a21bo_1 _20401_ (.A1(_12187_),
    .A2(_12197_),
    .B1_N(_12198_),
    .X(_12199_));
 sky130_fd_sc_hd__xor2_1 _20402_ (.A(net811),
    .B(_12199_),
    .X(_12200_));
 sky130_fd_sc_hd__a21oi_1 _20403_ (.A1(net1466),
    .A2(_12200_),
    .B1(net3355),
    .Y(_12201_));
 sky130_fd_sc_hd__or3_1 _20404_ (.A(\cordic0.slte0.opA[9] ),
    .B(net1915),
    .C(_12200_),
    .X(_12202_));
 sky130_fd_sc_hd__o21ai_1 _20405_ (.A1(_12191_),
    .A2(_12201_),
    .B1(_12202_),
    .Y(_00492_));
 sky130_fd_sc_hd__a21o_1 _20406_ (.A1(net6485),
    .A2(net4050),
    .B1(_12109_),
    .X(_12203_));
 sky130_fd_sc_hd__nand2_1 _20407_ (.A(_09082_),
    .B(_12203_),
    .Y(_12204_));
 sky130_fd_sc_hd__xnor2_2 _20408_ (.A(_12145_),
    .B(net2089),
    .Y(_12205_));
 sky130_fd_sc_hd__and2b_1 _20409_ (.A_N(net811),
    .B(_12197_),
    .X(_12206_));
 sky130_fd_sc_hd__and2_1 _20410_ (.A(_12191_),
    .B(_12197_),
    .X(_12207_));
 sky130_fd_sc_hd__o211ai_1 _20411_ (.A1(_12206_),
    .A2(_12207_),
    .B1(_12182_),
    .C1(net603),
    .Y(_12208_));
 sky130_fd_sc_hd__a21o_1 _20412_ (.A1(\cordic0.slte0.opA[9] ),
    .A2(_12198_),
    .B1(net811),
    .X(_12209_));
 sky130_fd_sc_hd__o211a_1 _20413_ (.A1(\cordic0.slte0.opA[9] ),
    .A2(_12198_),
    .B1(_12208_),
    .C1(_12209_),
    .X(_12210_));
 sky130_fd_sc_hd__xnor2_1 _20414_ (.A(_12205_),
    .B(_12210_),
    .Y(_12211_));
 sky130_fd_sc_hd__a21o_1 _20415_ (.A1(_06506_),
    .A2(_12211_),
    .B1(net4239),
    .X(_12212_));
 sky130_fd_sc_hd__nor2_1 _20416_ (.A(net1915),
    .B(_12211_),
    .Y(_12213_));
 sky130_fd_sc_hd__mux2_1 _20417_ (.A0(_12212_),
    .A1(_12213_),
    .S(_08865_),
    .X(_12214_));
 sky130_fd_sc_hd__clkbuf_1 _20418_ (.A(_12214_),
    .X(_00493_));
 sky130_fd_sc_hd__or2_1 _20419_ (.A(_12090_),
    .B(net1500),
    .X(_12215_));
 sky130_fd_sc_hd__or3_1 _20420_ (.A(net6467),
    .B(_12118_),
    .C(_12175_),
    .X(_12216_));
 sky130_fd_sc_hd__a21o_1 _20421_ (.A1(_12174_),
    .A2(_12192_),
    .B1(net3313),
    .X(_12217_));
 sky130_fd_sc_hd__a31oi_1 _20422_ (.A1(_12215_),
    .A2(_12216_),
    .A3(_12217_),
    .B1(net6459),
    .Y(_12218_));
 sky130_fd_sc_hd__o21a_1 _20423_ (.A1(_12205_),
    .A2(_12210_),
    .B1(\cordic0.slte0.opA[10] ),
    .X(_12219_));
 sky130_fd_sc_hd__a21oi_1 _20424_ (.A1(_12205_),
    .A2(_12210_),
    .B1(_12219_),
    .Y(_12220_));
 sky130_fd_sc_hd__xnor2_1 _20425_ (.A(net863),
    .B(_12220_),
    .Y(_12221_));
 sky130_fd_sc_hd__o21ai_1 _20426_ (.A1(net1832),
    .A2(_12221_),
    .B1(net8045),
    .Y(_12222_));
 sky130_fd_sc_hd__nor2_1 _20427_ (.A(\cordic0.slte0.opA[11] ),
    .B(net1559),
    .Y(_12223_));
 sky130_fd_sc_hd__a22o_1 _20428_ (.A1(\cordic0.slte0.opA[11] ),
    .A2(_12222_),
    .B1(_12223_),
    .B2(_12221_),
    .X(_00494_));
 sky130_fd_sc_hd__inv_2 _20429_ (.A(_12133_),
    .Y(_12224_));
 sky130_fd_sc_hd__and2_1 _20430_ (.A(net2596),
    .B(net2166),
    .X(_12225_));
 sky130_fd_sc_hd__mux2_2 _20431_ (.A0(net950),
    .A1(_12224_),
    .S(_12225_),
    .X(_12226_));
 sky130_fd_sc_hd__a221o_1 _20432_ (.A1(_12205_),
    .A2(_12210_),
    .B1(net863),
    .B2(\cordic0.slte0.opA[11] ),
    .C1(_12219_),
    .X(_12227_));
 sky130_fd_sc_hd__o21a_1 _20433_ (.A1(\cordic0.slte0.opA[11] ),
    .A2(net863),
    .B1(_12227_),
    .X(_12228_));
 sky130_fd_sc_hd__xor2_1 _20434_ (.A(_12226_),
    .B(_12228_),
    .X(_12229_));
 sky130_fd_sc_hd__a21o_1 _20435_ (.A1(net1487),
    .A2(_12229_),
    .B1(net3315),
    .X(_12230_));
 sky130_fd_sc_hd__or3_1 _20436_ (.A(\cordic0.slte0.opA[12] ),
    .B(net2279),
    .C(_12229_),
    .X(_12231_));
 sky130_fd_sc_hd__a21bo_1 _20437_ (.A1(net6370),
    .A2(_12230_),
    .B1_N(_12231_),
    .X(_00495_));
 sky130_fd_sc_hd__nand2_1 _20438_ (.A(net6493),
    .B(net2166),
    .Y(_12232_));
 sky130_fd_sc_hd__nor2_1 _20439_ (.A(net6511),
    .B(_12232_),
    .Y(_12233_));
 sky130_fd_sc_hd__xnor2_1 _20440_ (.A(net6369),
    .B(_12233_),
    .Y(_12234_));
 sky130_fd_sc_hd__xnor2_1 _20441_ (.A(net950),
    .B(_12234_),
    .Y(_12235_));
 sky130_fd_sc_hd__inv_2 _20442_ (.A(_12228_),
    .Y(_12236_));
 sky130_fd_sc_hd__o21a_1 _20443_ (.A1(_12226_),
    .A2(_12236_),
    .B1(_08857_),
    .X(_12237_));
 sky130_fd_sc_hd__a21oi_1 _20444_ (.A1(_12226_),
    .A2(_12236_),
    .B1(_12237_),
    .Y(_12238_));
 sky130_fd_sc_hd__xnor2_1 _20445_ (.A(_12235_),
    .B(_12238_),
    .Y(_12239_));
 sky130_fd_sc_hd__a22o_1 _20446_ (.A1(net3354),
    .A2(net6369),
    .B1(net1229),
    .B2(_12239_),
    .X(_00496_));
 sky130_fd_sc_hd__xnor2_1 _20447_ (.A(_08857_),
    .B(_12226_),
    .Y(_12240_));
 sky130_fd_sc_hd__a22o_1 _20448_ (.A1(net6511),
    .A2(_12133_),
    .B1(_12145_),
    .B2(_12233_),
    .X(_12241_));
 sky130_fd_sc_hd__a21oi_1 _20449_ (.A1(net6370),
    .A2(_12232_),
    .B1(net6369),
    .Y(_12242_));
 sky130_fd_sc_hd__a221o_1 _20450_ (.A1(net950),
    .A2(_12232_),
    .B1(_12241_),
    .B2(_08857_),
    .C1(_12242_),
    .X(_12243_));
 sky130_fd_sc_hd__o31a_1 _20451_ (.A1(_12236_),
    .A2(_12235_),
    .A3(_12240_),
    .B1(_12243_),
    .X(_12244_));
 sky130_fd_sc_hd__a31oi_1 _20452_ (.A1(net6515),
    .A2(net1501),
    .A3(net2586),
    .B1(_12136_),
    .Y(_12245_));
 sky130_fd_sc_hd__xor2_1 _20453_ (.A(_12244_),
    .B(net809),
    .X(_12246_));
 sky130_fd_sc_hd__o21ai_1 _20454_ (.A1(net1830),
    .A2(_12246_),
    .B1(net8044),
    .Y(_12247_));
 sky130_fd_sc_hd__nor2_1 _20455_ (.A(\cordic0.slte0.opA[14] ),
    .B(_06509_),
    .Y(_12248_));
 sky130_fd_sc_hd__a22o_1 _20456_ (.A1(net9191),
    .A2(_12247_),
    .B1(_12248_),
    .B2(_12246_),
    .X(_00497_));
 sky130_fd_sc_hd__o21a_1 _20457_ (.A1(net3667),
    .A2(net967),
    .B1(net2607),
    .X(_12249_));
 sky130_fd_sc_hd__nand2_1 _20458_ (.A(net8044),
    .B(\cordic0.slte0.opA[15] ),
    .Y(_12250_));
 sky130_fd_sc_hd__a21bo_1 _20459_ (.A1(_12244_),
    .A2(net809),
    .B1_N(\cordic0.slte0.opA[14] ),
    .X(_12251_));
 sky130_fd_sc_hd__o21a_1 _20460_ (.A1(_12244_),
    .A2(net809),
    .B1(_12251_),
    .X(_12252_));
 sky130_fd_sc_hd__mux2_1 _20461_ (.A0(_12250_),
    .A1(\cordic0.slte0.opA[15] ),
    .S(_12252_),
    .X(_12253_));
 sky130_fd_sc_hd__mux2_1 _20462_ (.A0(\cordic0.slte0.opA[15] ),
    .A1(_12250_),
    .S(_12252_),
    .X(_12254_));
 sky130_fd_sc_hd__o21bai_1 _20463_ (.A1(net3667),
    .A2(_12224_),
    .B1_N(_12254_),
    .Y(_12255_));
 sky130_fd_sc_hd__o221a_1 _20464_ (.A1(net8044),
    .A2(\cordic0.slte0.opA[15] ),
    .B1(_12249_),
    .B2(_12253_),
    .C1(_12255_),
    .X(_00498_));
 sky130_fd_sc_hd__nand2_1 _20465_ (.A(\cordic0.slte0.opA[15] ),
    .B(_12249_),
    .Y(_12256_));
 sky130_fd_sc_hd__nor2_1 _20466_ (.A(\cordic0.slte0.opA[15] ),
    .B(_12249_),
    .Y(_12257_));
 sky130_fd_sc_hd__a21o_1 _20467_ (.A1(_12252_),
    .A2(_12256_),
    .B1(_12257_),
    .X(_12258_));
 sky130_fd_sc_hd__xnor2_1 _20468_ (.A(_12133_),
    .B(_12258_),
    .Y(_12259_));
 sky130_fd_sc_hd__and3_1 _20469_ (.A(\cordic0.slte0.opA[16] ),
    .B(net1810),
    .C(_12259_),
    .X(_12260_));
 sky130_fd_sc_hd__and3b_1 _20470_ (.A_N(_12259_),
    .B(_08900_),
    .C(net1810),
    .X(_12261_));
 sky130_fd_sc_hd__a211o_1 _20471_ (.A1(net3353),
    .A2(net9153),
    .B1(_12260_),
    .C1(_12261_),
    .X(_00499_));
 sky130_fd_sc_hd__a32o_1 _20472_ (.A1(net8044),
    .A2(_12224_),
    .A3(_12258_),
    .B1(\cordic0.slte0.opA[17] ),
    .B2(net2178),
    .X(_12262_));
 sky130_fd_sc_hd__a21o_1 _20473_ (.A1(net2178),
    .A2(_12258_),
    .B1(net3353),
    .X(_12263_));
 sky130_fd_sc_hd__a22o_1 _20474_ (.A1(net4054),
    .A2(_12262_),
    .B1(_12263_),
    .B2(net9216),
    .X(_00500_));
 sky130_fd_sc_hd__mux4_1 _20475_ (.A0(net6890),
    .A1(net6853),
    .A2(net6840),
    .A3(net6824),
    .S0(net6521),
    .S1(net6488),
    .X(_12264_));
 sky130_fd_sc_hd__mux4_1 _20476_ (.A0(net7056),
    .A1(net7010),
    .A2(net7042),
    .A3(net6983),
    .S0(net6489),
    .S1(net6512),
    .X(_12265_));
 sky130_fd_sc_hd__mux4_1 _20477_ (.A0(net6962),
    .A1(net6917),
    .A2(net6937),
    .A3(net6904),
    .S0(net6491),
    .S1(net6521),
    .X(_12266_));
 sky130_fd_sc_hd__mux4_1 _20478_ (.A0(net7147),
    .A1(net7129),
    .A2(net7113),
    .A3(net7088),
    .S0(net6512),
    .S1(net6489),
    .X(_12267_));
 sky130_fd_sc_hd__mux4_1 _20479_ (.A0(net3854),
    .A1(net3853),
    .A2(net3852),
    .A3(net3851),
    .S0(net3335),
    .S1(net4060),
    .X(_12268_));
 sky130_fd_sc_hd__mux2_1 _20480_ (.A0(net6804),
    .A1(net6763),
    .S(net6523),
    .X(_12269_));
 sky130_fd_sc_hd__mux2_1 _20481_ (.A0(net6758),
    .A1(net3849),
    .S(_08836_),
    .X(_12270_));
 sky130_fd_sc_hd__mux2_1 _20482_ (.A0(_12268_),
    .A1(_12270_),
    .S(net6461),
    .X(_12271_));
 sky130_fd_sc_hd__or2_1 _20483_ (.A(net2192),
    .B(net2087),
    .X(_12272_));
 sky130_fd_sc_hd__a21oi_1 _20484_ (.A1(net1237),
    .A2(net2087),
    .B1(net3170),
    .Y(_12273_));
 sky130_fd_sc_hd__a31o_1 _20485_ (.A1(net8057),
    .A2(net3170),
    .A3(_12272_),
    .B1(_12273_),
    .X(_00501_));
 sky130_fd_sc_hd__mux4_1 _20486_ (.A0(net6853),
    .A1(net6824),
    .A2(net6840),
    .A3(net6790),
    .S0(net6491),
    .S1(net6521),
    .X(_12274_));
 sky130_fd_sc_hd__mux4_1 _20487_ (.A0(net7042),
    .A1(net7010),
    .A2(net6983),
    .A3(net6971),
    .S0(net6514),
    .S1(net6489),
    .X(_12275_));
 sky130_fd_sc_hd__mux4_1 _20488_ (.A0(net6935),
    .A1(net6917),
    .A2(net6904),
    .A3(net6890),
    .S0(net6513),
    .S1(net6491),
    .X(_12276_));
 sky130_fd_sc_hd__mux4_1 _20489_ (.A0(net7129),
    .A1(net7113),
    .A2(net7088),
    .A3(net7056),
    .S0(net6507),
    .S1(net6489),
    .X(_12277_));
 sky130_fd_sc_hd__mux4_1 _20490_ (.A0(net3848),
    .A1(_12275_),
    .A2(net3847),
    .A3(_12277_),
    .S0(net3334),
    .S1(net3333),
    .X(_12278_));
 sky130_fd_sc_hd__mux2_1 _20491_ (.A0(net6758),
    .A1(net2492),
    .S(net3345),
    .X(_12279_));
 sky130_fd_sc_hd__nand2_1 _20492_ (.A(net6363),
    .B(net970),
    .Y(_12280_));
 sky130_fd_sc_hd__nand2_1 _20493_ (.A(net3169),
    .B(net1499),
    .Y(_12281_));
 sky130_fd_sc_hd__inv_2 _20494_ (.A(net2088),
    .Y(_12282_));
 sky130_fd_sc_hd__a21oi_1 _20495_ (.A1(_12280_),
    .A2(_12281_),
    .B1(_12282_),
    .Y(_12283_));
 sky130_fd_sc_hd__xnor2_1 _20496_ (.A(net2086),
    .B(_12283_),
    .Y(_12284_));
 sky130_fd_sc_hd__nand2_1 _20497_ (.A(net6350),
    .B(net1471),
    .Y(_12285_));
 sky130_fd_sc_hd__a21oi_1 _20498_ (.A1(net2183),
    .A2(_12284_),
    .B1(net3359),
    .Y(_12286_));
 sky130_fd_sc_hd__o22a_1 _20499_ (.A1(_12284_),
    .A2(_12285_),
    .B1(_12286_),
    .B2(net6350),
    .X(_00502_));
 sky130_fd_sc_hd__inv_2 _20500_ (.A(net2086),
    .Y(_12287_));
 sky130_fd_sc_hd__a21oi_1 _20501_ (.A1(net1484),
    .A2(_12287_),
    .B1(net3169),
    .Y(_12288_));
 sky130_fd_sc_hd__or4_1 _20502_ (.A(net6363),
    .B(net1823),
    .C(_12282_),
    .D(net2086),
    .X(_12289_));
 sky130_fd_sc_hd__a21boi_1 _20503_ (.A1(net3169),
    .A2(net2088),
    .B1_N(net6350),
    .Y(_12290_));
 sky130_fd_sc_hd__a211o_1 _20504_ (.A1(net1484),
    .A2(net2088),
    .B1(_12287_),
    .C1(_12290_),
    .X(_12291_));
 sky130_fd_sc_hd__o311a_1 _20505_ (.A1(net6350),
    .A2(_12282_),
    .A3(_12288_),
    .B1(_12289_),
    .C1(_12291_),
    .X(_12292_));
 sky130_fd_sc_hd__a211o_1 _20506_ (.A1(_08836_),
    .A2(net3849),
    .B1(net3345),
    .C1(net6766),
    .X(_12293_));
 sky130_fd_sc_hd__o31a_1 _20507_ (.A1(net6461),
    .A2(_12268_),
    .A3(net2492),
    .B1(_12293_),
    .X(_12294_));
 sky130_fd_sc_hd__mux4_2 _20508_ (.A0(net6841),
    .A1(net6824),
    .A2(net6790),
    .A3(net6762),
    .S0(net6521),
    .S1(net6491),
    .X(_12295_));
 sky130_fd_sc_hd__mux4_1 _20509_ (.A0(net6917),
    .A1(net6890),
    .A2(net6904),
    .A3(net6871),
    .S0(net6491),
    .S1(net6521),
    .X(_12296_));
 sky130_fd_sc_hd__mux4_1 _20510_ (.A0(net7010),
    .A1(net6983),
    .A2(net6962),
    .A3(net6938),
    .S0(net6514),
    .S1(net6490),
    .X(_12297_));
 sky130_fd_sc_hd__mux4_1 _20511_ (.A0(net7113),
    .A1(net7088),
    .A2(net7056),
    .A3(net7042),
    .S0(net6514),
    .S1(net6489),
    .X(_12298_));
 sky130_fd_sc_hd__mux4_1 _20512_ (.A0(_12295_),
    .A1(net3846),
    .A2(_12297_),
    .A3(net3845),
    .S0(net4060),
    .S1(net3334),
    .X(_12299_));
 sky130_fd_sc_hd__mux2_1 _20513_ (.A0(net6766),
    .A1(net2491),
    .S(net3345),
    .X(_12300_));
 sky130_fd_sc_hd__a21o_1 _20514_ (.A1(net1484),
    .A2(net2084),
    .B1(net2082),
    .X(_12301_));
 sky130_fd_sc_hd__nand3_1 _20515_ (.A(net1484),
    .B(net2082),
    .C(net2084),
    .Y(_12302_));
 sky130_fd_sc_hd__nand2_1 _20516_ (.A(_12301_),
    .B(_12302_),
    .Y(_12303_));
 sky130_fd_sc_hd__or2_1 _20517_ (.A(net1053),
    .B(_12303_),
    .X(_12304_));
 sky130_fd_sc_hd__nand2_1 _20518_ (.A(net1053),
    .B(_12303_),
    .Y(_12305_));
 sky130_fd_sc_hd__nand2_1 _20519_ (.A(_12304_),
    .B(_12305_),
    .Y(_12306_));
 sky130_fd_sc_hd__nand2_1 _20520_ (.A(net6324),
    .B(net1470),
    .Y(_12307_));
 sky130_fd_sc_hd__a21oi_1 _20521_ (.A1(net1470),
    .A2(_12306_),
    .B1(_08909_),
    .Y(_12308_));
 sky130_fd_sc_hd__o22a_1 _20522_ (.A1(_12306_),
    .A2(_12307_),
    .B1(_12308_),
    .B2(net6324),
    .X(_00503_));
 sky130_fd_sc_hd__nand2_1 _20523_ (.A(net6324),
    .B(_12304_),
    .Y(_12309_));
 sky130_fd_sc_hd__or2_1 _20524_ (.A(net2082),
    .B(net2084),
    .X(_12310_));
 sky130_fd_sc_hd__nand2_1 _20525_ (.A(net1479),
    .B(_12310_),
    .Y(_12311_));
 sky130_fd_sc_hd__mux2_1 _20526_ (.A0(net6823),
    .A1(net6767),
    .S(net6502),
    .X(_12312_));
 sky130_fd_sc_hd__a22o_1 _20527_ (.A1(net6804),
    .A2(_08945_),
    .B1(_12312_),
    .B2(_08824_),
    .X(_12313_));
 sky130_fd_sc_hd__mux4_1 _20528_ (.A0(net6983),
    .A1(net6938),
    .A2(net6962),
    .A3(net6923),
    .S0(net6490),
    .S1(net6513),
    .X(_12314_));
 sky130_fd_sc_hd__mux4_2 _20529_ (.A0(net6901),
    .A1(net6853),
    .A2(net6890),
    .A3(net6840),
    .S0(net6490),
    .S1(net6513),
    .X(_12315_));
 sky130_fd_sc_hd__mux4_1 _20530_ (.A0(net7088),
    .A1(net7042),
    .A2(net7074),
    .A3(net7010),
    .S0(net6489),
    .S1(net6514),
    .X(_12316_));
 sky130_fd_sc_hd__mux4_1 _20531_ (.A0(net3124),
    .A1(_12314_),
    .A2(_12315_),
    .A3(_12316_),
    .S0(net3334),
    .S1(net3332),
    .X(_12317_));
 sky130_fd_sc_hd__a22oi_1 _20532_ (.A1(net6756),
    .A2(_08944_),
    .B1(net2490),
    .B2(_08924_),
    .Y(_12318_));
 sky130_fd_sc_hd__xnor2_1 _20533_ (.A(net3193),
    .B(net2079),
    .Y(_12319_));
 sky130_fd_sc_hd__xnor2_1 _20534_ (.A(_12311_),
    .B(_12319_),
    .Y(_12320_));
 sky130_fd_sc_hd__a21oi_1 _20535_ (.A1(_12305_),
    .A2(_12309_),
    .B1(_12320_),
    .Y(_12321_));
 sky130_fd_sc_hd__and3_1 _20536_ (.A(_12305_),
    .B(_12320_),
    .C(_12309_),
    .X(_12322_));
 sky130_fd_sc_hd__o32a_1 _20537_ (.A1(net1398),
    .A2(_12321_),
    .A3(_12322_),
    .B1(net6306),
    .B2(net8056),
    .X(_00504_));
 sky130_fd_sc_hd__a21o_1 _20538_ (.A1(net1479),
    .A2(_12310_),
    .B1(net6326),
    .X(_12323_));
 sky130_fd_sc_hd__mux2_1 _20539_ (.A0(net6310),
    .A1(net1484),
    .S(net2082),
    .X(_12324_));
 sky130_fd_sc_hd__a21o_1 _20540_ (.A1(_12323_),
    .A2(_12324_),
    .B1(net2079),
    .X(_12325_));
 sky130_fd_sc_hd__a31o_1 _20541_ (.A1(net1484),
    .A2(net2082),
    .A3(net2079),
    .B1(net3193),
    .X(_12326_));
 sky130_fd_sc_hd__or2b_1 _20542_ (.A(net6326),
    .B_N(_12326_),
    .X(_12327_));
 sky130_fd_sc_hd__or4bb_1 _20543_ (.A(net1822),
    .B(net2082),
    .C_N(net2084),
    .D_N(net2079),
    .X(_12328_));
 sky130_fd_sc_hd__inv_2 _20544_ (.A(net2079),
    .Y(_12329_));
 sky130_fd_sc_hd__a21o_1 _20545_ (.A1(net2084),
    .A2(_12329_),
    .B1(net6310),
    .X(_12330_));
 sky130_fd_sc_hd__or3_1 _20546_ (.A(net1822),
    .B(net2084),
    .C(_12329_),
    .X(_12331_));
 sky130_fd_sc_hd__a21bo_1 _20547_ (.A1(_12330_),
    .A2(_12331_),
    .B1_N(net2082),
    .X(_12332_));
 sky130_fd_sc_hd__nand4_2 _20548_ (.A(_12325_),
    .B(_12327_),
    .C(_12328_),
    .D(_12332_),
    .Y(_12333_));
 sky130_fd_sc_hd__a21oi_1 _20549_ (.A1(_12301_),
    .A2(_12302_),
    .B1(net6326),
    .Y(_12334_));
 sky130_fd_sc_hd__and3_1 _20550_ (.A(net6326),
    .B(_12301_),
    .C(_12302_),
    .X(_12335_));
 sky130_fd_sc_hd__o211ai_2 _20551_ (.A1(_12334_),
    .A2(_12335_),
    .B1(net1053),
    .C1(_12320_),
    .Y(_12336_));
 sky130_fd_sc_hd__nand2_1 _20552_ (.A(_12333_),
    .B(_12336_),
    .Y(_12337_));
 sky130_fd_sc_hd__mux2_1 _20553_ (.A0(net3854),
    .A1(net3853),
    .S(net3335),
    .X(_12338_));
 sky130_fd_sc_hd__or2_1 _20554_ (.A(net6480),
    .B(_12338_),
    .X(_12339_));
 sky130_fd_sc_hd__a221o_1 _20555_ (.A1(net2600),
    .A2(net3852),
    .B1(net3849),
    .B2(_08970_),
    .C1(_08971_),
    .X(_12340_));
 sky130_fd_sc_hd__a32o_1 _20556_ (.A1(net3345),
    .A2(_12339_),
    .A3(_12340_),
    .B1(net6766),
    .B2(_08973_),
    .X(_12341_));
 sky130_fd_sc_hd__or3_1 _20557_ (.A(net2082),
    .B(net2084),
    .C(_12329_),
    .X(_12342_));
 sky130_fd_sc_hd__nand2_1 _20558_ (.A(net1480),
    .B(_12342_),
    .Y(_12343_));
 sky130_fd_sc_hd__xnor2_2 _20559_ (.A(net1745),
    .B(_12343_),
    .Y(_12344_));
 sky130_fd_sc_hd__xnor2_1 _20560_ (.A(_12337_),
    .B(_12344_),
    .Y(_12345_));
 sky130_fd_sc_hd__or2_1 _20561_ (.A(net2192),
    .B(_12345_),
    .X(_12346_));
 sky130_fd_sc_hd__a21oi_1 _20562_ (.A1(net1237),
    .A2(_12345_),
    .B1(net2516),
    .Y(_12347_));
 sky130_fd_sc_hd__a31o_1 _20563_ (.A1(net8057),
    .A2(net2516),
    .A3(_12346_),
    .B1(_12347_),
    .X(_00505_));
 sky130_fd_sc_hd__a21o_1 _20564_ (.A1(_12333_),
    .A2(_12336_),
    .B1(_12344_),
    .X(_12348_));
 sky130_fd_sc_hd__a31o_1 _20565_ (.A1(_12333_),
    .A2(_12336_),
    .A3(_12344_),
    .B1(net2516),
    .X(_12349_));
 sky130_fd_sc_hd__mux2_1 _20566_ (.A0(net3848),
    .A1(_12275_),
    .S(net2602),
    .X(_12350_));
 sky130_fd_sc_hd__nand2_1 _20567_ (.A(net6470),
    .B(net3927),
    .Y(_12351_));
 sky130_fd_sc_hd__o21a_1 _20568_ (.A1(net3325),
    .A2(net3847),
    .B1(_12351_),
    .X(_12352_));
 sky130_fd_sc_hd__nand2_1 _20569_ (.A(net6464),
    .B(net3927),
    .Y(_12353_));
 sky130_fd_sc_hd__o221a_1 _20570_ (.A1(_09008_),
    .A2(_12350_),
    .B1(_12352_),
    .B2(net3333),
    .C1(_12353_),
    .X(_12354_));
 sky130_fd_sc_hd__o21a_1 _20571_ (.A1(net1745),
    .A2(_12342_),
    .B1(net1480),
    .X(_12355_));
 sky130_fd_sc_hd__xnor2_1 _20572_ (.A(net1742),
    .B(_12355_),
    .Y(_12356_));
 sky130_fd_sc_hd__a21boi_1 _20573_ (.A1(_12348_),
    .A2(_12349_),
    .B1_N(_12356_),
    .Y(_12357_));
 sky130_fd_sc_hd__nand3b_1 _20574_ (.A_N(_12356_),
    .B(_12348_),
    .C(_12349_),
    .Y(_12358_));
 sky130_fd_sc_hd__and2b_1 _20575_ (.A_N(_12357_),
    .B(_12358_),
    .X(_12359_));
 sky130_fd_sc_hd__o21ai_1 _20576_ (.A1(net1398),
    .A2(_12359_),
    .B1(net8056),
    .Y(_12360_));
 sky130_fd_sc_hd__and3_1 _20577_ (.A(net6253),
    .B(net1492),
    .C(_12359_),
    .X(_12361_));
 sky130_fd_sc_hd__a21oi_1 _20578_ (.A1(net3174),
    .A2(_12360_),
    .B1(_12361_),
    .Y(_00506_));
 sky130_fd_sc_hd__o21ai_1 _20579_ (.A1(net6255),
    .A2(_12357_),
    .B1(_12358_),
    .Y(_12362_));
 sky130_fd_sc_hd__o21a_1 _20580_ (.A1(net3325),
    .A2(net3846),
    .B1(_12351_),
    .X(_12363_));
 sky130_fd_sc_hd__mux2_1 _20581_ (.A0(_12295_),
    .A1(_12297_),
    .S(net2602),
    .X(_12364_));
 sky130_fd_sc_hd__o221a_1 _20582_ (.A1(net2594),
    .A2(_12363_),
    .B1(_12364_),
    .B2(_09008_),
    .C1(_12353_),
    .X(_12365_));
 sky130_fd_sc_hd__inv_2 _20583_ (.A(net1740),
    .Y(_12366_));
 sky130_fd_sc_hd__or3_2 _20584_ (.A(net1745),
    .B(_12342_),
    .C(net1742),
    .X(_12367_));
 sky130_fd_sc_hd__nand2_1 _20585_ (.A(_08991_),
    .B(_12367_),
    .Y(_12368_));
 sky130_fd_sc_hd__xnor2_2 _20586_ (.A(_12366_),
    .B(_12368_),
    .Y(_12369_));
 sky130_fd_sc_hd__and2b_1 _20587_ (.A_N(_12362_),
    .B(_12369_),
    .X(_12370_));
 sky130_fd_sc_hd__or2b_1 _20588_ (.A(_12369_),
    .B_N(_12362_),
    .X(_12371_));
 sky130_fd_sc_hd__and2b_1 _20589_ (.A_N(_12370_),
    .B(_12371_),
    .X(_12372_));
 sky130_fd_sc_hd__or2_1 _20590_ (.A(net2192),
    .B(_12372_),
    .X(_12373_));
 sky130_fd_sc_hd__a21oi_1 _20591_ (.A1(net1237),
    .A2(_12372_),
    .B1(net3164),
    .Y(_12374_));
 sky130_fd_sc_hd__a31o_1 _20592_ (.A1(net8057),
    .A2(net3164),
    .A3(_12373_),
    .B1(_12374_),
    .X(_00507_));
 sky130_fd_sc_hd__o21ai_1 _20593_ (.A1(net1740),
    .A2(_12367_),
    .B1(net1226),
    .Y(_12375_));
 sky130_fd_sc_hd__mux2_1 _20594_ (.A0(net3124),
    .A1(_12314_),
    .S(_09004_),
    .X(_12376_));
 sky130_fd_sc_hd__a22o_1 _20595_ (.A1(_09069_),
    .A2(_12376_),
    .B1(_12315_),
    .B2(_09029_),
    .X(_12377_));
 sky130_fd_sc_hd__a22oi_1 _20596_ (.A1(net6756),
    .A2(_09035_),
    .B1(_12377_),
    .B2(net2609),
    .Y(_12378_));
 sky130_fd_sc_hd__xnor2_1 _20597_ (.A(net6196),
    .B(net1396),
    .Y(_12379_));
 sky130_fd_sc_hd__xnor2_1 _20598_ (.A(_12375_),
    .B(_12379_),
    .Y(_12380_));
 sky130_fd_sc_hd__a21o_1 _20599_ (.A1(net6239),
    .A2(_12371_),
    .B1(_12370_),
    .X(_12381_));
 sky130_fd_sc_hd__xnor2_1 _20600_ (.A(_12380_),
    .B(_12381_),
    .Y(_12382_));
 sky130_fd_sc_hd__o22a_1 _20601_ (.A1(net8057),
    .A2(net6212),
    .B1(net1554),
    .B2(_12382_),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _20602_ (.A0(net3914),
    .A1(net1822),
    .S(net1740),
    .X(_12383_));
 sky130_fd_sc_hd__a21oi_1 _20603_ (.A1(net3163),
    .A2(_12375_),
    .B1(_12383_),
    .Y(_12384_));
 sky130_fd_sc_hd__inv_2 _20604_ (.A(_12367_),
    .Y(_12385_));
 sky130_fd_sc_hd__nor2_1 _20605_ (.A(_12385_),
    .B(net1396),
    .Y(_12386_));
 sky130_fd_sc_hd__nand2_1 _20606_ (.A(net1480),
    .B(net1396),
    .Y(_12387_));
 sky130_fd_sc_hd__o22a_1 _20607_ (.A1(net6195),
    .A2(_12386_),
    .B1(_12387_),
    .B2(_12367_),
    .X(_12388_));
 sky130_fd_sc_hd__o21a_1 _20608_ (.A1(_12366_),
    .A2(_12387_),
    .B1(net6195),
    .X(_12389_));
 sky130_fd_sc_hd__o32a_1 _20609_ (.A1(net1740),
    .A2(_12385_),
    .A3(_12387_),
    .B1(_12389_),
    .B2(net6216),
    .X(_12390_));
 sky130_fd_sc_hd__o221a_1 _20610_ (.A1(net1396),
    .A2(_12384_),
    .B1(_12388_),
    .B2(_12366_),
    .C1(_12390_),
    .X(_12391_));
 sky130_fd_sc_hd__xnor2_1 _20611_ (.A(net6217),
    .B(_12369_),
    .Y(_12392_));
 sky130_fd_sc_hd__nor3_1 _20612_ (.A(_12362_),
    .B(_12380_),
    .C(_12392_),
    .Y(_12393_));
 sky130_fd_sc_hd__o22a_1 _20613_ (.A1(net6766),
    .A2(net4038),
    .B1(_09055_),
    .B2(net3849),
    .X(_12394_));
 sky130_fd_sc_hd__mux2_1 _20614_ (.A0(net3854),
    .A1(net3852),
    .S(net2594),
    .X(_12395_));
 sky130_fd_sc_hd__o221a_1 _20615_ (.A1(net2601),
    .A2(_12394_),
    .B1(_12395_),
    .B2(net3325),
    .C1(_12353_),
    .X(_12396_));
 sky130_fd_sc_hd__or3b_1 _20616_ (.A(net1740),
    .B(_12367_),
    .C_N(net1396),
    .X(_12397_));
 sky130_fd_sc_hd__nand2_1 _20617_ (.A(net1226),
    .B(_12397_),
    .Y(_12398_));
 sky130_fd_sc_hd__xor2_1 _20618_ (.A(net1395),
    .B(_12398_),
    .X(_12399_));
 sky130_fd_sc_hd__o21a_1 _20619_ (.A1(_12391_),
    .A2(net707),
    .B1(_12399_),
    .X(_12400_));
 sky130_fd_sc_hd__or3_1 _20620_ (.A(_12399_),
    .B(_12391_),
    .C(net707),
    .X(_12401_));
 sky130_fd_sc_hd__and2b_1 _20621_ (.A_N(_12400_),
    .B(_12401_),
    .X(_12402_));
 sky130_fd_sc_hd__o21a_1 _20622_ (.A1(net2191),
    .A2(_12402_),
    .B1(net8054),
    .X(_12403_));
 sky130_fd_sc_hd__nand2_1 _20623_ (.A(net1494),
    .B(_12402_),
    .Y(_12404_));
 sky130_fd_sc_hd__mux2_1 _20624_ (.A0(_12403_),
    .A1(_12404_),
    .S(net6173),
    .X(_12405_));
 sky130_fd_sc_hd__clkbuf_1 _20625_ (.A(_12405_),
    .X(_00509_));
 sky130_fd_sc_hd__o21ai_1 _20626_ (.A1(net6173),
    .A2(_12400_),
    .B1(_12401_),
    .Y(_12406_));
 sky130_fd_sc_hd__mux2_1 _20627_ (.A0(net3848),
    .A1(net3847),
    .S(net2593),
    .X(_12407_));
 sky130_fd_sc_hd__mux2_1 _20628_ (.A0(net6755),
    .A1(_12407_),
    .S(net3305),
    .X(_12408_));
 sky130_fd_sc_hd__o21a_1 _20629_ (.A1(net1395),
    .A2(_12397_),
    .B1(_08992_),
    .X(_12409_));
 sky130_fd_sc_hd__xnor2_1 _20630_ (.A(net1739),
    .B(_12409_),
    .Y(_12410_));
 sky130_fd_sc_hd__and2b_1 _20631_ (.A_N(_12406_),
    .B(_12410_),
    .X(_12411_));
 sky130_fd_sc_hd__or2b_1 _20632_ (.A(_12410_),
    .B_N(_12406_),
    .X(_12412_));
 sky130_fd_sc_hd__and2b_1 _20633_ (.A_N(_12411_),
    .B(_12412_),
    .X(_12413_));
 sky130_fd_sc_hd__o21a_1 _20634_ (.A1(net2190),
    .A2(_12413_),
    .B1(net8054),
    .X(_12414_));
 sky130_fd_sc_hd__nand2_1 _20635_ (.A(net1495),
    .B(_12413_),
    .Y(_12415_));
 sky130_fd_sc_hd__mux2_1 _20636_ (.A0(_12414_),
    .A1(_12415_),
    .S(net6164),
    .X(_12416_));
 sky130_fd_sc_hd__clkbuf_1 _20637_ (.A(_12416_),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _20638_ (.A0(_12295_),
    .A1(net3846),
    .S(net2592),
    .X(_12417_));
 sky130_fd_sc_hd__mux2_1 _20639_ (.A0(net6755),
    .A1(_12417_),
    .S(net3305),
    .X(_12418_));
 sky130_fd_sc_hd__or3_1 _20640_ (.A(net1395),
    .B(_12397_),
    .C(net1739),
    .X(_12419_));
 sky130_fd_sc_hd__nand2_1 _20641_ (.A(_08992_),
    .B(_12419_),
    .Y(_12420_));
 sky130_fd_sc_hd__xor2_2 _20642_ (.A(net1738),
    .B(_12420_),
    .X(_12421_));
 sky130_fd_sc_hd__a21oi_1 _20643_ (.A1(net6164),
    .A2(_12412_),
    .B1(_12411_),
    .Y(_12422_));
 sky130_fd_sc_hd__xnor2_1 _20644_ (.A(_12421_),
    .B(_12422_),
    .Y(_12423_));
 sky130_fd_sc_hd__or2_1 _20645_ (.A(net2190),
    .B(_12423_),
    .X(_12424_));
 sky130_fd_sc_hd__a21oi_1 _20646_ (.A1(net1239),
    .A2(_12423_),
    .B1(net3147),
    .Y(_12425_));
 sky130_fd_sc_hd__a31o_1 _20647_ (.A1(net8058),
    .A2(net3147),
    .A3(_12424_),
    .B1(_12425_),
    .X(_00511_));
 sky130_fd_sc_hd__a22o_1 _20648_ (.A1(net6757),
    .A2(net2597),
    .B1(_09082_),
    .B2(net3124),
    .X(_12426_));
 sky130_fd_sc_hd__a22o_1 _20649_ (.A1(net6757),
    .A2(net3327),
    .B1(net2168),
    .B2(_12315_),
    .X(_12427_));
 sky130_fd_sc_hd__a21o_1 _20650_ (.A1(net6484),
    .A2(_12426_),
    .B1(_12427_),
    .X(_12428_));
 sky130_fd_sc_hd__or2_1 _20651_ (.A(net1738),
    .B(_12419_),
    .X(_12429_));
 sky130_fd_sc_hd__nand2_1 _20652_ (.A(net1077),
    .B(_12429_),
    .Y(_12430_));
 sky130_fd_sc_hd__xor2_1 _20653_ (.A(net1394),
    .B(_12430_),
    .X(_12431_));
 sky130_fd_sc_hd__nand2_1 _20654_ (.A(net6133),
    .B(_12421_),
    .Y(_12432_));
 sky130_fd_sc_hd__nor2_1 _20655_ (.A(net6132),
    .B(_12421_),
    .Y(_12433_));
 sky130_fd_sc_hd__a21oi_1 _20656_ (.A1(_12422_),
    .A2(_12432_),
    .B1(_12433_),
    .Y(_12434_));
 sky130_fd_sc_hd__and2_1 _20657_ (.A(_12431_),
    .B(_12434_),
    .X(_12435_));
 sky130_fd_sc_hd__nor2_1 _20658_ (.A(_12431_),
    .B(_12434_),
    .Y(_12436_));
 sky130_fd_sc_hd__nor2_1 _20659_ (.A(_12435_),
    .B(_12436_),
    .Y(_12437_));
 sky130_fd_sc_hd__o21a_1 _20660_ (.A1(net1837),
    .A2(_12437_),
    .B1(net8061),
    .X(_12438_));
 sky130_fd_sc_hd__or3b_1 _20661_ (.A(net3152),
    .B(net1816),
    .C_N(_12437_),
    .X(_12439_));
 sky130_fd_sc_hd__o21a_1 _20662_ (.A1(net6109),
    .A2(_12438_),
    .B1(_12439_),
    .X(_00512_));
 sky130_fd_sc_hd__or3_1 _20663_ (.A(net6502),
    .B(net3325),
    .C(net3850),
    .X(_12440_));
 sky130_fd_sc_hd__o21ai_1 _20664_ (.A1(net4039),
    .A2(net6757),
    .B1(_12440_),
    .Y(_12441_));
 sky130_fd_sc_hd__nand2_1 _20665_ (.A(net6483),
    .B(_12441_),
    .Y(_12442_));
 sky130_fd_sc_hd__o221a_1 _20666_ (.A1(net6755),
    .A2(net3305),
    .B1(_09143_),
    .B2(_12264_),
    .C1(_12442_),
    .X(_12443_));
 sky130_fd_sc_hd__o21a_1 _20667_ (.A1(net1394),
    .A2(_12429_),
    .B1(net1077),
    .X(_12444_));
 sky130_fd_sc_hd__xnor2_1 _20668_ (.A(_12443_),
    .B(_12444_),
    .Y(_12445_));
 sky130_fd_sc_hd__o21a_1 _20669_ (.A1(_12431_),
    .A2(_12434_),
    .B1(net6109),
    .X(_12446_));
 sky130_fd_sc_hd__or2_1 _20670_ (.A(_12435_),
    .B(_12446_),
    .X(_12447_));
 sky130_fd_sc_hd__xnor2_1 _20671_ (.A(_12445_),
    .B(_12447_),
    .Y(_12448_));
 sky130_fd_sc_hd__nand2_1 _20672_ (.A(net6091),
    .B(net1473),
    .Y(_12449_));
 sky130_fd_sc_hd__a21oi_1 _20673_ (.A1(net1473),
    .A2(_12448_),
    .B1(net3357),
    .Y(_12450_));
 sky130_fd_sc_hd__o22a_1 _20674_ (.A1(_12448_),
    .A2(_12449_),
    .B1(_12450_),
    .B2(net6091),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _20675_ (.A0(net6762),
    .A1(_12274_),
    .S(_09096_),
    .X(_12451_));
 sky130_fd_sc_hd__or3_1 _20676_ (.A(net1394),
    .B(_12429_),
    .C(_12443_),
    .X(_12452_));
 sky130_fd_sc_hd__nand2_1 _20677_ (.A(net1077),
    .B(_12452_),
    .Y(_12453_));
 sky130_fd_sc_hd__xor2_1 _20678_ (.A(_12451_),
    .B(_12453_),
    .X(_12454_));
 sky130_fd_sc_hd__and2_1 _20679_ (.A(net6091),
    .B(_12445_),
    .X(_12455_));
 sky130_fd_sc_hd__or2_1 _20680_ (.A(net6091),
    .B(_12445_),
    .X(_12456_));
 sky130_fd_sc_hd__o31a_1 _20681_ (.A1(_12435_),
    .A2(_12446_),
    .A3(_12455_),
    .B1(_12456_),
    .X(_12457_));
 sky130_fd_sc_hd__and2_1 _20682_ (.A(_12454_),
    .B(_12457_),
    .X(_12458_));
 sky130_fd_sc_hd__nor2_1 _20683_ (.A(_12454_),
    .B(_12457_),
    .Y(_12459_));
 sky130_fd_sc_hd__nor2_1 _20684_ (.A(_12458_),
    .B(_12459_),
    .Y(_12460_));
 sky130_fd_sc_hd__o21ai_1 _20685_ (.A1(net1403),
    .A2(_12460_),
    .B1(net8061),
    .Y(_12461_));
 sky130_fd_sc_hd__and3_1 _20686_ (.A(net6077),
    .B(net1496),
    .C(_12460_),
    .X(_12462_));
 sky130_fd_sc_hd__a21oi_1 _20687_ (.A1(net3143),
    .A2(_12461_),
    .B1(_12462_),
    .Y(_00514_));
 sky130_fd_sc_hd__mux2_2 _20688_ (.A0(net6762),
    .A1(_12295_),
    .S(_09096_),
    .X(_12463_));
 sky130_fd_sc_hd__or2_1 _20689_ (.A(_12451_),
    .B(_12452_),
    .X(_12464_));
 sky130_fd_sc_hd__nand2_1 _20690_ (.A(_08993_),
    .B(_12464_),
    .Y(_12465_));
 sky130_fd_sc_hd__xnor2_2 _20691_ (.A(_12463_),
    .B(_12465_),
    .Y(_12466_));
 sky130_fd_sc_hd__o21ba_1 _20692_ (.A1(net3143),
    .A2(_12459_),
    .B1_N(_12458_),
    .X(_12467_));
 sky130_fd_sc_hd__xor2_1 _20693_ (.A(_12466_),
    .B(_12467_),
    .X(_12468_));
 sky130_fd_sc_hd__o21ai_1 _20694_ (.A1(_12142_),
    .A2(_12468_),
    .B1(net8060),
    .Y(_12469_));
 sky130_fd_sc_hd__and3_1 _20695_ (.A(net6058),
    .B(net1496),
    .C(_12468_),
    .X(_12470_));
 sky130_fd_sc_hd__a21oi_1 _20696_ (.A1(net3132),
    .A2(_12469_),
    .B1(_12470_),
    .Y(_00515_));
 sky130_fd_sc_hd__a21o_1 _20697_ (.A1(_12466_),
    .A2(_12467_),
    .B1(net3132),
    .X(_12471_));
 sky130_fd_sc_hd__o21a_1 _20698_ (.A1(_12466_),
    .A2(_12467_),
    .B1(_12471_),
    .X(_12472_));
 sky130_fd_sc_hd__a22o_1 _20699_ (.A1(net6763),
    .A2(_09144_),
    .B1(_12313_),
    .B2(_09096_),
    .X(_12473_));
 sky130_fd_sc_hd__o21ai_1 _20700_ (.A1(_12463_),
    .A2(_12464_),
    .B1(_08993_),
    .Y(_12474_));
 sky130_fd_sc_hd__xor2_2 _20701_ (.A(_12473_),
    .B(_12474_),
    .X(_12475_));
 sky130_fd_sc_hd__xnor2_1 _20702_ (.A(_12472_),
    .B(_12475_),
    .Y(_12476_));
 sky130_fd_sc_hd__o21ai_1 _20703_ (.A1(_12142_),
    .A2(_12476_),
    .B1(net8060),
    .Y(_12477_));
 sky130_fd_sc_hd__and3_1 _20704_ (.A(net6056),
    .B(net1496),
    .C(_12476_),
    .X(_12478_));
 sky130_fd_sc_hd__a21oi_1 _20705_ (.A1(net3139),
    .A2(_12477_),
    .B1(_12478_),
    .Y(_00516_));
 sky130_fd_sc_hd__o31a_1 _20706_ (.A1(_12463_),
    .A2(_12464_),
    .A3(_12473_),
    .B1(_08993_),
    .X(_12479_));
 sky130_fd_sc_hd__mux2_1 _20707_ (.A0(net6763),
    .A1(_12269_),
    .S(net2583),
    .X(_12480_));
 sky130_fd_sc_hd__xnor2_2 _20708_ (.A(_12479_),
    .B(_12480_),
    .Y(_12481_));
 sky130_fd_sc_hd__nand2_1 _20709_ (.A(net6051),
    .B(_12475_),
    .Y(_12482_));
 sky130_fd_sc_hd__nor2_1 _20710_ (.A(net6051),
    .B(_12475_),
    .Y(_12483_));
 sky130_fd_sc_hd__a21o_1 _20711_ (.A1(_12472_),
    .A2(_12482_),
    .B1(_12483_),
    .X(_12484_));
 sky130_fd_sc_hd__xor2_1 _20712_ (.A(_12481_),
    .B(_12484_),
    .X(_12485_));
 sky130_fd_sc_hd__a21o_1 _20713_ (.A1(net2186),
    .A2(_12485_),
    .B1(_09023_),
    .X(_12486_));
 sky130_fd_sc_hd__or3_1 _20714_ (.A(net6023),
    .B(net2284),
    .C(_12485_),
    .X(_12487_));
 sky130_fd_sc_hd__a21bo_1 _20715_ (.A1(net6023),
    .A2(_12486_),
    .B1_N(_12487_),
    .X(_00517_));
 sky130_fd_sc_hd__xnor2_1 _20716_ (.A(net6764),
    .B(net5998),
    .Y(_12488_));
 sky130_fd_sc_hd__a21o_1 _20717_ (.A1(net2583),
    .A2(_12269_),
    .B1(_12479_),
    .X(_12489_));
 sky130_fd_sc_hd__nand2_1 _20718_ (.A(net966),
    .B(_12489_),
    .Y(_12490_));
 sky130_fd_sc_hd__xnor2_1 _20719_ (.A(_12488_),
    .B(_12490_),
    .Y(_12491_));
 sky130_fd_sc_hd__nand2_1 _20720_ (.A(net6023),
    .B(_12481_),
    .Y(_12492_));
 sky130_fd_sc_hd__and3_1 _20721_ (.A(_08915_),
    .B(_12482_),
    .C(_12492_),
    .X(_12493_));
 sky130_fd_sc_hd__nor2_1 _20722_ (.A(net6035),
    .B(_12481_),
    .Y(_12494_));
 sky130_fd_sc_hd__nor4_1 _20723_ (.A(net1817),
    .B(_12484_),
    .C(_12491_),
    .D(_12494_),
    .Y(_12495_));
 sky130_fd_sc_hd__a21oi_1 _20724_ (.A1(_12483_),
    .A2(_12492_),
    .B1(_12494_),
    .Y(_12496_));
 sky130_fd_sc_hd__mux2_1 _20725_ (.A0(_12492_),
    .A1(_12496_),
    .S(_12491_),
    .X(_12497_));
 sky130_fd_sc_hd__a2bb2o_1 _20726_ (.A1_N(net2284),
    .A2_N(_12497_),
    .B1(net4246),
    .B2(net5994),
    .X(_12498_));
 sky130_fd_sc_hd__a311o_1 _20727_ (.A1(_12472_),
    .A2(_12491_),
    .A3(_12493_),
    .B1(_12495_),
    .C1(_12498_),
    .X(_00518_));
 sky130_fd_sc_hd__o31a_1 _20728_ (.A1(net4390),
    .A2(net4346),
    .A3(net4324),
    .B1(net8906),
    .X(_12499_));
 sky130_fd_sc_hd__buf_1 _20729_ (.A(net3843),
    .X(_12500_));
 sky130_fd_sc_hd__inv_2 _20730_ (.A(_12499_),
    .Y(_12501_));
 sky130_fd_sc_hd__o31a_1 _20731_ (.A1(_04873_),
    .A2(_00005_),
    .A3(_00002_),
    .B1(_12501_),
    .X(_12502_));
 sky130_fd_sc_hd__clkbuf_1 _20732_ (.A(net2487),
    .X(_12503_));
 sky130_fd_sc_hd__nand2_1 _20733_ (.A(net5509),
    .B(net5867),
    .Y(_12504_));
 sky130_fd_sc_hd__nand2_1 _20734_ (.A(net5524),
    .B(net5838),
    .Y(_12505_));
 sky130_fd_sc_hd__nand2_1 _20735_ (.A(net5544),
    .B(net5810),
    .Y(_12506_));
 sky130_fd_sc_hd__xor2_1 _20736_ (.A(_12505_),
    .B(_12506_),
    .X(_12507_));
 sky130_fd_sc_hd__xnor2_2 _20737_ (.A(_12504_),
    .B(_12507_),
    .Y(_12508_));
 sky130_fd_sc_hd__nand2_1 _20738_ (.A(net5525),
    .B(net5867),
    .Y(_12509_));
 sky130_fd_sc_hd__nand2_1 _20739_ (.A(net5545),
    .B(net5838),
    .Y(_12510_));
 sky130_fd_sc_hd__nand2_1 _20740_ (.A(net5557),
    .B(net5823),
    .Y(_12511_));
 sky130_fd_sc_hd__o21a_1 _20741_ (.A1(_12509_),
    .A2(_12510_),
    .B1(_12511_),
    .X(_12512_));
 sky130_fd_sc_hd__a21o_1 _20742_ (.A1(_12509_),
    .A2(_12510_),
    .B1(_12512_),
    .X(_12513_));
 sky130_fd_sc_hd__nand2_2 _20743_ (.A(net5914),
    .B(net5473),
    .Y(_12514_));
 sky130_fd_sc_hd__nand2_2 _20744_ (.A(net5940),
    .B(net5454),
    .Y(_12515_));
 sky130_fd_sc_hd__nand2_1 _20745_ (.A(net5953),
    .B(net5424),
    .Y(_12516_));
 sky130_fd_sc_hd__xnor2_1 _20746_ (.A(_12515_),
    .B(_12516_),
    .Y(_12517_));
 sky130_fd_sc_hd__xnor2_2 _20747_ (.A(_12514_),
    .B(_12517_),
    .Y(_12518_));
 sky130_fd_sc_hd__xor2_1 _20748_ (.A(_12513_),
    .B(_12518_),
    .X(_12519_));
 sky130_fd_sc_hd__xnor2_2 _20749_ (.A(_12508_),
    .B(_12519_),
    .Y(_12520_));
 sky130_fd_sc_hd__nand2_1 _20750_ (.A(net5558),
    .B(net5836),
    .Y(_12521_));
 sky130_fd_sc_hd__nand2_1 _20751_ (.A(net5546),
    .B(net5873),
    .Y(_12522_));
 sky130_fd_sc_hd__nand2_1 _20752_ (.A(_12521_),
    .B(_12522_),
    .Y(_12523_));
 sky130_fd_sc_hd__nor2_1 _20753_ (.A(_12521_),
    .B(_12522_),
    .Y(_12524_));
 sky130_fd_sc_hd__a31o_1 _20754_ (.A1(net5579),
    .A2(net5822),
    .A3(_12523_),
    .B1(_12524_),
    .X(_12525_));
 sky130_fd_sc_hd__nand2_2 _20755_ (.A(net5931),
    .B(net5472),
    .Y(_12526_));
 sky130_fd_sc_hd__nand2_1 _20756_ (.A(net5491),
    .B(net5906),
    .Y(_12527_));
 sky130_fd_sc_hd__nand2_1 _20757_ (.A(net5954),
    .B(net5454),
    .Y(_12528_));
 sky130_fd_sc_hd__xnor2_1 _20758_ (.A(_12527_),
    .B(_12528_),
    .Y(_12529_));
 sky130_fd_sc_hd__xnor2_1 _20759_ (.A(_12526_),
    .B(_12529_),
    .Y(_12530_));
 sky130_fd_sc_hd__xnor2_1 _20760_ (.A(_12509_),
    .B(_12510_),
    .Y(_12531_));
 sky130_fd_sc_hd__xnor2_1 _20761_ (.A(_12511_),
    .B(_12531_),
    .Y(_12532_));
 sky130_fd_sc_hd__nor2_1 _20762_ (.A(_12530_),
    .B(net2485),
    .Y(_12533_));
 sky130_fd_sc_hd__nand2_1 _20763_ (.A(_12530_),
    .B(net2485),
    .Y(_12534_));
 sky130_fd_sc_hd__o21a_1 _20764_ (.A1(net2486),
    .A2(_12533_),
    .B1(_12534_),
    .X(_12535_));
 sky130_fd_sc_hd__xor2_2 _20765_ (.A(_12520_),
    .B(_12535_),
    .X(_12536_));
 sky130_fd_sc_hd__nand2_1 _20766_ (.A(net5612),
    .B(net5776),
    .Y(_12537_));
 sky130_fd_sc_hd__nand2_1 _20767_ (.A(net5596),
    .B(net5794),
    .Y(_12538_));
 sky130_fd_sc_hd__nand2_1 _20768_ (.A(net5627),
    .B(net5760),
    .Y(_12539_));
 sky130_fd_sc_hd__o21ai_1 _20769_ (.A1(_12537_),
    .A2(_12538_),
    .B1(_12539_),
    .Y(_12540_));
 sky130_fd_sc_hd__a21bo_1 _20770_ (.A1(_12537_),
    .A2(_12538_),
    .B1_N(_12540_),
    .X(_12541_));
 sky130_fd_sc_hd__nand2_1 _20771_ (.A(net5612),
    .B(net5760),
    .Y(_12542_));
 sky130_fd_sc_hd__nand2_1 _20772_ (.A(net5578),
    .B(net5794),
    .Y(_12543_));
 sky130_fd_sc_hd__nand2_1 _20773_ (.A(net5596),
    .B(net5776),
    .Y(_12544_));
 sky130_fd_sc_hd__xnor2_1 _20774_ (.A(_12543_),
    .B(_12544_),
    .Y(_12545_));
 sky130_fd_sc_hd__xnor2_1 _20775_ (.A(_12542_),
    .B(_12545_),
    .Y(_12546_));
 sky130_fd_sc_hd__or2_1 _20776_ (.A(_12541_),
    .B(_12546_),
    .X(_12547_));
 sky130_fd_sc_hd__nand2_2 _20777_ (.A(net5557),
    .B(net5795),
    .Y(_12548_));
 sky130_fd_sc_hd__nand2_1 _20778_ (.A(net5577),
    .B(net5774),
    .Y(_12549_));
 sky130_fd_sc_hd__nand2_1 _20779_ (.A(net5597),
    .B(net5761),
    .Y(_12550_));
 sky130_fd_sc_hd__xnor2_1 _20780_ (.A(_12549_),
    .B(_12550_),
    .Y(_12551_));
 sky130_fd_sc_hd__xnor2_2 _20781_ (.A(_12548_),
    .B(_12551_),
    .Y(_12552_));
 sky130_fd_sc_hd__nand4_1 _20782_ (.A(net5596),
    .B(net5578),
    .C(net5776),
    .D(net5794),
    .Y(_12553_));
 sky130_fd_sc_hd__a22oi_1 _20783_ (.A1(net5596),
    .A2(net5776),
    .B1(net5794),
    .B2(net5578),
    .Y(_12554_));
 sky130_fd_sc_hd__a21oi_1 _20784_ (.A1(_12542_),
    .A2(_12553_),
    .B1(_12554_),
    .Y(_12555_));
 sky130_fd_sc_hd__and2_1 _20785_ (.A(net5636),
    .B(net5625),
    .X(_12556_));
 sky130_fd_sc_hd__and3_1 _20786_ (.A(net5730),
    .B(net5740),
    .C(_12556_),
    .X(_12557_));
 sky130_fd_sc_hd__xnor2_1 _20787_ (.A(_12555_),
    .B(_12557_),
    .Y(_12558_));
 sky130_fd_sc_hd__xnor2_2 _20788_ (.A(_12552_),
    .B(_12558_),
    .Y(_12559_));
 sky130_fd_sc_hd__nand2_1 _20789_ (.A(net5615),
    .B(net5741),
    .Y(_12560_));
 sky130_fd_sc_hd__nand2_1 _20790_ (.A(net5626),
    .B(net5730),
    .Y(_12561_));
 sky130_fd_sc_hd__nand2_1 _20791_ (.A(net5637),
    .B(net5702),
    .Y(_12562_));
 sky130_fd_sc_hd__xnor2_1 _20792_ (.A(_12561_),
    .B(_12562_),
    .Y(_12563_));
 sky130_fd_sc_hd__xnor2_1 _20793_ (.A(_12560_),
    .B(_12563_),
    .Y(_00809_));
 sky130_fd_sc_hd__xnor2_2 _20794_ (.A(_12559_),
    .B(net2484),
    .Y(_00810_));
 sky130_fd_sc_hd__nand2_1 _20795_ (.A(net5627),
    .B(net5740),
    .Y(_00811_));
 sky130_fd_sc_hd__nand2_1 _20796_ (.A(net5635),
    .B(net5730),
    .Y(_00812_));
 sky130_fd_sc_hd__xor2_1 _20797_ (.A(_00811_),
    .B(_00812_),
    .X(_00813_));
 sky130_fd_sc_hd__a21bo_1 _20798_ (.A1(_12541_),
    .A2(_12546_),
    .B1_N(_00813_),
    .X(_00814_));
 sky130_fd_sc_hd__nand2_1 _20799_ (.A(_00810_),
    .B(_00814_),
    .Y(_00815_));
 sky130_fd_sc_hd__and2_1 _20800_ (.A(_12547_),
    .B(_00814_),
    .X(_00816_));
 sky130_fd_sc_hd__o21ai_1 _20801_ (.A1(_00810_),
    .A2(_00816_),
    .B1(_12536_),
    .Y(_00817_));
 sky130_fd_sc_hd__o211a_1 _20802_ (.A1(_12536_),
    .A2(_12547_),
    .B1(_00815_),
    .C1(_00817_),
    .X(_00818_));
 sky130_fd_sc_hd__nand2_1 _20803_ (.A(net5913),
    .B(net5455),
    .Y(_00819_));
 sky130_fd_sc_hd__nand2_2 _20804_ (.A(net5936),
    .B(net5425),
    .Y(_00820_));
 sky130_fd_sc_hd__nand2_1 _20805_ (.A(net5960),
    .B(net5414),
    .Y(_00821_));
 sky130_fd_sc_hd__xnor2_1 _20806_ (.A(_00820_),
    .B(_00821_),
    .Y(_00822_));
 sky130_fd_sc_hd__xnor2_1 _20807_ (.A(_00819_),
    .B(_00822_),
    .Y(_00823_));
 sky130_fd_sc_hd__o21ai_1 _20808_ (.A1(_12504_),
    .A2(_12505_),
    .B1(_12506_),
    .Y(_00824_));
 sky130_fd_sc_hd__a21bo_1 _20809_ (.A1(_12504_),
    .A2(_12505_),
    .B1_N(_00824_),
    .X(_00825_));
 sky130_fd_sc_hd__nand2_2 _20810_ (.A(net5861),
    .B(net5494),
    .Y(_00826_));
 sky130_fd_sc_hd__nand2_1 _20811_ (.A(net5830),
    .B(net5510),
    .Y(_00827_));
 sky130_fd_sc_hd__nand2_1 _20812_ (.A(net5810),
    .B(net5524),
    .Y(_00828_));
 sky130_fd_sc_hd__xnor2_1 _20813_ (.A(_00827_),
    .B(_00828_),
    .Y(_00829_));
 sky130_fd_sc_hd__xnor2_2 _20814_ (.A(_00826_),
    .B(_00829_),
    .Y(_00830_));
 sky130_fd_sc_hd__xnor2_1 _20815_ (.A(_00825_),
    .B(_00830_),
    .Y(_00831_));
 sky130_fd_sc_hd__xnor2_1 _20816_ (.A(_00823_),
    .B(_00831_),
    .Y(_00832_));
 sky130_fd_sc_hd__o21ba_1 _20817_ (.A1(_12513_),
    .A2(_12518_),
    .B1_N(_12508_),
    .X(_00833_));
 sky130_fd_sc_hd__a21oi_1 _20818_ (.A1(_12513_),
    .A2(_12518_),
    .B1(_00833_),
    .Y(_00834_));
 sky130_fd_sc_hd__o21ba_1 _20819_ (.A1(_12555_),
    .A2(_12557_),
    .B1_N(_12552_),
    .X(_00835_));
 sky130_fd_sc_hd__a21oi_1 _20820_ (.A1(_12555_),
    .A2(_12557_),
    .B1(_00835_),
    .Y(_00836_));
 sky130_fd_sc_hd__xor2_1 _20821_ (.A(_00834_),
    .B(net1736),
    .X(_00837_));
 sky130_fd_sc_hd__xnor2_2 _20822_ (.A(net1737),
    .B(_00837_),
    .Y(_00838_));
 sky130_fd_sc_hd__nor2_1 _20823_ (.A(_12559_),
    .B(net2484),
    .Y(_00839_));
 sky130_fd_sc_hd__nand2_2 _20824_ (.A(net5795),
    .B(net5544),
    .Y(_00840_));
 sky130_fd_sc_hd__nand2_1 _20825_ (.A(net5774),
    .B(net5570),
    .Y(_00841_));
 sky130_fd_sc_hd__nand2_1 _20826_ (.A(net5761),
    .B(net5577),
    .Y(_00842_));
 sky130_fd_sc_hd__xnor2_1 _20827_ (.A(_00841_),
    .B(_00842_),
    .Y(_00843_));
 sky130_fd_sc_hd__xnor2_2 _20828_ (.A(_00840_),
    .B(_00843_),
    .Y(_00844_));
 sky130_fd_sc_hd__o21a_1 _20829_ (.A1(_12560_),
    .A2(_12561_),
    .B1(_12562_),
    .X(_00845_));
 sky130_fd_sc_hd__a21o_1 _20830_ (.A1(_12560_),
    .A2(_12561_),
    .B1(_00845_),
    .X(_00846_));
 sky130_fd_sc_hd__o21a_1 _20831_ (.A1(_12548_),
    .A2(_12549_),
    .B1(_12550_),
    .X(_00847_));
 sky130_fd_sc_hd__a21o_1 _20832_ (.A1(_12548_),
    .A2(_12549_),
    .B1(_00847_),
    .X(_00848_));
 sky130_fd_sc_hd__xnor2_1 _20833_ (.A(net2483),
    .B(_00848_),
    .Y(_00849_));
 sky130_fd_sc_hd__xnor2_1 _20834_ (.A(_00844_),
    .B(_00849_),
    .Y(_00850_));
 sky130_fd_sc_hd__nand2_1 _20835_ (.A(net5687),
    .B(net5637),
    .Y(_00851_));
 sky130_fd_sc_hd__nand2_1 _20836_ (.A(net5741),
    .B(net5597),
    .Y(_00852_));
 sky130_fd_sc_hd__nand2_1 _20837_ (.A(net5731),
    .B(net5615),
    .Y(_00853_));
 sky130_fd_sc_hd__nand2_1 _20838_ (.A(net5702),
    .B(net5626),
    .Y(_00854_));
 sky130_fd_sc_hd__xnor2_1 _20839_ (.A(_00853_),
    .B(_00854_),
    .Y(_00855_));
 sky130_fd_sc_hd__xnor2_1 _20840_ (.A(_00852_),
    .B(_00855_),
    .Y(_00856_));
 sky130_fd_sc_hd__xnor2_1 _20841_ (.A(net3842),
    .B(_00856_),
    .Y(_00857_));
 sky130_fd_sc_hd__xnor2_1 _20842_ (.A(_00850_),
    .B(_00857_),
    .Y(_00858_));
 sky130_fd_sc_hd__xor2_1 _20843_ (.A(net1735),
    .B(net1393),
    .X(_00859_));
 sky130_fd_sc_hd__xnor2_2 _20844_ (.A(_00838_),
    .B(_00859_),
    .Y(_00860_));
 sky130_fd_sc_hd__o21bai_1 _20845_ (.A1(_12520_),
    .A2(_12547_),
    .B1_N(_12535_),
    .Y(_00861_));
 sky130_fd_sc_hd__a21bo_2 _20846_ (.A1(_12520_),
    .A2(_12547_),
    .B1_N(_00861_),
    .X(_00862_));
 sky130_fd_sc_hd__o21a_1 _20847_ (.A1(_12514_),
    .A2(_12515_),
    .B1(_12516_),
    .X(_00863_));
 sky130_fd_sc_hd__a21oi_2 _20848_ (.A1(_12514_),
    .A2(_12515_),
    .B1(_00863_),
    .Y(_00864_));
 sky130_fd_sc_hd__nand2_1 _20849_ (.A(_12526_),
    .B(_12528_),
    .Y(_00865_));
 sky130_fd_sc_hd__nor2_1 _20850_ (.A(_12526_),
    .B(_12528_),
    .Y(_00866_));
 sky130_fd_sc_hd__a21o_1 _20851_ (.A1(net5906),
    .A2(_00865_),
    .B1(_00866_),
    .X(_00867_));
 sky130_fd_sc_hd__nand2_1 _20852_ (.A(net5492),
    .B(_00867_),
    .Y(_00868_));
 sky130_fd_sc_hd__nand2_1 _20853_ (.A(net5473),
    .B(_00868_),
    .Y(_00869_));
 sky130_fd_sc_hd__or2_1 _20854_ (.A(net5473),
    .B(_00868_),
    .X(_00870_));
 sky130_fd_sc_hd__inv_2 _20855_ (.A(net5879),
    .Y(_00871_));
 sky130_fd_sc_hd__clkbuf_1 _20856_ (.A(net3840),
    .X(_00872_));
 sky130_fd_sc_hd__a21o_1 _20857_ (.A1(_00869_),
    .A2(_00870_),
    .B1(net3119),
    .X(_00873_));
 sky130_fd_sc_hd__xor2_1 _20858_ (.A(_00864_),
    .B(_00873_),
    .X(_00874_));
 sky130_fd_sc_hd__xnor2_2 _20859_ (.A(_00862_),
    .B(_00874_),
    .Y(_00875_));
 sky130_fd_sc_hd__xnor2_1 _20860_ (.A(_00860_),
    .B(_00875_),
    .Y(_00876_));
 sky130_fd_sc_hd__xnor2_2 _20861_ (.A(net1052),
    .B(_00876_),
    .Y(_00877_));
 sky130_fd_sc_hd__nand2_1 _20862_ (.A(net5642),
    .B(net5740),
    .Y(_00878_));
 sky130_fd_sc_hd__xnor2_1 _20863_ (.A(_12537_),
    .B(_12538_),
    .Y(_00879_));
 sky130_fd_sc_hd__xnor2_1 _20864_ (.A(_12539_),
    .B(_00879_),
    .Y(_00880_));
 sky130_fd_sc_hd__inv_2 _20865_ (.A(net5613),
    .Y(_00881_));
 sky130_fd_sc_hd__inv_2 _20866_ (.A(net5802),
    .Y(_00882_));
 sky130_fd_sc_hd__nand2_1 _20867_ (.A(net5627),
    .B(net5775),
    .Y(_00883_));
 sky130_fd_sc_hd__o21ai_1 _20868_ (.A1(_00881_),
    .A2(net3836),
    .B1(_00883_),
    .Y(_00884_));
 sky130_fd_sc_hd__and4_1 _20869_ (.A(net5627),
    .B(net5613),
    .C(net5775),
    .D(net5792),
    .X(_00885_));
 sky130_fd_sc_hd__a31oi_1 _20870_ (.A1(net5635),
    .A2(net5759),
    .A3(_00884_),
    .B1(_00885_),
    .Y(_00886_));
 sky130_fd_sc_hd__and2_1 _20871_ (.A(_00880_),
    .B(net2482),
    .X(_00887_));
 sky130_fd_sc_hd__xnor2_1 _20872_ (.A(_12541_),
    .B(_00813_),
    .Y(_00888_));
 sky130_fd_sc_hd__xnor2_1 _20873_ (.A(_12546_),
    .B(_00888_),
    .Y(_00889_));
 sky130_fd_sc_hd__o21bai_1 _20874_ (.A1(_00878_),
    .A2(_00887_),
    .B1_N(_00889_),
    .Y(_00890_));
 sky130_fd_sc_hd__or2_1 _20875_ (.A(_00880_),
    .B(net2482),
    .X(_00891_));
 sky130_fd_sc_hd__a21oi_1 _20876_ (.A1(_00891_),
    .A2(_00878_),
    .B1(_00887_),
    .Y(_00892_));
 sky130_fd_sc_hd__and2_1 _20877_ (.A(_00889_),
    .B(_00892_),
    .X(_00893_));
 sky130_fd_sc_hd__xor2_1 _20878_ (.A(net2486),
    .B(net2485),
    .X(_00894_));
 sky130_fd_sc_hd__xnor2_1 _20879_ (.A(_12530_),
    .B(_00894_),
    .Y(_00895_));
 sky130_fd_sc_hd__and2_1 _20880_ (.A(net5954),
    .B(net5472),
    .X(_00896_));
 sky130_fd_sc_hd__nand2_1 _20881_ (.A(net5507),
    .B(net5905),
    .Y(_00897_));
 sky130_fd_sc_hd__and2_1 _20882_ (.A(net5491),
    .B(net5935),
    .X(_00898_));
 sky130_fd_sc_hd__xnor2_1 _20883_ (.A(_00897_),
    .B(_00898_),
    .Y(_00899_));
 sky130_fd_sc_hd__xnor2_1 _20884_ (.A(_00896_),
    .B(_00899_),
    .Y(_00900_));
 sky130_fd_sc_hd__nand2_1 _20885_ (.A(net5575),
    .B(net5832),
    .Y(_00901_));
 sky130_fd_sc_hd__nand2_1 _20886_ (.A(net5558),
    .B(net5869),
    .Y(_00902_));
 sky130_fd_sc_hd__nand2_1 _20887_ (.A(net5601),
    .B(net5821),
    .Y(_00903_));
 sky130_fd_sc_hd__o21ai_1 _20888_ (.A1(_00901_),
    .A2(_00902_),
    .B1(_00903_),
    .Y(_00904_));
 sky130_fd_sc_hd__a21bo_1 _20889_ (.A1(_00901_),
    .A2(_00902_),
    .B1_N(_00904_),
    .X(_00905_));
 sky130_fd_sc_hd__or2_1 _20890_ (.A(_00900_),
    .B(net2481),
    .X(_00906_));
 sky130_fd_sc_hd__nand2_1 _20891_ (.A(net5579),
    .B(net5822),
    .Y(_00907_));
 sky130_fd_sc_hd__xnor2_1 _20892_ (.A(_12521_),
    .B(_12522_),
    .Y(_00908_));
 sky130_fd_sc_hd__xnor2_1 _20893_ (.A(_00907_),
    .B(_00908_),
    .Y(_00909_));
 sky130_fd_sc_hd__a21o_1 _20894_ (.A1(_00900_),
    .A2(net2481),
    .B1(_00909_),
    .X(_00910_));
 sky130_fd_sc_hd__nand2_1 _20895_ (.A(_00906_),
    .B(_00910_),
    .Y(_00911_));
 sky130_fd_sc_hd__xor2_1 _20896_ (.A(_00895_),
    .B(_00911_),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _20897_ (.A0(_00891_),
    .A1(_00893_),
    .S(_00912_),
    .X(_00913_));
 sky130_fd_sc_hd__a21o_1 _20898_ (.A1(_00906_),
    .A2(_00910_),
    .B1(_00891_),
    .X(_00914_));
 sky130_fd_sc_hd__and3_1 _20899_ (.A(_00906_),
    .B(_00910_),
    .C(_00891_),
    .X(_00915_));
 sky130_fd_sc_hd__a21o_1 _20900_ (.A1(_00895_),
    .A2(_00914_),
    .B1(_00915_),
    .X(_00916_));
 sky130_fd_sc_hd__inv_2 _20901_ (.A(net5513),
    .Y(_00917_));
 sky130_fd_sc_hd__nor2_1 _20902_ (.A(net3830),
    .B(net3840),
    .Y(_00918_));
 sky130_fd_sc_hd__o21a_1 _20903_ (.A1(net5906),
    .A2(_00896_),
    .B1(_00898_),
    .X(_00919_));
 sky130_fd_sc_hd__a21o_1 _20904_ (.A1(net5906),
    .A2(_00896_),
    .B1(_00919_),
    .X(_00920_));
 sky130_fd_sc_hd__and2_1 _20905_ (.A(_00918_),
    .B(_00920_),
    .X(_00921_));
 sky130_fd_sc_hd__a21o_1 _20906_ (.A1(net5906),
    .A2(_00865_),
    .B1(net5883),
    .X(_00922_));
 sky130_fd_sc_hd__a21oi_1 _20907_ (.A1(net5491),
    .A2(_00922_),
    .B1(_00866_),
    .Y(_00923_));
 sky130_fd_sc_hd__a31oi_2 _20908_ (.A1(net5492),
    .A2(net5883),
    .A3(_00867_),
    .B1(_00923_),
    .Y(_00924_));
 sky130_fd_sc_hd__xor2_1 _20909_ (.A(_00921_),
    .B(_00924_),
    .X(_00925_));
 sky130_fd_sc_hd__xnor2_1 _20910_ (.A(_00916_),
    .B(_00925_),
    .Y(_00926_));
 sky130_fd_sc_hd__a21oi_1 _20911_ (.A1(net1392),
    .A2(net1187),
    .B1(_00926_),
    .Y(_00927_));
 sky130_fd_sc_hd__xnor2_1 _20912_ (.A(_00810_),
    .B(_00816_),
    .Y(_00928_));
 sky130_fd_sc_hd__xnor2_1 _20913_ (.A(_12536_),
    .B(_00928_),
    .Y(_00929_));
 sky130_fd_sc_hd__and3_1 _20914_ (.A(_00926_),
    .B(net1392),
    .C(net1187),
    .X(_00930_));
 sky130_fd_sc_hd__o21ba_1 _20915_ (.A1(_00927_),
    .A2(net1186),
    .B1_N(_00930_),
    .X(_00931_));
 sky130_fd_sc_hd__o21ba_1 _20916_ (.A1(_00921_),
    .A2(_00924_),
    .B1_N(_00916_),
    .X(_00932_));
 sky130_fd_sc_hd__a21o_1 _20917_ (.A1(_00921_),
    .A2(_00924_),
    .B1(_00932_),
    .X(_00933_));
 sky130_fd_sc_hd__xor2_1 _20918_ (.A(_00931_),
    .B(_00933_),
    .X(_00934_));
 sky130_fd_sc_hd__xnor2_1 _20919_ (.A(_00877_),
    .B(_00934_),
    .Y(_00935_));
 sky130_fd_sc_hd__nand2_1 _20920_ (.A(net1392),
    .B(net1187),
    .Y(_00936_));
 sky130_fd_sc_hd__xor2_1 _20921_ (.A(_00926_),
    .B(net1186),
    .X(_00937_));
 sky130_fd_sc_hd__xnor2_2 _20922_ (.A(_00936_),
    .B(_00937_),
    .Y(_00938_));
 sky130_fd_sc_hd__nand2_2 _20923_ (.A(net5491),
    .B(net5954),
    .Y(_00939_));
 sky130_fd_sc_hd__nand2_1 _20924_ (.A(net5507),
    .B(net5935),
    .Y(_00940_));
 sky130_fd_sc_hd__nand2_1 _20925_ (.A(net5527),
    .B(net5905),
    .Y(_00941_));
 sky130_fd_sc_hd__o21ai_1 _20926_ (.A1(_00939_),
    .A2(_00940_),
    .B1(_00941_),
    .Y(_00942_));
 sky130_fd_sc_hd__a21boi_2 _20927_ (.A1(_00939_),
    .A2(_00940_),
    .B1_N(_00942_),
    .Y(_00943_));
 sky130_fd_sc_hd__and3_1 _20928_ (.A(net5527),
    .B(net5884),
    .C(_00943_),
    .X(_00944_));
 sky130_fd_sc_hd__nand2_1 _20929_ (.A(net5601),
    .B(net5832),
    .Y(_00945_));
 sky130_fd_sc_hd__nand2_1 _20930_ (.A(net5575),
    .B(net5869),
    .Y(_00946_));
 sky130_fd_sc_hd__nand2_1 _20931_ (.A(_00945_),
    .B(_00946_),
    .Y(_00947_));
 sky130_fd_sc_hd__nor2_1 _20932_ (.A(_00945_),
    .B(_00946_),
    .Y(_00948_));
 sky130_fd_sc_hd__a31o_1 _20933_ (.A1(net5621),
    .A2(net5821),
    .A3(_00947_),
    .B1(_00948_),
    .X(_00949_));
 sky130_fd_sc_hd__xor2_1 _20934_ (.A(_00901_),
    .B(_00902_),
    .X(_00950_));
 sky130_fd_sc_hd__xnor2_1 _20935_ (.A(_00903_),
    .B(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__or2_1 _20936_ (.A(_00949_),
    .B(_00951_),
    .X(_00952_));
 sky130_fd_sc_hd__xor2_1 _20937_ (.A(_00939_),
    .B(_00940_),
    .X(_00953_));
 sky130_fd_sc_hd__xnor2_1 _20938_ (.A(_00953_),
    .B(_00941_),
    .Y(_00954_));
 sky130_fd_sc_hd__a21o_1 _20939_ (.A1(_00949_),
    .A2(_00951_),
    .B1(_00954_),
    .X(_00955_));
 sky130_fd_sc_hd__nand2_1 _20940_ (.A(_00952_),
    .B(_00955_),
    .Y(_00956_));
 sky130_fd_sc_hd__xnor2_1 _20941_ (.A(_00900_),
    .B(net2481),
    .Y(_00957_));
 sky130_fd_sc_hd__xnor2_1 _20942_ (.A(_00909_),
    .B(_00957_),
    .Y(_00958_));
 sky130_fd_sc_hd__xnor2_1 _20943_ (.A(net5613),
    .B(net5759),
    .Y(_00959_));
 sky130_fd_sc_hd__and2_1 _20944_ (.A(net5779),
    .B(net5804),
    .X(_00960_));
 sky130_fd_sc_hd__and3_1 _20945_ (.A(_12556_),
    .B(_00959_),
    .C(net3825),
    .X(_00961_));
 sky130_fd_sc_hd__o21ba_1 _20946_ (.A1(_00956_),
    .A2(net1734),
    .B1_N(net3111),
    .X(_00962_));
 sky130_fd_sc_hd__a21oi_2 _20947_ (.A1(_00956_),
    .A2(net1734),
    .B1(_00962_),
    .Y(_00963_));
 sky130_fd_sc_hd__o21ai_1 _20948_ (.A1(_00896_),
    .A2(_00898_),
    .B1(net5905),
    .Y(_00964_));
 sky130_fd_sc_hd__mux2_1 _20949_ (.A0(_00920_),
    .A1(_00964_),
    .S(net3840),
    .X(_00965_));
 sky130_fd_sc_hd__o32a_1 _20950_ (.A1(_12526_),
    .A2(_00918_),
    .A3(_00939_),
    .B1(_00965_),
    .B2(net3830),
    .X(_00966_));
 sky130_fd_sc_hd__a21bo_1 _20951_ (.A1(_00944_),
    .A2(_00963_),
    .B1_N(_00966_),
    .X(_00967_));
 sky130_fd_sc_hd__o21ai_2 _20952_ (.A1(_00944_),
    .A2(_00963_),
    .B1(_00967_),
    .Y(_00968_));
 sky130_fd_sc_hd__and3b_1 _20953_ (.A_N(net5635),
    .B(net5613),
    .C(net5797),
    .X(_00969_));
 sky130_fd_sc_hd__a31o_1 _20954_ (.A1(net5635),
    .A2(net5759),
    .A3(net3836),
    .B1(_00969_),
    .X(_00970_));
 sky130_fd_sc_hd__a21o_1 _20955_ (.A1(net5613),
    .A2(net5792),
    .B1(net5635),
    .X(_00971_));
 sky130_fd_sc_hd__o21ai_1 _20956_ (.A1(net5759),
    .A2(net5792),
    .B1(_00971_),
    .Y(_00972_));
 sky130_fd_sc_hd__mux2_1 _20957_ (.A0(_00970_),
    .A1(_00972_),
    .S(_00883_),
    .X(_00973_));
 sky130_fd_sc_hd__a31o_1 _20958_ (.A1(net5635),
    .A2(net5793),
    .A3(_00959_),
    .B1(_00973_),
    .X(_00974_));
 sky130_fd_sc_hd__xnor2_1 _20959_ (.A(_00949_),
    .B(_00951_),
    .Y(_00975_));
 sky130_fd_sc_hd__xnor2_1 _20960_ (.A(_00954_),
    .B(_00975_),
    .Y(_00976_));
 sky130_fd_sc_hd__inv_2 _20961_ (.A(net5553),
    .Y(_00977_));
 sky130_fd_sc_hd__inv_4 _20962_ (.A(net5924),
    .Y(_00978_));
 sky130_fd_sc_hd__nor2_1 _20963_ (.A(net3823),
    .B(net3808),
    .Y(_00979_));
 sky130_fd_sc_hd__nand2_1 _20964_ (.A(net5528),
    .B(net5930),
    .Y(_00980_));
 sky130_fd_sc_hd__nand2_1 _20965_ (.A(net5506),
    .B(net5950),
    .Y(_00981_));
 sky130_fd_sc_hd__xor2_1 _20966_ (.A(_00980_),
    .B(_00981_),
    .X(_00982_));
 sky130_fd_sc_hd__xnor2_2 _20967_ (.A(_00979_),
    .B(_00982_),
    .Y(_00983_));
 sky130_fd_sc_hd__nand2_1 _20968_ (.A(net5621),
    .B(net5821),
    .Y(_00984_));
 sky130_fd_sc_hd__xnor2_1 _20969_ (.A(_00945_),
    .B(_00946_),
    .Y(_00985_));
 sky130_fd_sc_hd__xnor2_2 _20970_ (.A(_00984_),
    .B(_00985_),
    .Y(_00986_));
 sky130_fd_sc_hd__nand2_1 _20971_ (.A(net5621),
    .B(net5831),
    .Y(_00987_));
 sky130_fd_sc_hd__nand2_1 _20972_ (.A(net5602),
    .B(net5868),
    .Y(_00988_));
 sky130_fd_sc_hd__nand2_1 _20973_ (.A(_00987_),
    .B(_00988_),
    .Y(_00989_));
 sky130_fd_sc_hd__nor2_1 _20974_ (.A(_00987_),
    .B(_00988_),
    .Y(_00990_));
 sky130_fd_sc_hd__a31o_1 _20975_ (.A1(net5631),
    .A2(net5821),
    .A3(_00989_),
    .B1(_00990_),
    .X(_00991_));
 sky130_fd_sc_hd__o21bai_1 _20976_ (.A1(_00983_),
    .A2(_00986_),
    .B1_N(_00991_),
    .Y(_00992_));
 sky130_fd_sc_hd__a21bo_1 _20977_ (.A1(_00983_),
    .A2(_00986_),
    .B1_N(_00992_),
    .X(_00993_));
 sky130_fd_sc_hd__xor2_1 _20978_ (.A(_00976_),
    .B(_00993_),
    .X(_00994_));
 sky130_fd_sc_hd__or2_1 _20979_ (.A(net2076),
    .B(_00994_),
    .X(_00995_));
 sky130_fd_sc_hd__or2b_1 _20980_ (.A(_00993_),
    .B_N(_00976_),
    .X(_00996_));
 sky130_fd_sc_hd__nand2_1 _20981_ (.A(net5527),
    .B(net5884),
    .Y(_00997_));
 sky130_fd_sc_hd__xnor2_2 _20982_ (.A(_00997_),
    .B(_00943_),
    .Y(_00998_));
 sky130_fd_sc_hd__nor2_1 _20983_ (.A(_00980_),
    .B(_00981_),
    .Y(_00999_));
 sky130_fd_sc_hd__nand2_1 _20984_ (.A(_00980_),
    .B(_00981_),
    .Y(_01000_));
 sky130_fd_sc_hd__o21a_2 _20985_ (.A1(_00979_),
    .A2(_00999_),
    .B1(_01000_),
    .X(_01001_));
 sky130_fd_sc_hd__and3_1 _20986_ (.A(net5547),
    .B(net5884),
    .C(_01001_),
    .X(_01002_));
 sky130_fd_sc_hd__xnor2_1 _20987_ (.A(_00998_),
    .B(_01002_),
    .Y(_01003_));
 sky130_fd_sc_hd__xnor2_1 _20988_ (.A(_00996_),
    .B(_01003_),
    .Y(_01004_));
 sky130_fd_sc_hd__xor2_1 _20989_ (.A(net2482),
    .B(_00878_),
    .X(_01005_));
 sky130_fd_sc_hd__xnor2_1 _20990_ (.A(_00880_),
    .B(_01005_),
    .Y(_01006_));
 sky130_fd_sc_hd__nand3_2 _20991_ (.A(_00952_),
    .B(_00955_),
    .C(net3111),
    .Y(_01007_));
 sky130_fd_sc_hd__a21o_1 _20992_ (.A1(_00952_),
    .A2(_00955_),
    .B1(net3111),
    .X(_01008_));
 sky130_fd_sc_hd__nand3b_1 _20993_ (.A_N(net1734),
    .B(_01007_),
    .C(_01008_),
    .Y(_01009_));
 sky130_fd_sc_hd__a21bo_1 _20994_ (.A1(_01007_),
    .A2(_01008_),
    .B1_N(net1734),
    .X(_01010_));
 sky130_fd_sc_hd__nand3_1 _20995_ (.A(net1732),
    .B(_01009_),
    .C(_01010_),
    .Y(_01011_));
 sky130_fd_sc_hd__a21o_1 _20996_ (.A1(_01009_),
    .A2(_01010_),
    .B1(net1732),
    .X(_01012_));
 sky130_fd_sc_hd__nand2_1 _20997_ (.A(_01011_),
    .B(_01012_),
    .Y(_01013_));
 sky130_fd_sc_hd__o21a_1 _20998_ (.A1(_00995_),
    .A2(_01004_),
    .B1(net1051),
    .X(_01014_));
 sky130_fd_sc_hd__a21o_1 _20999_ (.A1(_00995_),
    .A2(_01004_),
    .B1(_01014_),
    .X(_01015_));
 sky130_fd_sc_hd__nand2_1 _21000_ (.A(_00998_),
    .B(_01002_),
    .Y(_01016_));
 sky130_fd_sc_hd__nor2_1 _21001_ (.A(_00998_),
    .B(_01002_),
    .Y(_01017_));
 sky130_fd_sc_hd__a21oi_1 _21002_ (.A1(_00996_),
    .A2(_01016_),
    .B1(_01017_),
    .Y(_01018_));
 sky130_fd_sc_hd__xor2_1 _21003_ (.A(_00889_),
    .B(_00892_),
    .X(_01019_));
 sky130_fd_sc_hd__xnor2_1 _21004_ (.A(_00912_),
    .B(_01019_),
    .Y(_01020_));
 sky130_fd_sc_hd__xnor2_1 _21005_ (.A(_01011_),
    .B(net1183),
    .Y(_01021_));
 sky130_fd_sc_hd__xnor2_1 _21006_ (.A(_00966_),
    .B(_00944_),
    .Y(_01022_));
 sky130_fd_sc_hd__xnor2_1 _21007_ (.A(_01022_),
    .B(_00963_),
    .Y(_01023_));
 sky130_fd_sc_hd__xnor2_2 _21008_ (.A(_01021_),
    .B(_01023_),
    .Y(_01024_));
 sky130_fd_sc_hd__nand2_1 _21009_ (.A(net1185),
    .B(_01024_),
    .Y(_01025_));
 sky130_fd_sc_hd__nor2_1 _21010_ (.A(net1185),
    .B(_01024_),
    .Y(_01026_));
 sky130_fd_sc_hd__a21oi_2 _21011_ (.A1(net862),
    .A2(_01025_),
    .B1(_01026_),
    .Y(_01027_));
 sky130_fd_sc_hd__xnor2_1 _21012_ (.A(_00995_),
    .B(_01004_),
    .Y(_01028_));
 sky130_fd_sc_hd__xnor2_2 _21013_ (.A(net1051),
    .B(_01028_),
    .Y(_01029_));
 sky130_fd_sc_hd__nand2_1 _21014_ (.A(net2076),
    .B(_00994_),
    .Y(_01030_));
 sky130_fd_sc_hd__nand2_1 _21015_ (.A(_00995_),
    .B(_01030_),
    .Y(_01031_));
 sky130_fd_sc_hd__nand2_1 _21016_ (.A(net5556),
    .B(net5910),
    .Y(_01032_));
 sky130_fd_sc_hd__nand2_1 _21017_ (.A(net5528),
    .B(net5950),
    .Y(_01033_));
 sky130_fd_sc_hd__nand2_1 _21018_ (.A(net5541),
    .B(net5930),
    .Y(_01034_));
 sky130_fd_sc_hd__xnor2_1 _21019_ (.A(_01033_),
    .B(_01034_),
    .Y(_01035_));
 sky130_fd_sc_hd__xnor2_1 _21020_ (.A(_01032_),
    .B(_01035_),
    .Y(_01036_));
 sky130_fd_sc_hd__nand2_1 _21021_ (.A(net5631),
    .B(net5831),
    .Y(_01037_));
 sky130_fd_sc_hd__nand2_1 _21022_ (.A(net5622),
    .B(net5868),
    .Y(_01038_));
 sky130_fd_sc_hd__and2_1 _21023_ (.A(net5640),
    .B(net5820),
    .X(_01039_));
 sky130_fd_sc_hd__o21bai_1 _21024_ (.A1(_01037_),
    .A2(_01038_),
    .B1_N(_01039_),
    .Y(_01040_));
 sky130_fd_sc_hd__a21bo_1 _21025_ (.A1(_01037_),
    .A2(_01038_),
    .B1_N(_01040_),
    .X(_01041_));
 sky130_fd_sc_hd__or2_1 _21026_ (.A(_01036_),
    .B(_01041_),
    .X(_01042_));
 sky130_fd_sc_hd__nand2_1 _21027_ (.A(net5631),
    .B(net5820),
    .Y(_01043_));
 sky130_fd_sc_hd__xnor2_1 _21028_ (.A(_00987_),
    .B(_00988_),
    .Y(_01044_));
 sky130_fd_sc_hd__xnor2_2 _21029_ (.A(_01043_),
    .B(_01044_),
    .Y(_01045_));
 sky130_fd_sc_hd__a21o_1 _21030_ (.A1(_01036_),
    .A2(_01041_),
    .B1(_01045_),
    .X(_01046_));
 sky130_fd_sc_hd__xor2_1 _21031_ (.A(_00991_),
    .B(_00983_),
    .X(_01047_));
 sky130_fd_sc_hd__xnor2_1 _21032_ (.A(_00986_),
    .B(_01047_),
    .Y(_01048_));
 sky130_fd_sc_hd__inv_2 _21033_ (.A(net5629),
    .Y(_01049_));
 sky130_fd_sc_hd__o211a_1 _21034_ (.A1(_01049_),
    .A2(net3836),
    .B1(net5775),
    .C1(net5635),
    .X(_01050_));
 sky130_fd_sc_hd__a211o_1 _21035_ (.A1(net5641),
    .A2(net5775),
    .B1(net3836),
    .C1(_01049_),
    .X(_01051_));
 sky130_fd_sc_hd__and2b_1 _21036_ (.A_N(_01050_),
    .B(_01051_),
    .X(_01052_));
 sky130_fd_sc_hd__a22o_1 _21037_ (.A1(net5528),
    .A2(net5950),
    .B1(net5930),
    .B2(net5910),
    .X(_01053_));
 sky130_fd_sc_hd__or2_1 _21038_ (.A(net5929),
    .B(net5911),
    .X(_01054_));
 sky130_fd_sc_hd__a31o_1 _21039_ (.A1(net5556),
    .A2(_01053_),
    .A3(net3806),
    .B1(net3823),
    .X(_01055_));
 sky130_fd_sc_hd__or3_1 _21040_ (.A(net5541),
    .B(_01032_),
    .C(_01033_),
    .X(_01056_));
 sky130_fd_sc_hd__a21oi_1 _21041_ (.A1(_01055_),
    .A2(_01056_),
    .B1(net3841),
    .Y(_01057_));
 sky130_fd_sc_hd__xnor2_2 _21042_ (.A(_01001_),
    .B(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hd__a311o_1 _21043_ (.A1(net2075),
    .A2(net2074),
    .A3(net1731),
    .B1(net2480),
    .C1(_01058_),
    .X(_01059_));
 sky130_fd_sc_hd__a21oi_1 _21044_ (.A1(net2075),
    .A2(net2074),
    .B1(net1731),
    .Y(_01060_));
 sky130_fd_sc_hd__a21o_1 _21045_ (.A1(net2075),
    .A2(net2074),
    .B1(net2480),
    .X(_01061_));
 sky130_fd_sc_hd__and3_1 _21046_ (.A(net2075),
    .B(net2074),
    .C(net2480),
    .X(_01062_));
 sky130_fd_sc_hd__a21o_1 _21047_ (.A1(net1731),
    .A2(_01061_),
    .B1(_01062_),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _21048_ (.A0(_01060_),
    .A1(_01063_),
    .S(_01058_),
    .X(_01064_));
 sky130_fd_sc_hd__a21o_1 _21049_ (.A1(_01031_),
    .A2(_01059_),
    .B1(_01064_),
    .X(_01065_));
 sky130_fd_sc_hd__inv_2 _21050_ (.A(net5567),
    .Y(_01066_));
 sky130_fd_sc_hd__o21a_1 _21051_ (.A1(_01033_),
    .A2(_01034_),
    .B1(_01032_),
    .X(_01067_));
 sky130_fd_sc_hd__a21o_1 _21052_ (.A1(_01033_),
    .A2(_01034_),
    .B1(_01067_),
    .X(_01068_));
 sky130_fd_sc_hd__or2_1 _21053_ (.A(net3805),
    .B(_01068_),
    .X(_01069_));
 sky130_fd_sc_hd__and2b_1 _21054_ (.A_N(_01060_),
    .B(_01069_),
    .X(_01070_));
 sky130_fd_sc_hd__a21oi_1 _21055_ (.A1(net3823),
    .A2(_01001_),
    .B1(_01060_),
    .Y(_01071_));
 sky130_fd_sc_hd__o32a_1 _21056_ (.A1(net3823),
    .A2(_01001_),
    .A3(_01070_),
    .B1(_01071_),
    .B2(_01069_),
    .X(_01072_));
 sky130_fd_sc_hd__o211a_1 _21057_ (.A1(net3823),
    .A2(net3121),
    .B1(_01060_),
    .C1(_01001_),
    .X(_01073_));
 sky130_fd_sc_hd__o21ba_1 _21058_ (.A1(net3121),
    .A2(_01072_),
    .B1_N(_01073_),
    .X(_01074_));
 sky130_fd_sc_hd__a21o_1 _21059_ (.A1(_01029_),
    .A2(_01065_),
    .B1(_01074_),
    .X(_01075_));
 sky130_fd_sc_hd__o21ai_1 _21060_ (.A1(_01029_),
    .A2(_01065_),
    .B1(_01075_),
    .Y(_01076_));
 sky130_fd_sc_hd__xor2_1 _21061_ (.A(net1185),
    .B(_01024_),
    .X(_01077_));
 sky130_fd_sc_hd__xnor2_1 _21062_ (.A(net862),
    .B(_01077_),
    .Y(_01078_));
 sky130_fd_sc_hd__nand2_1 _21063_ (.A(net5581),
    .B(net5911),
    .Y(_01079_));
 sky130_fd_sc_hd__nand2_1 _21064_ (.A(net5552),
    .B(net5949),
    .Y(_01080_));
 sky130_fd_sc_hd__nand2_1 _21065_ (.A(net5564),
    .B(net5929),
    .Y(_01081_));
 sky130_fd_sc_hd__xor2_1 _21066_ (.A(_01080_),
    .B(_01081_),
    .X(_01082_));
 sky130_fd_sc_hd__xnor2_2 _21067_ (.A(_01079_),
    .B(_01082_),
    .Y(_01083_));
 sky130_fd_sc_hd__and3_1 _21068_ (.A(net5835),
    .B(net5871),
    .C(_12556_),
    .X(_01084_));
 sky130_fd_sc_hd__xnor2_1 _21069_ (.A(_01037_),
    .B(_01038_),
    .Y(_01085_));
 sky130_fd_sc_hd__xnor2_1 _21070_ (.A(_01039_),
    .B(_01085_),
    .Y(_01086_));
 sky130_fd_sc_hd__o21a_1 _21071_ (.A1(_01083_),
    .A2(_01084_),
    .B1(_01086_),
    .X(_01087_));
 sky130_fd_sc_hd__a21o_1 _21072_ (.A1(_01083_),
    .A2(_01084_),
    .B1(_01087_),
    .X(_01088_));
 sky130_fd_sc_hd__xor2_1 _21073_ (.A(_01036_),
    .B(_01041_),
    .X(_01089_));
 sky130_fd_sc_hd__xnor2_2 _21074_ (.A(_01045_),
    .B(_01089_),
    .Y(_01090_));
 sky130_fd_sc_hd__o21a_1 _21075_ (.A1(_01080_),
    .A2(_01081_),
    .B1(_01079_),
    .X(_01091_));
 sky130_fd_sc_hd__a21oi_2 _21076_ (.A1(_01080_),
    .A2(_01081_),
    .B1(_01091_),
    .Y(_01092_));
 sky130_fd_sc_hd__and2_1 _21077_ (.A(net5581),
    .B(_01092_),
    .X(_01093_));
 sky130_fd_sc_hd__a21o_1 _21078_ (.A1(_01088_),
    .A2(_01090_),
    .B1(_01093_),
    .X(_01094_));
 sky130_fd_sc_hd__nand2_1 _21079_ (.A(_01088_),
    .B(_01090_),
    .Y(_01095_));
 sky130_fd_sc_hd__o21ai_1 _21080_ (.A1(net5556),
    .A2(_01068_),
    .B1(_01095_),
    .Y(_01096_));
 sky130_fd_sc_hd__a32o_1 _21081_ (.A1(net5556),
    .A2(_01068_),
    .A3(_01094_),
    .B1(_01096_),
    .B2(_01093_),
    .X(_01097_));
 sky130_fd_sc_hd__a211o_1 _21082_ (.A1(net5562),
    .A2(net5879),
    .B1(_01095_),
    .C1(_01068_),
    .X(_01098_));
 sky130_fd_sc_hd__a21bo_1 _21083_ (.A1(net5879),
    .A2(_01097_),
    .B1_N(_01098_),
    .X(_01099_));
 sky130_fd_sc_hd__xor2_2 _21084_ (.A(_01088_),
    .B(_01090_),
    .X(_01100_));
 sky130_fd_sc_hd__a21oi_1 _21085_ (.A1(net2075),
    .A2(net2074),
    .B1(net2480),
    .Y(_01101_));
 sky130_fd_sc_hd__o21ba_1 _21086_ (.A1(_01101_),
    .A2(_01062_),
    .B1_N(net1731),
    .X(_01102_));
 sky130_fd_sc_hd__and3b_1 _21087_ (.A_N(_01062_),
    .B(net1731),
    .C(_01061_),
    .X(_01103_));
 sky130_fd_sc_hd__a311o_1 _21088_ (.A1(net5642),
    .A2(net5793),
    .A3(_01100_),
    .B1(_01102_),
    .C1(_01103_),
    .X(_01104_));
 sky130_fd_sc_hd__a22o_1 _21089_ (.A1(net5552),
    .A2(net5949),
    .B1(net5929),
    .B2(net5904),
    .X(_01105_));
 sky130_fd_sc_hd__a31o_1 _21090_ (.A1(net5581),
    .A2(_01054_),
    .A3(_01105_),
    .B1(net3805),
    .X(_01106_));
 sky130_fd_sc_hd__or3_1 _21091_ (.A(net5564),
    .B(_01079_),
    .C(_01080_),
    .X(_01107_));
 sky130_fd_sc_hd__a21oi_1 _21092_ (.A1(_01106_),
    .A2(_01107_),
    .B1(_00871_),
    .Y(_01108_));
 sky130_fd_sc_hd__xnor2_1 _21093_ (.A(_01068_),
    .B(_01108_),
    .Y(_01109_));
 sky130_fd_sc_hd__xnor2_1 _21094_ (.A(_01095_),
    .B(_01109_),
    .Y(_01110_));
 sky130_fd_sc_hd__o2111ai_2 _21095_ (.A1(_01103_),
    .A2(_01102_),
    .B1(_01100_),
    .C1(net5793),
    .D1(net5642),
    .Y(_01111_));
 sky130_fd_sc_hd__a21bo_1 _21096_ (.A1(_01104_),
    .A2(_01110_),
    .B1_N(_01111_),
    .X(_01112_));
 sky130_fd_sc_hd__xnor2_1 _21097_ (.A(_01063_),
    .B(_01058_),
    .Y(_01113_));
 sky130_fd_sc_hd__xnor2_1 _21098_ (.A(_01031_),
    .B(_01113_),
    .Y(_01114_));
 sky130_fd_sc_hd__a21boi_1 _21099_ (.A1(_01099_),
    .A2(_01112_),
    .B1_N(_01114_),
    .Y(_01115_));
 sky130_fd_sc_hd__nor2_1 _21100_ (.A(_01099_),
    .B(_01112_),
    .Y(_01116_));
 sky130_fd_sc_hd__nand2_1 _21101_ (.A(net5564),
    .B(net5949),
    .Y(_01117_));
 sky130_fd_sc_hd__nand2_1 _21102_ (.A(net5581),
    .B(net5929),
    .Y(_01118_));
 sky130_fd_sc_hd__nand2_2 _21103_ (.A(net5607),
    .B(net5911),
    .Y(_01119_));
 sky130_fd_sc_hd__o21a_1 _21104_ (.A1(_01117_),
    .A2(_01118_),
    .B1(_01119_),
    .X(_01120_));
 sky130_fd_sc_hd__a21oi_1 _21105_ (.A1(_01117_),
    .A2(_01118_),
    .B1(_01120_),
    .Y(_01121_));
 sky130_fd_sc_hd__and3_1 _21106_ (.A(net5605),
    .B(net5880),
    .C(_01121_),
    .X(_01122_));
 sky130_fd_sc_hd__nand2_1 _21107_ (.A(net5584),
    .B(net5880),
    .Y(_01123_));
 sky130_fd_sc_hd__xnor2_1 _21108_ (.A(_01092_),
    .B(_01123_),
    .Y(_01124_));
 sky130_fd_sc_hd__xnor2_1 _21109_ (.A(_01117_),
    .B(_01118_),
    .Y(_01125_));
 sky130_fd_sc_hd__xnor2_2 _21110_ (.A(_01119_),
    .B(_01125_),
    .Y(_01126_));
 sky130_fd_sc_hd__nand2_1 _21111_ (.A(net5630),
    .B(net5870),
    .Y(_01127_));
 sky130_fd_sc_hd__nand2_1 _21112_ (.A(net5644),
    .B(net5833),
    .Y(_01128_));
 sky130_fd_sc_hd__xor2_2 _21113_ (.A(_01127_),
    .B(_01128_),
    .X(_01129_));
 sky130_fd_sc_hd__or2b_1 _21114_ (.A(_01126_),
    .B_N(_01129_),
    .X(_01130_));
 sky130_fd_sc_hd__xnor2_1 _21115_ (.A(_01086_),
    .B(_01083_),
    .Y(_01131_));
 sky130_fd_sc_hd__xnor2_1 _21116_ (.A(_01084_),
    .B(_01131_),
    .Y(_01132_));
 sky130_fd_sc_hd__and2b_1 _21117_ (.A_N(_01130_),
    .B(_01132_),
    .X(_01133_));
 sky130_fd_sc_hd__a22o_1 _21118_ (.A1(net5564),
    .A2(net5949),
    .B1(net5929),
    .B2(net5911),
    .X(_01134_));
 sky130_fd_sc_hd__inv_2 _21119_ (.A(net5585),
    .Y(_01135_));
 sky130_fd_sc_hd__a31o_1 _21120_ (.A1(net5603),
    .A2(_01054_),
    .A3(_01134_),
    .B1(_01135_),
    .X(_01136_));
 sky130_fd_sc_hd__or3_1 _21121_ (.A(net5584),
    .B(_01119_),
    .C(_01117_),
    .X(_01137_));
 sky130_fd_sc_hd__a21oi_1 _21122_ (.A1(_01136_),
    .A2(_01137_),
    .B1(_00871_),
    .Y(_01138_));
 sky130_fd_sc_hd__xnor2_1 _21123_ (.A(_01092_),
    .B(_01138_),
    .Y(_01139_));
 sky130_fd_sc_hd__xnor2_1 _21124_ (.A(_01133_),
    .B(_01139_),
    .Y(_01140_));
 sky130_fd_sc_hd__nand2_1 _21125_ (.A(net5643),
    .B(net5796),
    .Y(_01141_));
 sky130_fd_sc_hd__xnor2_1 _21126_ (.A(_01141_),
    .B(_01100_),
    .Y(_01142_));
 sky130_fd_sc_hd__and2b_1 _21127_ (.A_N(_01139_),
    .B(_01133_),
    .X(_01143_));
 sky130_fd_sc_hd__a221o_1 _21128_ (.A1(_01122_),
    .A2(_01124_),
    .B1(_01140_),
    .B2(_01142_),
    .C1(_01143_),
    .X(_01144_));
 sky130_fd_sc_hd__and3_1 _21129_ (.A(_01104_),
    .B(_01111_),
    .C(_01110_),
    .X(_01145_));
 sky130_fd_sc_hd__a21oi_1 _21130_ (.A1(_01104_),
    .A2(_01111_),
    .B1(_01110_),
    .Y(_01146_));
 sky130_fd_sc_hd__nor2_1 _21131_ (.A(_01145_),
    .B(_01146_),
    .Y(_01147_));
 sky130_fd_sc_hd__xor2_1 _21132_ (.A(_01130_),
    .B(_01132_),
    .X(_01148_));
 sky130_fd_sc_hd__nand2_1 _21133_ (.A(net5614),
    .B(net5908),
    .Y(_01149_));
 sky130_fd_sc_hd__nand2_1 _21134_ (.A(net5583),
    .B(net5952),
    .Y(_01150_));
 sky130_fd_sc_hd__nand2_2 _21135_ (.A(net5603),
    .B(net5932),
    .Y(_01151_));
 sky130_fd_sc_hd__xnor2_1 _21136_ (.A(_01150_),
    .B(_01151_),
    .Y(_01152_));
 sky130_fd_sc_hd__xnor2_1 _21137_ (.A(_01149_),
    .B(_01152_),
    .Y(_01153_));
 sky130_fd_sc_hd__nand2_1 _21138_ (.A(net5634),
    .B(net5872),
    .Y(_01154_));
 sky130_fd_sc_hd__or2_1 _21139_ (.A(_01153_),
    .B(_01154_),
    .X(_01155_));
 sky130_fd_sc_hd__xor2_2 _21140_ (.A(_01126_),
    .B(_01129_),
    .X(_01156_));
 sky130_fd_sc_hd__nor2_1 _21141_ (.A(net2073),
    .B(_01156_),
    .Y(_01157_));
 sky130_fd_sc_hd__a21oi_1 _21142_ (.A1(net3816),
    .A2(_01151_),
    .B1(_01150_),
    .Y(_01158_));
 sky130_fd_sc_hd__nor2_1 _21143_ (.A(net3816),
    .B(_01151_),
    .Y(_01159_));
 sky130_fd_sc_hd__nand2_1 _21144_ (.A(net5617),
    .B(net5881),
    .Y(_01160_));
 sky130_fd_sc_hd__o21ba_1 _21145_ (.A1(_01158_),
    .A2(_01159_),
    .B1_N(_01160_),
    .X(_01161_));
 sky130_fd_sc_hd__nand2_1 _21146_ (.A(net5605),
    .B(net5880),
    .Y(_01162_));
 sky130_fd_sc_hd__xnor2_1 _21147_ (.A(_01121_),
    .B(_01162_),
    .Y(_01163_));
 sky130_fd_sc_hd__xnor2_1 _21148_ (.A(_01161_),
    .B(_01163_),
    .Y(_01164_));
 sky130_fd_sc_hd__xnor2_1 _21149_ (.A(_01157_),
    .B(_01164_),
    .Y(_01165_));
 sky130_fd_sc_hd__xnor2_1 _21150_ (.A(_01148_),
    .B(_01165_),
    .Y(_01166_));
 sky130_fd_sc_hd__xor2_1 _21151_ (.A(_01153_),
    .B(_01154_),
    .X(_01167_));
 sky130_fd_sc_hd__nand2_1 _21152_ (.A(net5618),
    .B(net5937),
    .Y(_01168_));
 sky130_fd_sc_hd__nand2_1 _21153_ (.A(net5599),
    .B(net5955),
    .Y(_01169_));
 sky130_fd_sc_hd__nand2_1 _21154_ (.A(net5628),
    .B(net5912),
    .Y(_01170_));
 sky130_fd_sc_hd__xor2_1 _21155_ (.A(_01169_),
    .B(_01170_),
    .X(_01171_));
 sky130_fd_sc_hd__xnor2_1 _21156_ (.A(_01168_),
    .B(_01171_),
    .Y(_01172_));
 sky130_fd_sc_hd__a22o_1 _21157_ (.A1(net5611),
    .A2(net5948),
    .B1(net5928),
    .B2(net5629),
    .X(_01173_));
 sky130_fd_sc_hd__and2_1 _21158_ (.A(net5956),
    .B(net5937),
    .X(_01174_));
 sky130_fd_sc_hd__a32o_1 _21159_ (.A1(net5625),
    .A2(net5611),
    .A3(_01174_),
    .B1(net5916),
    .B2(net5641),
    .X(_01175_));
 sky130_fd_sc_hd__nand2_1 _21160_ (.A(_01173_),
    .B(_01175_),
    .Y(_01176_));
 sky130_fd_sc_hd__or2_1 _21161_ (.A(net5611),
    .B(net5916),
    .X(_01177_));
 sky130_fd_sc_hd__nand2_1 _21162_ (.A(_01174_),
    .B(_12556_),
    .Y(_01178_));
 sky130_fd_sc_hd__a21o_1 _21163_ (.A1(_01149_),
    .A2(_01177_),
    .B1(_01178_),
    .X(_01179_));
 sky130_fd_sc_hd__nor2_1 _21164_ (.A(_01176_),
    .B(_01179_),
    .Y(_01180_));
 sky130_fd_sc_hd__or2_1 _21165_ (.A(_01168_),
    .B(_01169_),
    .X(_01181_));
 sky130_fd_sc_hd__nand2_1 _21166_ (.A(net5882),
    .B(_01181_),
    .Y(_01182_));
 sky130_fd_sc_hd__a21o_1 _21167_ (.A1(_01168_),
    .A2(_01169_),
    .B1(net3816),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _21168_ (.A0(net5882),
    .A1(_01182_),
    .S(_01183_),
    .X(_01184_));
 sky130_fd_sc_hd__a21o_1 _21169_ (.A1(net5628),
    .A2(net5882),
    .B1(_01181_),
    .X(_01185_));
 sky130_fd_sc_hd__o21ai_1 _21170_ (.A1(net3807),
    .A2(_01184_),
    .B1(_01185_),
    .Y(_01186_));
 sky130_fd_sc_hd__a41o_1 _21171_ (.A1(net5634),
    .A2(net5882),
    .A3(_01172_),
    .A4(_01180_),
    .B1(_01186_),
    .X(_01187_));
 sky130_fd_sc_hd__xor2_2 _21172_ (.A(net2073),
    .B(_01156_),
    .X(_01188_));
 sky130_fd_sc_hd__a21oi_1 _21173_ (.A1(_01181_),
    .A2(_01183_),
    .B1(net3807),
    .Y(_01189_));
 sky130_fd_sc_hd__xnor2_1 _21174_ (.A(net3839),
    .B(_01189_),
    .Y(_01190_));
 sky130_fd_sc_hd__nand2_1 _21175_ (.A(net5881),
    .B(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__nand2_1 _21176_ (.A(_01150_),
    .B(_01151_),
    .Y(_01192_));
 sky130_fd_sc_hd__nor2_1 _21177_ (.A(_01150_),
    .B(_01151_),
    .Y(_01193_));
 sky130_fd_sc_hd__a31o_1 _21178_ (.A1(net5619),
    .A2(net5909),
    .A3(_01192_),
    .B1(_01193_),
    .X(_01194_));
 sky130_fd_sc_hd__inv_2 _21179_ (.A(_01194_),
    .Y(_01195_));
 sky130_fd_sc_hd__xnor2_1 _21180_ (.A(_01191_),
    .B(_01195_),
    .Y(_01196_));
 sky130_fd_sc_hd__xnor2_1 _21181_ (.A(_01188_),
    .B(_01196_),
    .Y(_01197_));
 sky130_fd_sc_hd__nand2_1 _21182_ (.A(_01176_),
    .B(_01179_),
    .Y(_01198_));
 sky130_fd_sc_hd__a31o_1 _21183_ (.A1(net5634),
    .A2(net5882),
    .A3(_01172_),
    .B1(_01198_),
    .X(_01199_));
 sky130_fd_sc_hd__a211o_1 _21184_ (.A1(net5638),
    .A2(net5878),
    .B1(_01172_),
    .C1(_01180_),
    .X(_01200_));
 sky130_fd_sc_hd__a22o_1 _21185_ (.A1(_01167_),
    .A2(_01186_),
    .B1(_01199_),
    .B2(_01200_),
    .X(_01201_));
 sky130_fd_sc_hd__o211a_1 _21186_ (.A1(_01167_),
    .A2(_01187_),
    .B1(_01197_),
    .C1(_01201_),
    .X(_01202_));
 sky130_fd_sc_hd__a21bo_1 _21187_ (.A1(_01157_),
    .A2(_01161_),
    .B1_N(_01148_),
    .X(_01203_));
 sky130_fd_sc_hd__o21a_1 _21188_ (.A1(_01157_),
    .A2(_01161_),
    .B1(_01203_),
    .X(_01204_));
 sky130_fd_sc_hd__or3b_1 _21189_ (.A(_01157_),
    .B(_01161_),
    .C_N(_01148_),
    .X(_01205_));
 sky130_fd_sc_hd__o21a_1 _21190_ (.A1(_01163_),
    .A2(_01204_),
    .B1(_01205_),
    .X(_01206_));
 sky130_fd_sc_hd__xor2_1 _21191_ (.A(_01142_),
    .B(_01140_),
    .X(_01207_));
 sky130_fd_sc_hd__or2_1 _21192_ (.A(_01189_),
    .B(_01188_),
    .X(_01208_));
 sky130_fd_sc_hd__a21o_1 _21193_ (.A1(net3839),
    .A2(_01194_),
    .B1(_01188_),
    .X(_01209_));
 sky130_fd_sc_hd__a32o_1 _21194_ (.A1(net5617),
    .A2(_01195_),
    .A3(_01208_),
    .B1(_01209_),
    .B2(_01189_),
    .X(_01210_));
 sky130_fd_sc_hd__and3_1 _21195_ (.A(_01160_),
    .B(_01188_),
    .C(_01194_),
    .X(_01211_));
 sky130_fd_sc_hd__a221o_1 _21196_ (.A1(_01166_),
    .A2(_01202_),
    .B1(_01210_),
    .B2(net5881),
    .C1(_01211_),
    .X(_01212_));
 sky130_fd_sc_hd__o221a_1 _21197_ (.A1(_01166_),
    .A2(_01202_),
    .B1(_01206_),
    .B2(_01207_),
    .C1(_01212_),
    .X(_01213_));
 sky130_fd_sc_hd__a22o_1 _21198_ (.A1(_01144_),
    .A2(_01147_),
    .B1(_01206_),
    .B2(_01207_),
    .X(_01214_));
 sky130_fd_sc_hd__o22a_1 _21199_ (.A1(_01144_),
    .A2(_01147_),
    .B1(_01213_),
    .B2(_01214_),
    .X(_01215_));
 sky130_fd_sc_hd__o21bai_1 _21200_ (.A1(_01115_),
    .A2(_01116_),
    .B1_N(net807),
    .Y(_01216_));
 sky130_fd_sc_hd__xnor2_1 _21201_ (.A(_01065_),
    .B(_01074_),
    .Y(_01217_));
 sky130_fd_sc_hd__xnor2_1 _21202_ (.A(_01029_),
    .B(_01217_),
    .Y(_01218_));
 sky130_fd_sc_hd__a21oi_1 _21203_ (.A1(_01114_),
    .A2(_01116_),
    .B1(_01218_),
    .Y(_01219_));
 sky130_fd_sc_hd__and2_1 _21204_ (.A(net808),
    .B(_01078_),
    .X(_01220_));
 sky130_fd_sc_hd__a21o_1 _21205_ (.A1(net761),
    .A2(net760),
    .B1(_01220_),
    .X(_01221_));
 sky130_fd_sc_hd__o21a_1 _21206_ (.A1(net808),
    .A2(_01078_),
    .B1(_01221_),
    .X(_01222_));
 sky130_fd_sc_hd__inv_2 _21207_ (.A(net1732),
    .Y(_01223_));
 sky130_fd_sc_hd__a21bo_1 _21208_ (.A1(_01223_),
    .A2(net1734),
    .B1_N(net1183),
    .X(_01224_));
 sky130_fd_sc_hd__nor2_1 _21209_ (.A(_01223_),
    .B(net1734),
    .Y(_01225_));
 sky130_fd_sc_hd__o2bb2a_1 _21210_ (.A1_N(_01007_),
    .A2_N(_01224_),
    .B1(_01225_),
    .B2(_01008_),
    .X(_01226_));
 sky130_fd_sc_hd__a21o_1 _21211_ (.A1(net1183),
    .A2(_01225_),
    .B1(_01007_),
    .X(_01227_));
 sky130_fd_sc_hd__a21bo_1 _21212_ (.A1(_01009_),
    .A2(_01227_),
    .B1_N(_01022_),
    .X(_01228_));
 sky130_fd_sc_hd__a21o_1 _21213_ (.A1(net1732),
    .A2(_01010_),
    .B1(net1183),
    .X(_01229_));
 sky130_fd_sc_hd__o211a_1 _21214_ (.A1(_01022_),
    .A2(_01226_),
    .B1(_01228_),
    .C1(_01229_),
    .X(_01230_));
 sky130_fd_sc_hd__o21a_1 _21215_ (.A1(_01027_),
    .A2(_01222_),
    .B1(net861),
    .X(_01231_));
 sky130_fd_sc_hd__a21oi_1 _21216_ (.A1(_01027_),
    .A2(_01222_),
    .B1(_01231_),
    .Y(_01232_));
 sky130_fd_sc_hd__xnor2_1 _21217_ (.A(_00938_),
    .B(_00968_),
    .Y(_01233_));
 sky130_fd_sc_hd__xnor2_1 _21218_ (.A(net861),
    .B(_01233_),
    .Y(_01234_));
 sky130_fd_sc_hd__o22a_1 _21219_ (.A1(net808),
    .A2(_01078_),
    .B1(_01027_),
    .B2(_01234_),
    .X(_01235_));
 sky130_fd_sc_hd__nor2_1 _21220_ (.A(_00938_),
    .B(_00968_),
    .Y(_01236_));
 sky130_fd_sc_hd__nand2_1 _21221_ (.A(_00938_),
    .B(_00968_),
    .Y(_01237_));
 sky130_fd_sc_hd__o21a_1 _21222_ (.A1(net861),
    .A2(_01236_),
    .B1(_01237_),
    .X(_01238_));
 sky130_fd_sc_hd__and2_1 _21223_ (.A(_01027_),
    .B(_01234_),
    .X(_01239_));
 sky130_fd_sc_hd__a211o_1 _21224_ (.A1(_01221_),
    .A2(_01235_),
    .B1(_01238_),
    .C1(_01239_),
    .X(_01240_));
 sky130_fd_sc_hd__o31a_1 _21225_ (.A1(_00938_),
    .A2(_00968_),
    .A3(_01232_),
    .B1(_01240_),
    .X(_01241_));
 sky130_fd_sc_hd__xor2_1 _21226_ (.A(_00935_),
    .B(_01241_),
    .X(_01242_));
 sky130_fd_sc_hd__xor2_1 _21227_ (.A(net5987),
    .B(net4392),
    .X(_01243_));
 sky130_fd_sc_hd__xnor2_1 _21228_ (.A(\pid_d.prev_error[0] ),
    .B(net5973),
    .Y(_01244_));
 sky130_fd_sc_hd__nor2_1 _21229_ (.A(net4298),
    .B(_01244_),
    .Y(_01245_));
 sky130_fd_sc_hd__a221o_1 _21230_ (.A1(net4320),
    .A2(net480),
    .B1(_01243_),
    .B2(net4384),
    .C1(_01245_),
    .X(_01246_));
 sky130_fd_sc_hd__a22o_1 _21231_ (.A1(net5987),
    .A2(net3122),
    .B1(net2077),
    .B2(_01246_),
    .X(_00519_));
 sky130_fd_sc_hd__nand2_1 _21232_ (.A(net5987),
    .B(net4392),
    .Y(_01247_));
 sky130_fd_sc_hd__xor2_1 _21233_ (.A(net5985),
    .B(\pid_d.prev_int[1] ),
    .X(_01248_));
 sky130_fd_sc_hd__xnor2_1 _21234_ (.A(_01247_),
    .B(_01248_),
    .Y(_01249_));
 sky130_fd_sc_hd__and2_1 _21235_ (.A(_00935_),
    .B(_01238_),
    .X(_01250_));
 sky130_fd_sc_hd__a211o_1 _21236_ (.A1(net761),
    .A2(net760),
    .B1(_01220_),
    .C1(_01239_),
    .X(_01251_));
 sky130_fd_sc_hd__o22a_1 _21237_ (.A1(_00935_),
    .A2(_01238_),
    .B1(_01239_),
    .B2(_01235_),
    .X(_01252_));
 sky130_fd_sc_hd__and2_1 _21238_ (.A(net705),
    .B(net703),
    .X(_01253_));
 sky130_fd_sc_hd__nor2_1 _21239_ (.A(net759),
    .B(_01253_),
    .Y(_01254_));
 sky130_fd_sc_hd__o21ba_1 _21240_ (.A1(_00838_),
    .A2(net1393),
    .B1_N(net1735),
    .X(_01255_));
 sky130_fd_sc_hd__a21o_1 _21241_ (.A1(_00838_),
    .A2(net1393),
    .B1(_01255_),
    .X(_01256_));
 sky130_fd_sc_hd__nand2_2 _21242_ (.A(net5861),
    .B(net5475),
    .Y(_01257_));
 sky130_fd_sc_hd__nand2_1 _21243_ (.A(net5844),
    .B(net5495),
    .Y(_01258_));
 sky130_fd_sc_hd__nand2_1 _21244_ (.A(net5811),
    .B(net5510),
    .Y(_01259_));
 sky130_fd_sc_hd__xnor2_1 _21245_ (.A(_01258_),
    .B(_01259_),
    .Y(_01260_));
 sky130_fd_sc_hd__xnor2_2 _21246_ (.A(_01257_),
    .B(_01260_),
    .Y(_01261_));
 sky130_fd_sc_hd__o21ai_1 _21247_ (.A1(_00826_),
    .A2(_00827_),
    .B1(_00828_),
    .Y(_01262_));
 sky130_fd_sc_hd__a21bo_1 _21248_ (.A1(_00826_),
    .A2(_00827_),
    .B1_N(_01262_),
    .X(_01263_));
 sky130_fd_sc_hd__and2_1 _21249_ (.A(net5962),
    .B(net5399),
    .X(_01264_));
 sky130_fd_sc_hd__nand2_1 _21250_ (.A(net5426),
    .B(net5922),
    .Y(_01265_));
 sky130_fd_sc_hd__nand2_1 _21251_ (.A(net5415),
    .B(net5945),
    .Y(_01266_));
 sky130_fd_sc_hd__xor2_1 _21252_ (.A(_01265_),
    .B(_01266_),
    .X(_01267_));
 sky130_fd_sc_hd__xnor2_2 _21253_ (.A(_01264_),
    .B(_01267_),
    .Y(_01268_));
 sky130_fd_sc_hd__xnor2_1 _21254_ (.A(_01263_),
    .B(_01268_),
    .Y(_01269_));
 sky130_fd_sc_hd__xnor2_2 _21255_ (.A(_01261_),
    .B(_01269_),
    .Y(_01270_));
 sky130_fd_sc_hd__o21a_1 _21256_ (.A1(_00844_),
    .A2(_00848_),
    .B1(net2483),
    .X(_01271_));
 sky130_fd_sc_hd__a21o_1 _21257_ (.A1(_00844_),
    .A2(_00848_),
    .B1(_01271_),
    .X(_01272_));
 sky130_fd_sc_hd__o21a_1 _21258_ (.A1(_00825_),
    .A2(_00830_),
    .B1(_00823_),
    .X(_01273_));
 sky130_fd_sc_hd__a21o_1 _21259_ (.A1(_00825_),
    .A2(_00830_),
    .B1(_01273_),
    .X(_01274_));
 sky130_fd_sc_hd__xnor2_1 _21260_ (.A(net1730),
    .B(_01274_),
    .Y(_01275_));
 sky130_fd_sc_hd__xnor2_2 _21261_ (.A(_01270_),
    .B(_01275_),
    .Y(_01276_));
 sky130_fd_sc_hd__nor2_1 _21262_ (.A(_00850_),
    .B(_00857_),
    .Y(_01277_));
 sky130_fd_sc_hd__nand2_1 _21263_ (.A(net5803),
    .B(net5535),
    .Y(_01278_));
 sky130_fd_sc_hd__nand2_1 _21264_ (.A(net5778),
    .B(net5543),
    .Y(_01279_));
 sky130_fd_sc_hd__nand2_1 _21265_ (.A(net5761),
    .B(net5570),
    .Y(_01280_));
 sky130_fd_sc_hd__xnor2_1 _21266_ (.A(_01279_),
    .B(_01280_),
    .Y(_01281_));
 sky130_fd_sc_hd__xnor2_1 _21267_ (.A(_01278_),
    .B(_01281_),
    .Y(_01282_));
 sky130_fd_sc_hd__o21a_1 _21268_ (.A1(_00852_),
    .A2(_00853_),
    .B1(_00854_),
    .X(_01283_));
 sky130_fd_sc_hd__a21oi_2 _21269_ (.A1(_00852_),
    .A2(_00853_),
    .B1(_01283_),
    .Y(_01284_));
 sky130_fd_sc_hd__o21a_1 _21270_ (.A1(_00840_),
    .A2(_00841_),
    .B1(_00842_),
    .X(_01285_));
 sky130_fd_sc_hd__a21oi_2 _21271_ (.A1(_00840_),
    .A2(_00841_),
    .B1(_01285_),
    .Y(_01286_));
 sky130_fd_sc_hd__xor2_1 _21272_ (.A(_01284_),
    .B(_01286_),
    .X(_01287_));
 sky130_fd_sc_hd__xnor2_1 _21273_ (.A(_01282_),
    .B(_01287_),
    .Y(_01288_));
 sky130_fd_sc_hd__nor2_1 _21274_ (.A(net3842),
    .B(_00856_),
    .Y(_01289_));
 sky130_fd_sc_hd__nand2_1 _21275_ (.A(net5637),
    .B(net5674),
    .Y(_01290_));
 sky130_fd_sc_hd__nand2_1 _21276_ (.A(net5687),
    .B(net5626),
    .Y(_01291_));
 sky130_fd_sc_hd__xor2_1 _21277_ (.A(_01290_),
    .B(_01291_),
    .X(_01292_));
 sky130_fd_sc_hd__nand2_1 _21278_ (.A(net5741),
    .B(net5590),
    .Y(_01293_));
 sky130_fd_sc_hd__nand2_1 _21279_ (.A(net5731),
    .B(net5598),
    .Y(_01294_));
 sky130_fd_sc_hd__nand2_1 _21280_ (.A(net5702),
    .B(net5615),
    .Y(_01295_));
 sky130_fd_sc_hd__xor2_1 _21281_ (.A(_01294_),
    .B(_01295_),
    .X(_01296_));
 sky130_fd_sc_hd__xnor2_1 _21282_ (.A(_01293_),
    .B(_01296_),
    .Y(_01297_));
 sky130_fd_sc_hd__xor2_1 _21283_ (.A(_01292_),
    .B(_01297_),
    .X(_01298_));
 sky130_fd_sc_hd__xor2_1 _21284_ (.A(_01289_),
    .B(_01298_),
    .X(_01299_));
 sky130_fd_sc_hd__xnor2_1 _21285_ (.A(_01288_),
    .B(_01299_),
    .Y(_01300_));
 sky130_fd_sc_hd__xor2_1 _21286_ (.A(net1391),
    .B(net1390),
    .X(_01301_));
 sky130_fd_sc_hd__xnor2_1 _21287_ (.A(_01276_),
    .B(_01301_),
    .Y(_01302_));
 sky130_fd_sc_hd__a21bo_1 _21288_ (.A1(net1737),
    .A2(net1736),
    .B1_N(_00834_),
    .X(_01303_));
 sky130_fd_sc_hd__o21a_2 _21289_ (.A1(net1737),
    .A2(net1736),
    .B1(_01303_),
    .X(_01304_));
 sky130_fd_sc_hd__o21a_1 _21290_ (.A1(_00819_),
    .A2(_00820_),
    .B1(_00821_),
    .X(_01305_));
 sky130_fd_sc_hd__a21oi_2 _21291_ (.A1(_00819_),
    .A2(_00820_),
    .B1(_01305_),
    .Y(_01306_));
 sky130_fd_sc_hd__a21o_1 _21292_ (.A1(net3811),
    .A2(_12515_),
    .B1(_12516_),
    .X(_01307_));
 sky130_fd_sc_hd__o21ai_1 _21293_ (.A1(net3811),
    .A2(_12515_),
    .B1(_01307_),
    .Y(_01308_));
 sky130_fd_sc_hd__nand2_1 _21294_ (.A(net5473),
    .B(_01308_),
    .Y(_01309_));
 sky130_fd_sc_hd__xnor2_1 _21295_ (.A(net5455),
    .B(_01309_),
    .Y(_01310_));
 sky130_fd_sc_hd__nand2_1 _21296_ (.A(net5889),
    .B(_01310_),
    .Y(_01311_));
 sky130_fd_sc_hd__xor2_1 _21297_ (.A(_01306_),
    .B(_01311_),
    .X(_01312_));
 sky130_fd_sc_hd__xnor2_2 _21298_ (.A(_01304_),
    .B(_01312_),
    .Y(_01313_));
 sky130_fd_sc_hd__xor2_1 _21299_ (.A(net1050),
    .B(_01313_),
    .X(_01314_));
 sky130_fd_sc_hd__xnor2_1 _21300_ (.A(_01256_),
    .B(_01314_),
    .Y(_01315_));
 sky130_fd_sc_hd__o31a_1 _21301_ (.A1(net5473),
    .A2(_12515_),
    .A3(_12516_),
    .B1(_00862_),
    .X(_01316_));
 sky130_fd_sc_hd__inv_2 _21302_ (.A(net5487),
    .Y(_01317_));
 sky130_fd_sc_hd__a211o_1 _21303_ (.A1(_00862_),
    .A2(_00868_),
    .B1(_00864_),
    .C1(net3796),
    .X(_01318_));
 sky130_fd_sc_hd__o21a_1 _21304_ (.A1(_00868_),
    .A2(_01316_),
    .B1(_01318_),
    .X(_01319_));
 sky130_fd_sc_hd__o21ai_1 _21305_ (.A1(net3796),
    .A2(net3119),
    .B1(_00864_),
    .Y(_01320_));
 sky130_fd_sc_hd__o22a_1 _21306_ (.A1(net3119),
    .A2(_01319_),
    .B1(_01320_),
    .B2(_00862_),
    .X(_01321_));
 sky130_fd_sc_hd__a21bo_1 _21307_ (.A1(_00860_),
    .A2(_00875_),
    .B1_N(net1052),
    .X(_01322_));
 sky130_fd_sc_hd__o21a_1 _21308_ (.A1(_00860_),
    .A2(_00875_),
    .B1(_01322_),
    .X(_01323_));
 sky130_fd_sc_hd__xor2_1 _21309_ (.A(_01321_),
    .B(_01323_),
    .X(_01324_));
 sky130_fd_sc_hd__xnor2_1 _21310_ (.A(_01315_),
    .B(_01324_),
    .Y(_01325_));
 sky130_fd_sc_hd__a21bo_1 _21311_ (.A1(_00877_),
    .A2(_00933_),
    .B1_N(_00931_),
    .X(_01326_));
 sky130_fd_sc_hd__o21ai_1 _21312_ (.A1(_00877_),
    .A2(_00933_),
    .B1(_01326_),
    .Y(_01327_));
 sky130_fd_sc_hd__nor2_1 _21313_ (.A(_01325_),
    .B(net758),
    .Y(_01328_));
 sky130_fd_sc_hd__nand2_1 _21314_ (.A(_01325_),
    .B(net758),
    .Y(_01329_));
 sky130_fd_sc_hd__and2b_1 _21315_ (.A_N(_01328_),
    .B(_01329_),
    .X(_01330_));
 sky130_fd_sc_hd__xnor2_1 _21316_ (.A(_01254_),
    .B(_01330_),
    .Y(_01331_));
 sky130_fd_sc_hd__xnor2_1 _21317_ (.A(\pid_d.prev_error[1] ),
    .B(net5972),
    .Y(_01332_));
 sky130_fd_sc_hd__and3_1 _21318_ (.A(\pid_d.prev_error[0] ),
    .B(net5973),
    .C(_01332_),
    .X(_01333_));
 sky130_fd_sc_hd__a21oi_1 _21319_ (.A1(\pid_d.prev_error[0] ),
    .A2(net5973),
    .B1(_01332_),
    .Y(_01334_));
 sky130_fd_sc_hd__o21a_1 _21320_ (.A1(_01333_),
    .A2(_01334_),
    .B1(net4356),
    .X(_01335_));
 sky130_fd_sc_hd__a221o_1 _21321_ (.A1(net4384),
    .A2(_01249_),
    .B1(net561),
    .B2(net4320),
    .C1(_01335_),
    .X(_01336_));
 sky130_fd_sc_hd__a22o_1 _21322_ (.A1(net9009),
    .A2(net3122),
    .B1(net2077),
    .B2(_01336_),
    .X(_00520_));
 sky130_fd_sc_hd__or2_1 _21323_ (.A(net5984),
    .B(\pid_d.prev_int[1] ),
    .X(_01337_));
 sky130_fd_sc_hd__a22o_1 _21324_ (.A1(\pid_d.curr_int[0] ),
    .A2(\pid_d.prev_int[0] ),
    .B1(\pid_d.prev_int[1] ),
    .B2(net5984),
    .X(_01338_));
 sky130_fd_sc_hd__nand2_1 _21325_ (.A(_01337_),
    .B(_01338_),
    .Y(_01339_));
 sky130_fd_sc_hd__xnor2_1 _21326_ (.A(net5983),
    .B(\pid_d.prev_int[2] ),
    .Y(_01340_));
 sky130_fd_sc_hd__xnor2_1 _21327_ (.A(_01339_),
    .B(_01340_),
    .Y(_01341_));
 sky130_fd_sc_hd__o31ai_2 _21328_ (.A1(net759),
    .A2(_01253_),
    .A3(_01328_),
    .B1(_01329_),
    .Y(_01342_));
 sky130_fd_sc_hd__nand2_1 _21329_ (.A(net5739),
    .B(net5560),
    .Y(_01343_));
 sky130_fd_sc_hd__nand2_1 _21330_ (.A(net5705),
    .B(net5598),
    .Y(_01344_));
 sky130_fd_sc_hd__nand2_1 _21331_ (.A(net5731),
    .B(net5576),
    .Y(_01345_));
 sky130_fd_sc_hd__xnor2_1 _21332_ (.A(_01344_),
    .B(_01345_),
    .Y(_01346_));
 sky130_fd_sc_hd__xnor2_1 _21333_ (.A(_01343_),
    .B(_01346_),
    .Y(_01347_));
 sky130_fd_sc_hd__and2_1 _21334_ (.A(net5687),
    .B(net5616),
    .X(_01348_));
 sky130_fd_sc_hd__nand2_4 _21335_ (.A(net5626),
    .B(net5674),
    .Y(_01349_));
 sky130_fd_sc_hd__xor2_1 _21336_ (.A(net5654),
    .B(_01349_),
    .X(_01350_));
 sky130_fd_sc_hd__nand2_1 _21337_ (.A(_01348_),
    .B(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hd__nor2_1 _21338_ (.A(net5687),
    .B(_01349_),
    .Y(_01352_));
 sky130_fd_sc_hd__o21ai_1 _21339_ (.A1(_01348_),
    .A2(_01352_),
    .B1(net5638),
    .Y(_01353_));
 sky130_fd_sc_hd__or2b_1 _21340_ (.A(net5638),
    .B_N(net5654),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _21341_ (.A0(net5654),
    .A1(_01354_),
    .S(_01349_),
    .X(_01355_));
 sky130_fd_sc_hd__o32a_1 _21342_ (.A1(net5638),
    .A2(net5616),
    .A3(_01350_),
    .B1(_01355_),
    .B2(net5687),
    .X(_01356_));
 sky130_fd_sc_hd__and3_1 _21343_ (.A(_01351_),
    .B(_01353_),
    .C(_01356_),
    .X(_01357_));
 sky130_fd_sc_hd__xnor2_1 _21344_ (.A(_01347_),
    .B(_01357_),
    .Y(_01358_));
 sky130_fd_sc_hd__nand2_1 _21345_ (.A(_01292_),
    .B(_01297_),
    .Y(_01359_));
 sky130_fd_sc_hd__nand2_2 _21346_ (.A(net5807),
    .B(net5511),
    .Y(_01360_));
 sky130_fd_sc_hd__nand2_1 _21347_ (.A(net5758),
    .B(net5543),
    .Y(_01361_));
 sky130_fd_sc_hd__nand2_1 _21348_ (.A(net5777),
    .B(net5535),
    .Y(_01362_));
 sky130_fd_sc_hd__xnor2_1 _21349_ (.A(_01361_),
    .B(_01362_),
    .Y(_01363_));
 sky130_fd_sc_hd__xnor2_2 _21350_ (.A(_01360_),
    .B(_01363_),
    .Y(_01364_));
 sky130_fd_sc_hd__o21a_1 _21351_ (.A1(_01293_),
    .A2(_01294_),
    .B1(_01295_),
    .X(_01365_));
 sky130_fd_sc_hd__a21oi_2 _21352_ (.A1(_01293_),
    .A2(_01294_),
    .B1(_01365_),
    .Y(_01366_));
 sky130_fd_sc_hd__o21a_1 _21353_ (.A1(_01278_),
    .A2(_01279_),
    .B1(_01280_),
    .X(_01367_));
 sky130_fd_sc_hd__a21oi_2 _21354_ (.A1(_01278_),
    .A2(_01279_),
    .B1(_01367_),
    .Y(_01368_));
 sky130_fd_sc_hd__xnor2_1 _21355_ (.A(_01366_),
    .B(_01368_),
    .Y(_01369_));
 sky130_fd_sc_hd__xnor2_2 _21356_ (.A(_01364_),
    .B(_01369_),
    .Y(_01370_));
 sky130_fd_sc_hd__xor2_1 _21357_ (.A(_01359_),
    .B(_01370_),
    .X(_01371_));
 sky130_fd_sc_hd__xnor2_1 _21358_ (.A(net1729),
    .B(_01371_),
    .Y(_01372_));
 sky130_fd_sc_hd__nand2_1 _21359_ (.A(net5844),
    .B(net5476),
    .Y(_01373_));
 sky130_fd_sc_hd__nand2_1 _21360_ (.A(net5811),
    .B(net5495),
    .Y(_01374_));
 sky130_fd_sc_hd__nand2_1 _21361_ (.A(net5865),
    .B(net5457),
    .Y(_01375_));
 sky130_fd_sc_hd__xnor2_1 _21362_ (.A(_01374_),
    .B(_01375_),
    .Y(_01376_));
 sky130_fd_sc_hd__xnor2_1 _21363_ (.A(_01373_),
    .B(_01376_),
    .Y(_01377_));
 sky130_fd_sc_hd__o21ai_1 _21364_ (.A1(_01257_),
    .A2(_01258_),
    .B1(_01259_),
    .Y(_01378_));
 sky130_fd_sc_hd__a21bo_1 _21365_ (.A1(_01257_),
    .A2(_01258_),
    .B1_N(_01378_),
    .X(_01379_));
 sky130_fd_sc_hd__and2_1 _21366_ (.A(net5963),
    .B(net5382),
    .X(_01380_));
 sky130_fd_sc_hd__nand2_1 _21367_ (.A(net5416),
    .B(net5922),
    .Y(_01381_));
 sky130_fd_sc_hd__nand2_1 _21368_ (.A(net5944),
    .B(net5399),
    .Y(_01382_));
 sky130_fd_sc_hd__xor2_1 _21369_ (.A(_01381_),
    .B(_01382_),
    .X(_01383_));
 sky130_fd_sc_hd__xnor2_1 _21370_ (.A(_01380_),
    .B(_01383_),
    .Y(_01384_));
 sky130_fd_sc_hd__xnor2_1 _21371_ (.A(_01379_),
    .B(_01384_),
    .Y(_01385_));
 sky130_fd_sc_hd__xnor2_1 _21372_ (.A(_01377_),
    .B(_01385_),
    .Y(_01386_));
 sky130_fd_sc_hd__a21bo_1 _21373_ (.A1(_01284_),
    .A2(_01286_),
    .B1_N(_01282_),
    .X(_01387_));
 sky130_fd_sc_hd__o21ai_1 _21374_ (.A1(_01284_),
    .A2(_01286_),
    .B1(_01387_),
    .Y(_01388_));
 sky130_fd_sc_hd__o21a_1 _21375_ (.A1(_01263_),
    .A2(_01268_),
    .B1(_01261_),
    .X(_01389_));
 sky130_fd_sc_hd__a21o_1 _21376_ (.A1(_01263_),
    .A2(_01268_),
    .B1(_01389_),
    .X(_01390_));
 sky130_fd_sc_hd__xnor2_1 _21377_ (.A(net1728),
    .B(_01390_),
    .Y(_01391_));
 sky130_fd_sc_hd__xnor2_1 _21378_ (.A(_01386_),
    .B(_01391_),
    .Y(_01392_));
 sky130_fd_sc_hd__a21o_1 _21379_ (.A1(_01288_),
    .A2(_01289_),
    .B1(_01298_),
    .X(_01393_));
 sky130_fd_sc_hd__o21a_1 _21380_ (.A1(_01288_),
    .A2(_01289_),
    .B1(_01393_),
    .X(_01394_));
 sky130_fd_sc_hd__xor2_1 _21381_ (.A(_01392_),
    .B(net1181),
    .X(_01395_));
 sky130_fd_sc_hd__xnor2_2 _21382_ (.A(net1182),
    .B(_01395_),
    .Y(_01396_));
 sky130_fd_sc_hd__o21ba_1 _21383_ (.A1(_01276_),
    .A2(net1390),
    .B1_N(net1391),
    .X(_01397_));
 sky130_fd_sc_hd__a21o_1 _21384_ (.A1(_01276_),
    .A2(net1390),
    .B1(_01397_),
    .X(_01398_));
 sky130_fd_sc_hd__a21o_1 _21385_ (.A1(_01270_),
    .A2(_01274_),
    .B1(net1730),
    .X(_01399_));
 sky130_fd_sc_hd__o21ai_1 _21386_ (.A1(_01270_),
    .A2(_01274_),
    .B1(_01399_),
    .Y(_01400_));
 sky130_fd_sc_hd__o21ba_1 _21387_ (.A1(_01265_),
    .A2(_01266_),
    .B1_N(_01264_),
    .X(_01401_));
 sky130_fd_sc_hd__a21oi_2 _21388_ (.A1(_01265_),
    .A2(_01266_),
    .B1(_01401_),
    .Y(_01402_));
 sky130_fd_sc_hd__xnor2_2 _21389_ (.A(net5651),
    .B(_01402_),
    .Y(_01403_));
 sky130_fd_sc_hd__a21bo_1 _21390_ (.A1(net5456),
    .A2(net2479),
    .B1_N(net5426),
    .X(_01404_));
 sky130_fd_sc_hd__inv_2 _21391_ (.A(net5462),
    .Y(_01405_));
 sky130_fd_sc_hd__or4_1 _21392_ (.A(net5444),
    .B(net3812),
    .C(net3789),
    .D(_00821_),
    .X(_01406_));
 sky130_fd_sc_hd__a21o_1 _21393_ (.A1(_01404_),
    .A2(_01406_),
    .B1(net3117),
    .X(_01407_));
 sky130_fd_sc_hd__xnor2_1 _21394_ (.A(_01403_),
    .B(_01407_),
    .Y(_01408_));
 sky130_fd_sc_hd__xnor2_1 _21395_ (.A(_01400_),
    .B(_01408_),
    .Y(_01409_));
 sky130_fd_sc_hd__xnor2_1 _21396_ (.A(_01398_),
    .B(_01409_),
    .Y(_01410_));
 sky130_fd_sc_hd__xnor2_1 _21397_ (.A(_01396_),
    .B(_01410_),
    .Y(_01411_));
 sky130_fd_sc_hd__o31a_1 _21398_ (.A1(net5455),
    .A2(_00820_),
    .A3(_00821_),
    .B1(_01304_),
    .X(_01412_));
 sky130_fd_sc_hd__a211o_1 _21399_ (.A1(_01304_),
    .A2(_01309_),
    .B1(_01306_),
    .C1(net3789),
    .X(_01413_));
 sky130_fd_sc_hd__o21a_1 _21400_ (.A1(_01309_),
    .A2(_01412_),
    .B1(_01413_),
    .X(_01414_));
 sky130_fd_sc_hd__o21ai_1 _21401_ (.A1(net3789),
    .A2(net3118),
    .B1(_01306_),
    .Y(_01415_));
 sky130_fd_sc_hd__o22a_1 _21402_ (.A1(net3118),
    .A2(_01414_),
    .B1(_01415_),
    .B2(_01304_),
    .X(_01416_));
 sky130_fd_sc_hd__a221o_1 _21403_ (.A1(_00838_),
    .A2(net1393),
    .B1(net1050),
    .B2(_01313_),
    .C1(_01255_),
    .X(_01417_));
 sky130_fd_sc_hd__o21a_2 _21404_ (.A1(net1050),
    .A2(_01313_),
    .B1(_01417_),
    .X(_01418_));
 sky130_fd_sc_hd__xnor2_1 _21405_ (.A(net860),
    .B(_01418_),
    .Y(_01419_));
 sky130_fd_sc_hd__xnor2_1 _21406_ (.A(net806),
    .B(_01419_),
    .Y(_01420_));
 sky130_fd_sc_hd__a21bo_1 _21407_ (.A1(_01321_),
    .A2(_01323_),
    .B1_N(_01315_),
    .X(_01421_));
 sky130_fd_sc_hd__o21a_1 _21408_ (.A1(_01321_),
    .A2(_01323_),
    .B1(_01421_),
    .X(_01422_));
 sky130_fd_sc_hd__nand2_1 _21409_ (.A(_01420_),
    .B(net757),
    .Y(_01423_));
 sky130_fd_sc_hd__or2_1 _21410_ (.A(_01420_),
    .B(net757),
    .X(_01424_));
 sky130_fd_sc_hd__nand2_1 _21411_ (.A(_01423_),
    .B(_01424_),
    .Y(_01425_));
 sky130_fd_sc_hd__xor2_1 _21412_ (.A(_01342_),
    .B(_01425_),
    .X(_01426_));
 sky130_fd_sc_hd__nand2_1 _21413_ (.A(net4320),
    .B(net555),
    .Y(_01427_));
 sky130_fd_sc_hd__or2_1 _21414_ (.A(\pid_d.prev_error[1] ),
    .B(net5972),
    .X(_01428_));
 sky130_fd_sc_hd__a22o_1 _21415_ (.A1(\pid_d.prev_error[0] ),
    .A2(net5973),
    .B1(\pid_d.prev_error[1] ),
    .B2(net5972),
    .X(_01429_));
 sky130_fd_sc_hd__and2_1 _21416_ (.A(_01428_),
    .B(_01429_),
    .X(_01430_));
 sky130_fd_sc_hd__xor2_1 _21417_ (.A(\pid_d.prev_error[2] ),
    .B(net5971),
    .X(_01431_));
 sky130_fd_sc_hd__nor2_1 _21418_ (.A(_01430_),
    .B(_01431_),
    .Y(_01432_));
 sky130_fd_sc_hd__and3_1 _21419_ (.A(_01428_),
    .B(_01429_),
    .C(_01431_),
    .X(_01433_));
 sky130_fd_sc_hd__or3_1 _21420_ (.A(net4298),
    .B(_01432_),
    .C(_01433_),
    .X(_01434_));
 sky130_fd_sc_hd__o211ai_1 _21421_ (.A1(_04875_),
    .A2(net2478),
    .B1(_01427_),
    .C1(_01434_),
    .Y(_01435_));
 sky130_fd_sc_hd__a22o_1 _21422_ (.A1(net9079),
    .A2(net3122),
    .B1(net2077),
    .B2(_01435_),
    .X(_00521_));
 sky130_fd_sc_hd__a21o_1 _21423_ (.A1(_01337_),
    .A2(_01338_),
    .B1(\pid_d.prev_int[2] ),
    .X(_01436_));
 sky130_fd_sc_hd__a31o_1 _21424_ (.A1(\pid_d.prev_int[2] ),
    .A2(_01337_),
    .A3(_01338_),
    .B1(net5983),
    .X(_01437_));
 sky130_fd_sc_hd__and2_1 _21425_ (.A(_01436_),
    .B(_01437_),
    .X(_01438_));
 sky130_fd_sc_hd__xnor2_1 _21426_ (.A(\pid_d.curr_int[3] ),
    .B(\pid_d.prev_int[3] ),
    .Y(_01439_));
 sky130_fd_sc_hd__xnor2_1 _21427_ (.A(_01438_),
    .B(_01439_),
    .Y(_01440_));
 sky130_fd_sc_hd__o21ba_1 _21428_ (.A1(_01396_),
    .A2(_01409_),
    .B1_N(_01398_),
    .X(_01441_));
 sky130_fd_sc_hd__a21o_1 _21429_ (.A1(_01396_),
    .A2(_01409_),
    .B1(_01441_),
    .X(_01442_));
 sky130_fd_sc_hd__nand2_1 _21430_ (.A(net5426),
    .B(net5894),
    .Y(_01443_));
 sky130_fd_sc_hd__xor2_1 _21431_ (.A(_01403_),
    .B(_01443_),
    .X(_01444_));
 sky130_fd_sc_hd__and3_1 _21432_ (.A(net5456),
    .B(net5890),
    .C(net2479),
    .X(_01445_));
 sky130_fd_sc_hd__a21o_1 _21433_ (.A1(_01444_),
    .A2(_01445_),
    .B1(_01400_),
    .X(_01446_));
 sky130_fd_sc_hd__o21a_1 _21434_ (.A1(_01444_),
    .A2(_01445_),
    .B1(_01446_),
    .X(_01447_));
 sky130_fd_sc_hd__nand2_1 _21435_ (.A(net3807),
    .B(net5654),
    .Y(_01448_));
 sky130_fd_sc_hd__nand2_1 _21436_ (.A(net5685),
    .B(net5608),
    .Y(_01449_));
 sky130_fd_sc_hd__nand2_1 _21437_ (.A(net5618),
    .B(net5673),
    .Y(_01450_));
 sky130_fd_sc_hd__xnor2_1 _21438_ (.A(_01449_),
    .B(_01450_),
    .Y(_01451_));
 sky130_fd_sc_hd__xnor2_1 _21439_ (.A(_01448_),
    .B(_01451_),
    .Y(_01452_));
 sky130_fd_sc_hd__a21bo_1 _21440_ (.A1(_01349_),
    .A2(_01354_),
    .B1_N(_01348_),
    .X(_01453_));
 sky130_fd_sc_hd__o21ai_2 _21441_ (.A1(_01349_),
    .A2(_01354_),
    .B1(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__nand2_2 _21442_ (.A(net5739),
    .B(net5542),
    .Y(_01455_));
 sky130_fd_sc_hd__nand2_1 _21443_ (.A(net5705),
    .B(net5582),
    .Y(_01456_));
 sky130_fd_sc_hd__nand2_1 _21444_ (.A(net5724),
    .B(net5565),
    .Y(_01457_));
 sky130_fd_sc_hd__xor2_1 _21445_ (.A(_01456_),
    .B(_01457_),
    .X(_01458_));
 sky130_fd_sc_hd__xnor2_2 _21446_ (.A(_01455_),
    .B(_01458_),
    .Y(_01459_));
 sky130_fd_sc_hd__xor2_1 _21447_ (.A(_01454_),
    .B(_01459_),
    .X(_01460_));
 sky130_fd_sc_hd__xnor2_1 _21448_ (.A(_01452_),
    .B(_01460_),
    .Y(_01461_));
 sky130_fd_sc_hd__inv_2 _21449_ (.A(_01349_),
    .Y(_01462_));
 sky130_fd_sc_hd__o21ai_1 _21450_ (.A1(_01348_),
    .A2(_01462_),
    .B1(net5638),
    .Y(_01463_));
 sky130_fd_sc_hd__o211a_1 _21451_ (.A1(_01348_),
    .A2(_01355_),
    .B1(_01463_),
    .C1(_01351_),
    .X(_01464_));
 sky130_fd_sc_hd__o32a_1 _21452_ (.A1(net5616),
    .A2(_00851_),
    .A3(_01349_),
    .B1(_01464_),
    .B2(_01347_),
    .X(_01465_));
 sky130_fd_sc_hd__nand2_1 _21453_ (.A(net5807),
    .B(net5490),
    .Y(_01466_));
 sky130_fd_sc_hd__nand2_1 _21454_ (.A(net5766),
    .B(net5529),
    .Y(_01467_));
 sky130_fd_sc_hd__nand2_1 _21455_ (.A(net5777),
    .B(net5511),
    .Y(_01468_));
 sky130_fd_sc_hd__xnor2_1 _21456_ (.A(_01467_),
    .B(_01468_),
    .Y(_01469_));
 sky130_fd_sc_hd__xnor2_1 _21457_ (.A(_01466_),
    .B(_01469_),
    .Y(_01470_));
 sky130_fd_sc_hd__o21a_1 _21458_ (.A1(_01343_),
    .A2(_01345_),
    .B1(_01344_),
    .X(_01471_));
 sky130_fd_sc_hd__a21oi_2 _21459_ (.A1(_01343_),
    .A2(_01345_),
    .B1(_01471_),
    .Y(_01472_));
 sky130_fd_sc_hd__o21a_1 _21460_ (.A1(_01360_),
    .A2(_01362_),
    .B1(_01361_),
    .X(_01473_));
 sky130_fd_sc_hd__a21oi_2 _21461_ (.A1(_01360_),
    .A2(_01362_),
    .B1(_01473_),
    .Y(_01474_));
 sky130_fd_sc_hd__xnor2_1 _21462_ (.A(_01472_),
    .B(_01474_),
    .Y(_01475_));
 sky130_fd_sc_hd__xnor2_1 _21463_ (.A(_01470_),
    .B(_01475_),
    .Y(_01476_));
 sky130_fd_sc_hd__nor2_1 _21464_ (.A(net1726),
    .B(_01476_),
    .Y(_01477_));
 sky130_fd_sc_hd__nand2_1 _21465_ (.A(net1726),
    .B(_01476_),
    .Y(_01478_));
 sky130_fd_sc_hd__and2b_1 _21466_ (.A_N(_01477_),
    .B(_01478_),
    .X(_01479_));
 sky130_fd_sc_hd__xor2_1 _21467_ (.A(net1727),
    .B(_01479_),
    .X(_01480_));
 sky130_fd_sc_hd__o21a_1 _21468_ (.A1(net1729),
    .A2(_01370_),
    .B1(_01359_),
    .X(_01481_));
 sky130_fd_sc_hd__a21o_1 _21469_ (.A1(net1729),
    .A2(_01370_),
    .B1(_01481_),
    .X(_01482_));
 sky130_fd_sc_hd__nand2_1 _21470_ (.A(net5814),
    .B(net5482),
    .Y(_01483_));
 sky130_fd_sc_hd__nand2_1 _21471_ (.A(net5864),
    .B(net5429),
    .Y(_01484_));
 sky130_fd_sc_hd__nand2_1 _21472_ (.A(net5843),
    .B(net5458),
    .Y(_01485_));
 sky130_fd_sc_hd__xor2_1 _21473_ (.A(_01484_),
    .B(_01485_),
    .X(_01486_));
 sky130_fd_sc_hd__xnor2_2 _21474_ (.A(_01483_),
    .B(_01486_),
    .Y(_01487_));
 sky130_fd_sc_hd__o21a_1 _21475_ (.A1(_01373_),
    .A2(_01375_),
    .B1(_01374_),
    .X(_01488_));
 sky130_fd_sc_hd__a21oi_2 _21476_ (.A1(_01373_),
    .A2(_01375_),
    .B1(_01488_),
    .Y(_01489_));
 sky130_fd_sc_hd__xor2_1 _21477_ (.A(net5961),
    .B(net5943),
    .X(_01490_));
 sky130_fd_sc_hd__nand2_1 _21478_ (.A(net5383),
    .B(_01490_),
    .Y(_01491_));
 sky130_fd_sc_hd__nand2_1 _21479_ (.A(net5920),
    .B(net5400),
    .Y(_01492_));
 sky130_fd_sc_hd__xor2_2 _21480_ (.A(_01491_),
    .B(_01492_),
    .X(_01493_));
 sky130_fd_sc_hd__xnor2_1 _21481_ (.A(_01489_),
    .B(_01493_),
    .Y(_01494_));
 sky130_fd_sc_hd__xnor2_2 _21482_ (.A(_01487_),
    .B(_01494_),
    .Y(_01495_));
 sky130_fd_sc_hd__a21bo_1 _21483_ (.A1(_01366_),
    .A2(_01368_),
    .B1_N(_01364_),
    .X(_01496_));
 sky130_fd_sc_hd__o21ai_1 _21484_ (.A1(_01366_),
    .A2(_01368_),
    .B1(_01496_),
    .Y(_01497_));
 sky130_fd_sc_hd__o21a_1 _21485_ (.A1(_01379_),
    .A2(_01384_),
    .B1(_01377_),
    .X(_01498_));
 sky130_fd_sc_hd__a21o_1 _21486_ (.A1(_01379_),
    .A2(_01384_),
    .B1(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__xnor2_1 _21487_ (.A(net1725),
    .B(_01499_),
    .Y(_01500_));
 sky130_fd_sc_hd__xnor2_2 _21488_ (.A(_01495_),
    .B(_01500_),
    .Y(_01501_));
 sky130_fd_sc_hd__xor2_1 _21489_ (.A(net1180),
    .B(_01501_),
    .X(_01502_));
 sky130_fd_sc_hd__xnor2_1 _21490_ (.A(net1049),
    .B(_01502_),
    .Y(_01503_));
 sky130_fd_sc_hd__o21a_1 _21491_ (.A1(net1728),
    .A2(_01390_),
    .B1(_01386_),
    .X(_01504_));
 sky130_fd_sc_hd__a21o_1 _21492_ (.A1(net1728),
    .A2(_01390_),
    .B1(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__or2_1 _21493_ (.A(net5651),
    .B(_01402_),
    .X(_01506_));
 sky130_fd_sc_hd__a21o_1 _21494_ (.A1(net5427),
    .A2(_01506_),
    .B1(net5416),
    .X(_01507_));
 sky130_fd_sc_hd__and2_1 _21495_ (.A(net5651),
    .B(_01402_),
    .X(_01508_));
 sky130_fd_sc_hd__o211ai_1 _21496_ (.A1(net5427),
    .A2(_01508_),
    .B1(_01506_),
    .C1(net5416),
    .Y(_01509_));
 sky130_fd_sc_hd__nand2_1 _21497_ (.A(net5416),
    .B(net5894),
    .Y(_01510_));
 sky130_fd_sc_hd__a32o_1 _21498_ (.A1(net5894),
    .A2(_01507_),
    .A3(_01509_),
    .B1(_01510_),
    .B2(_01508_),
    .X(_01511_));
 sky130_fd_sc_hd__o21ba_1 _21499_ (.A1(_01381_),
    .A2(_01382_),
    .B1_N(_01380_),
    .X(_01512_));
 sky130_fd_sc_hd__a21oi_1 _21500_ (.A1(_01381_),
    .A2(_01382_),
    .B1(_01512_),
    .Y(_01513_));
 sky130_fd_sc_hd__xor2_1 _21501_ (.A(_01511_),
    .B(_01513_),
    .X(_01514_));
 sky130_fd_sc_hd__xnor2_2 _21502_ (.A(net1179),
    .B(_01514_),
    .Y(_01515_));
 sky130_fd_sc_hd__o21ba_1 _21503_ (.A1(net1182),
    .A2(net1181),
    .B1_N(_01392_),
    .X(_01516_));
 sky130_fd_sc_hd__a21oi_1 _21504_ (.A1(net1182),
    .A2(net1181),
    .B1(_01516_),
    .Y(_01517_));
 sky130_fd_sc_hd__xor2_1 _21505_ (.A(_01515_),
    .B(net947),
    .X(_01518_));
 sky130_fd_sc_hd__xnor2_2 _21506_ (.A(net948),
    .B(_01518_),
    .Y(_01519_));
 sky130_fd_sc_hd__xor2_1 _21507_ (.A(_01447_),
    .B(_01519_),
    .X(_01520_));
 sky130_fd_sc_hd__xnor2_1 _21508_ (.A(_01442_),
    .B(_01520_),
    .Y(_01521_));
 sky130_fd_sc_hd__or2_1 _21509_ (.A(net806),
    .B(net757),
    .X(_01522_));
 sky130_fd_sc_hd__and2_1 _21510_ (.A(net806),
    .B(net757),
    .X(_01523_));
 sky130_fd_sc_hd__a21oi_1 _21511_ (.A1(net860),
    .A2(_01522_),
    .B1(_01523_),
    .Y(_01524_));
 sky130_fd_sc_hd__inv_2 _21512_ (.A(_01524_),
    .Y(_01525_));
 sky130_fd_sc_hd__and3_1 _21513_ (.A(net860),
    .B(net806),
    .C(net757),
    .X(_01526_));
 sky130_fd_sc_hd__a21o_1 _21514_ (.A1(_01418_),
    .A2(_01525_),
    .B1(_01526_),
    .X(_01527_));
 sky130_fd_sc_hd__nor2_1 _21515_ (.A(net860),
    .B(_01522_),
    .Y(_01528_));
 sky130_fd_sc_hd__nor2_1 _21516_ (.A(_01418_),
    .B(_01525_),
    .Y(_01529_));
 sky130_fd_sc_hd__o21ba_1 _21517_ (.A1(_01528_),
    .A2(_01529_),
    .B1_N(_01342_),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _21518_ (.A0(_01528_),
    .A1(_01526_),
    .S(_01418_),
    .X(_01531_));
 sky130_fd_sc_hd__a211o_1 _21519_ (.A1(_01342_),
    .A2(_01527_),
    .B1(_01530_),
    .C1(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__xor2_1 _21520_ (.A(_01521_),
    .B(net478),
    .X(_01533_));
 sky130_fd_sc_hd__a31o_1 _21521_ (.A1(net5971),
    .A2(_01428_),
    .A3(_01429_),
    .B1(\pid_d.prev_error[2] ),
    .X(_01534_));
 sky130_fd_sc_hd__o21ai_2 _21522_ (.A1(net5971),
    .A2(_01430_),
    .B1(_01534_),
    .Y(_01535_));
 sky130_fd_sc_hd__xnor2_1 _21523_ (.A(\pid_d.prev_error[3] ),
    .B(net5970),
    .Y(_01536_));
 sky130_fd_sc_hd__nand2_1 _21524_ (.A(_01535_),
    .B(_01536_),
    .Y(_01537_));
 sky130_fd_sc_hd__or2_1 _21525_ (.A(_01535_),
    .B(_01536_),
    .X(_01538_));
 sky130_fd_sc_hd__and3_1 _21526_ (.A(net4357),
    .B(_01537_),
    .C(_01538_),
    .X(_01539_));
 sky130_fd_sc_hd__a221o_1 _21527_ (.A1(net4384),
    .A2(_01440_),
    .B1(net416),
    .B2(net4320),
    .C1(net1723),
    .X(_01540_));
 sky130_fd_sc_hd__a22o_1 _21528_ (.A1(\pid_d.curr_int[3] ),
    .A2(net3122),
    .B1(net2077),
    .B2(_01540_),
    .X(_00522_));
 sky130_fd_sc_hd__a31o_1 _21529_ (.A1(\pid_d.prev_int[3] ),
    .A2(_01436_),
    .A3(_01437_),
    .B1(net5982),
    .X(_01541_));
 sky130_fd_sc_hd__o21ai_2 _21530_ (.A1(\pid_d.prev_int[3] ),
    .A2(_01438_),
    .B1(_01541_),
    .Y(_01542_));
 sky130_fd_sc_hd__xor2_1 _21531_ (.A(\pid_d.curr_int[4] ),
    .B(\pid_d.prev_int[4] ),
    .X(_01543_));
 sky130_fd_sc_hd__xnor2_1 _21532_ (.A(_01542_),
    .B(_01543_),
    .Y(_01544_));
 sky130_fd_sc_hd__a21o_1 _21533_ (.A1(net860),
    .A2(net806),
    .B1(_01418_),
    .X(_01545_));
 sky130_fd_sc_hd__o21a_1 _21534_ (.A1(net860),
    .A2(net806),
    .B1(_01545_),
    .X(_01546_));
 sky130_fd_sc_hd__xor2_1 _21535_ (.A(net702),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__nor2_1 _21536_ (.A(_01420_),
    .B(net757),
    .Y(_01548_));
 sky130_fd_sc_hd__a2111o_1 _21537_ (.A1(net705),
    .A2(net703),
    .B1(_01328_),
    .C1(_01548_),
    .D1(net759),
    .X(_01549_));
 sky130_fd_sc_hd__a21o_1 _21538_ (.A1(_01329_),
    .A2(_01423_),
    .B1(_01548_),
    .X(_01550_));
 sky130_fd_sc_hd__nor2_1 _21539_ (.A(net702),
    .B(_01546_),
    .Y(_01551_));
 sky130_fd_sc_hd__a31o_1 _21540_ (.A1(_01547_),
    .A2(net652),
    .A3(_01550_),
    .B1(_01551_),
    .X(_01552_));
 sky130_fd_sc_hd__a21bo_1 _21541_ (.A1(_01501_),
    .A2(net1049),
    .B1_N(net1180),
    .X(_01553_));
 sky130_fd_sc_hd__o21ai_2 _21542_ (.A1(_01501_),
    .A2(net1049),
    .B1(_01553_),
    .Y(_01554_));
 sky130_fd_sc_hd__o21a_1 _21543_ (.A1(_01448_),
    .A2(_01450_),
    .B1(_01449_),
    .X(_01555_));
 sky130_fd_sc_hd__a21oi_2 _21544_ (.A1(_01448_),
    .A2(_01450_),
    .B1(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__nand2_1 _21545_ (.A(net3839),
    .B(net5653),
    .Y(_01557_));
 sky130_fd_sc_hd__nand2_1 _21546_ (.A(net5685),
    .B(net5592),
    .Y(_01558_));
 sky130_fd_sc_hd__nand2_1 _21547_ (.A(net5599),
    .B(net5680),
    .Y(_01559_));
 sky130_fd_sc_hd__xnor2_1 _21548_ (.A(_01558_),
    .B(_01559_),
    .Y(_01560_));
 sky130_fd_sc_hd__xnor2_1 _21549_ (.A(_01557_),
    .B(_01560_),
    .Y(_01561_));
 sky130_fd_sc_hd__nand2_2 _21550_ (.A(net5743),
    .B(net5537),
    .Y(_01562_));
 sky130_fd_sc_hd__nand2_1 _21551_ (.A(net5704),
    .B(net5565),
    .Y(_01563_));
 sky130_fd_sc_hd__nand2_1 _21552_ (.A(net5729),
    .B(net5549),
    .Y(_01564_));
 sky130_fd_sc_hd__xor2_1 _21553_ (.A(_01563_),
    .B(_01564_),
    .X(_01565_));
 sky130_fd_sc_hd__xnor2_2 _21554_ (.A(_01562_),
    .B(_01565_),
    .Y(_01566_));
 sky130_fd_sc_hd__xnor2_1 _21555_ (.A(_01561_),
    .B(_01566_),
    .Y(_01567_));
 sky130_fd_sc_hd__xnor2_1 _21556_ (.A(_01556_),
    .B(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__a21bo_1 _21557_ (.A1(_01454_),
    .A2(_01459_),
    .B1_N(_01452_),
    .X(_01569_));
 sky130_fd_sc_hd__o21a_1 _21558_ (.A1(_01454_),
    .A2(_01459_),
    .B1(_01569_),
    .X(_01570_));
 sky130_fd_sc_hd__nand2_1 _21559_ (.A(net5806),
    .B(net5471),
    .Y(_01571_));
 sky130_fd_sc_hd__nand2_1 _21560_ (.A(net5769),
    .B(net5505),
    .Y(_01572_));
 sky130_fd_sc_hd__nand2_1 _21561_ (.A(net5782),
    .B(net5501),
    .Y(_01573_));
 sky130_fd_sc_hd__xnor2_1 _21562_ (.A(_01572_),
    .B(_01573_),
    .Y(_01574_));
 sky130_fd_sc_hd__xnor2_1 _21563_ (.A(_01571_),
    .B(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__o21a_1 _21564_ (.A1(_01466_),
    .A2(_01468_),
    .B1(_01467_),
    .X(_01576_));
 sky130_fd_sc_hd__a21oi_2 _21565_ (.A1(_01466_),
    .A2(_01468_),
    .B1(_01576_),
    .Y(_01577_));
 sky130_fd_sc_hd__o21a_1 _21566_ (.A1(_01455_),
    .A2(_01457_),
    .B1(_01456_),
    .X(_01578_));
 sky130_fd_sc_hd__a21oi_2 _21567_ (.A1(_01455_),
    .A2(_01457_),
    .B1(_01578_),
    .Y(_01579_));
 sky130_fd_sc_hd__xor2_1 _21568_ (.A(_01577_),
    .B(_01579_),
    .X(_01580_));
 sky130_fd_sc_hd__xnor2_1 _21569_ (.A(_01575_),
    .B(_01580_),
    .Y(_01581_));
 sky130_fd_sc_hd__xor2_1 _21570_ (.A(_01570_),
    .B(_01581_),
    .X(_01582_));
 sky130_fd_sc_hd__xnor2_1 _21571_ (.A(net1722),
    .B(_01582_),
    .Y(_01583_));
 sky130_fd_sc_hd__o21ai_1 _21572_ (.A1(net1727),
    .A2(_01477_),
    .B1(_01478_),
    .Y(_01584_));
 sky130_fd_sc_hd__nand2_1 _21573_ (.A(net5816),
    .B(net5458),
    .Y(_01585_));
 sky130_fd_sc_hd__nand2_1 _21574_ (.A(net5856),
    .B(net5418),
    .Y(_01586_));
 sky130_fd_sc_hd__nand2_1 _21575_ (.A(net5851),
    .B(net5423),
    .Y(_01587_));
 sky130_fd_sc_hd__xnor2_1 _21576_ (.A(_01586_),
    .B(_01587_),
    .Y(_01588_));
 sky130_fd_sc_hd__xnor2_2 _21577_ (.A(_01585_),
    .B(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__o21ai_1 _21578_ (.A1(_01484_),
    .A2(_01485_),
    .B1(_01483_),
    .Y(_01590_));
 sky130_fd_sc_hd__a21bo_1 _21579_ (.A1(_01484_),
    .A2(_01485_),
    .B1_N(_01590_),
    .X(_01591_));
 sky130_fd_sc_hd__xnor2_1 _21580_ (.A(net3818),
    .B(_01490_),
    .Y(_01592_));
 sky130_fd_sc_hd__nand2_2 _21581_ (.A(net5384),
    .B(_01592_),
    .Y(_01593_));
 sky130_fd_sc_hd__xnor2_1 _21582_ (.A(_01591_),
    .B(_01593_),
    .Y(_01594_));
 sky130_fd_sc_hd__xnor2_2 _21583_ (.A(_01589_),
    .B(_01594_),
    .Y(_01595_));
 sky130_fd_sc_hd__a21bo_1 _21584_ (.A1(_01472_),
    .A2(_01474_),
    .B1_N(_01470_),
    .X(_01596_));
 sky130_fd_sc_hd__o21a_1 _21585_ (.A1(_01472_),
    .A2(_01474_),
    .B1(_01596_),
    .X(_01597_));
 sky130_fd_sc_hd__a21o_1 _21586_ (.A1(_01489_),
    .A2(_01493_),
    .B1(_01487_),
    .X(_01598_));
 sky130_fd_sc_hd__o21a_1 _21587_ (.A1(_01489_),
    .A2(_01493_),
    .B1(_01598_),
    .X(_01599_));
 sky130_fd_sc_hd__xnor2_1 _21588_ (.A(net1721),
    .B(_01599_),
    .Y(_01600_));
 sky130_fd_sc_hd__xnor2_2 _21589_ (.A(_01595_),
    .B(_01600_),
    .Y(_01601_));
 sky130_fd_sc_hd__xnor2_1 _21590_ (.A(net1177),
    .B(_01601_),
    .Y(_01602_));
 sky130_fd_sc_hd__xnor2_1 _21591_ (.A(net1178),
    .B(_01602_),
    .Y(_01603_));
 sky130_fd_sc_hd__o21ba_1 _21592_ (.A1(net1725),
    .A2(_01499_),
    .B1_N(_01495_),
    .X(_01604_));
 sky130_fd_sc_hd__a21o_1 _21593_ (.A1(net1725),
    .A2(_01499_),
    .B1(_01604_),
    .X(_01605_));
 sky130_fd_sc_hd__nand2_1 _21594_ (.A(net5892),
    .B(net5400),
    .Y(_01606_));
 sky130_fd_sc_hd__o211a_1 _21595_ (.A1(net5961),
    .A2(net5943),
    .B1(net5921),
    .C1(net3115),
    .X(_01607_));
 sky130_fd_sc_hd__a21o_1 _21596_ (.A1(net5928),
    .A2(net5909),
    .B1(net5951),
    .X(_01608_));
 sky130_fd_sc_hd__and2_1 _21597_ (.A(net3806),
    .B(_01608_),
    .X(_01609_));
 sky130_fd_sc_hd__nand2_1 _21598_ (.A(net5383),
    .B(net3106),
    .Y(_01610_));
 sky130_fd_sc_hd__a22o_1 _21599_ (.A1(net5383),
    .A2(_01607_),
    .B1(_01610_),
    .B2(net5897),
    .X(_01611_));
 sky130_fd_sc_hd__a32o_1 _21600_ (.A1(net5383),
    .A2(net3803),
    .A3(_01606_),
    .B1(_01611_),
    .B2(net5400),
    .X(_01612_));
 sky130_fd_sc_hd__and3_1 _21601_ (.A(net5416),
    .B(net5893),
    .C(_01513_),
    .X(_01613_));
 sky130_fd_sc_hd__xnor2_1 _21602_ (.A(_01612_),
    .B(_01613_),
    .Y(_01614_));
 sky130_fd_sc_hd__xnor2_2 _21603_ (.A(_01605_),
    .B(_01614_),
    .Y(_01615_));
 sky130_fd_sc_hd__xor2_1 _21604_ (.A(_01603_),
    .B(_01615_),
    .X(_01616_));
 sky130_fd_sc_hd__xnor2_1 _21605_ (.A(_01554_),
    .B(_01616_),
    .Y(_01617_));
 sky130_fd_sc_hd__o21ba_1 _21606_ (.A1(net948),
    .A2(_01515_),
    .B1_N(net947),
    .X(_01618_));
 sky130_fd_sc_hd__a21o_1 _21607_ (.A1(net948),
    .A2(_01515_),
    .B1(_01618_),
    .X(_01619_));
 sky130_fd_sc_hd__a21oi_1 _21608_ (.A1(net5416),
    .A2(net5893),
    .B1(_01513_),
    .Y(_01620_));
 sky130_fd_sc_hd__or2_1 _21609_ (.A(_01613_),
    .B(_01620_),
    .X(_01621_));
 sky130_fd_sc_hd__a21o_1 _21610_ (.A1(net5427),
    .A2(net5888),
    .B1(_01508_),
    .X(_01622_));
 sky130_fd_sc_hd__o2bb2a_1 _21611_ (.A1_N(_01506_),
    .A2_N(_01622_),
    .B1(_01621_),
    .B2(net1179),
    .X(_01623_));
 sky130_fd_sc_hd__a21oi_1 _21612_ (.A1(net1179),
    .A2(_01621_),
    .B1(_01623_),
    .Y(_01624_));
 sky130_fd_sc_hd__nand2_1 _21613_ (.A(_01619_),
    .B(_01624_),
    .Y(_01625_));
 sky130_fd_sc_hd__or2_1 _21614_ (.A(_01619_),
    .B(_01624_),
    .X(_01626_));
 sky130_fd_sc_hd__nand2_1 _21615_ (.A(_01625_),
    .B(_01626_),
    .Y(_01627_));
 sky130_fd_sc_hd__xor2_1 _21616_ (.A(_01617_),
    .B(_01627_),
    .X(_01628_));
 sky130_fd_sc_hd__a21o_1 _21617_ (.A1(_01447_),
    .A2(_01519_),
    .B1(_01442_),
    .X(_01629_));
 sky130_fd_sc_hd__o21a_1 _21618_ (.A1(_01447_),
    .A2(_01519_),
    .B1(_01629_),
    .X(_01630_));
 sky130_fd_sc_hd__or2_1 _21619_ (.A(_01628_),
    .B(net701),
    .X(_01631_));
 sky130_fd_sc_hd__and2_1 _21620_ (.A(_01628_),
    .B(net701),
    .X(_01632_));
 sky130_fd_sc_hd__inv_2 _21621_ (.A(_01632_),
    .Y(_01633_));
 sky130_fd_sc_hd__nand2_1 _21622_ (.A(_01631_),
    .B(_01633_),
    .Y(_01634_));
 sky130_fd_sc_hd__xnor2_1 _21623_ (.A(net600),
    .B(_01634_),
    .Y(_01635_));
 sky130_fd_sc_hd__inv_2 _21624_ (.A(net5970),
    .Y(_01636_));
 sky130_fd_sc_hd__o21ba_1 _21625_ (.A1(_01636_),
    .A2(_01535_),
    .B1_N(\pid_d.prev_error[3] ),
    .X(_01637_));
 sky130_fd_sc_hd__a21o_1 _21626_ (.A1(_01636_),
    .A2(_01535_),
    .B1(_01637_),
    .X(_01638_));
 sky130_fd_sc_hd__xnor2_1 _21627_ (.A(\pid_d.prev_error[4] ),
    .B(\pid_d.curr_error[4] ),
    .Y(_01639_));
 sky130_fd_sc_hd__nand2_1 _21628_ (.A(_01638_),
    .B(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hd__or2_1 _21629_ (.A(_01638_),
    .B(_01639_),
    .X(_01641_));
 sky130_fd_sc_hd__and3_1 _21630_ (.A(net4357),
    .B(_01640_),
    .C(_01641_),
    .X(_01642_));
 sky130_fd_sc_hd__a221o_1 _21631_ (.A1(net4385),
    .A2(_01544_),
    .B1(net476),
    .B2(net4318),
    .C1(net1175),
    .X(_01643_));
 sky130_fd_sc_hd__a22o_1 _21632_ (.A1(\pid_d.curr_int[4] ),
    .A2(net3122),
    .B1(net2077),
    .B2(_01643_),
    .X(_00523_));
 sky130_fd_sc_hd__inv_2 _21633_ (.A(\pid_d.prev_int[4] ),
    .Y(_01644_));
 sky130_fd_sc_hd__o21ba_1 _21634_ (.A1(_01644_),
    .A2(_01542_),
    .B1_N(\pid_d.curr_int[4] ),
    .X(_01645_));
 sky130_fd_sc_hd__a21o_1 _21635_ (.A1(_01644_),
    .A2(_01542_),
    .B1(_01645_),
    .X(_01646_));
 sky130_fd_sc_hd__xor2_1 _21636_ (.A(\pid_d.curr_int[5] ),
    .B(\pid_d.prev_int[5] ),
    .X(_01647_));
 sky130_fd_sc_hd__xnor2_1 _21637_ (.A(_01646_),
    .B(_01647_),
    .Y(_01648_));
 sky130_fd_sc_hd__a21o_1 _21638_ (.A1(net600),
    .A2(_01631_),
    .B1(_01632_),
    .X(_01649_));
 sky130_fd_sc_hd__nand2_1 _21639_ (.A(_01554_),
    .B(_01615_),
    .Y(_01650_));
 sky130_fd_sc_hd__nor2_1 _21640_ (.A(_01554_),
    .B(_01615_),
    .Y(_01651_));
 sky130_fd_sc_hd__a21o_1 _21641_ (.A1(_01603_),
    .A2(_01650_),
    .B1(_01651_),
    .X(_01652_));
 sky130_fd_sc_hd__o21ba_1 _21642_ (.A1(net1177),
    .A2(_01601_),
    .B1_N(net1178),
    .X(_01653_));
 sky130_fd_sc_hd__a21o_1 _21643_ (.A1(net1177),
    .A2(_01601_),
    .B1(_01653_),
    .X(_01654_));
 sky130_fd_sc_hd__a21bo_1 _21644_ (.A1(_01570_),
    .A2(_01581_),
    .B1_N(net1722),
    .X(_01655_));
 sky130_fd_sc_hd__o21a_1 _21645_ (.A1(_01570_),
    .A2(_01581_),
    .B1(_01655_),
    .X(_01656_));
 sky130_fd_sc_hd__a21bo_1 _21646_ (.A1(_01556_),
    .A2(_01566_),
    .B1_N(_01561_),
    .X(_01657_));
 sky130_fd_sc_hd__o21ai_2 _21647_ (.A1(_01556_),
    .A2(_01566_),
    .B1(_01657_),
    .Y(_01658_));
 sky130_fd_sc_hd__o21a_1 _21648_ (.A1(_01557_),
    .A2(_01559_),
    .B1(_01558_),
    .X(_01659_));
 sky130_fd_sc_hd__a21oi_2 _21649_ (.A1(_01557_),
    .A2(_01559_),
    .B1(_01659_),
    .Y(_01660_));
 sky130_fd_sc_hd__nand2b_1 _21650_ (.A_N(net5609),
    .B(net5653),
    .Y(_01661_));
 sky130_fd_sc_hd__nand2_1 _21651_ (.A(net5688),
    .B(net5566),
    .Y(_01662_));
 sky130_fd_sc_hd__nand2_1 _21652_ (.A(net5593),
    .B(net5680),
    .Y(_01663_));
 sky130_fd_sc_hd__xnor2_1 _21653_ (.A(_01662_),
    .B(_01663_),
    .Y(_01664_));
 sky130_fd_sc_hd__xnor2_1 _21654_ (.A(_01661_),
    .B(_01664_),
    .Y(_01665_));
 sky130_fd_sc_hd__nand2_1 _21655_ (.A(net5744),
    .B(net5516),
    .Y(_01666_));
 sky130_fd_sc_hd__nand2_1 _21656_ (.A(net5704),
    .B(net5550),
    .Y(_01667_));
 sky130_fd_sc_hd__nand2_1 _21657_ (.A(net5718),
    .B(net5538),
    .Y(_01668_));
 sky130_fd_sc_hd__xor2_1 _21658_ (.A(_01667_),
    .B(_01668_),
    .X(_01669_));
 sky130_fd_sc_hd__xnor2_2 _21659_ (.A(_01666_),
    .B(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__xor2_1 _21660_ (.A(_01665_),
    .B(_01670_),
    .X(_01671_));
 sky130_fd_sc_hd__xnor2_1 _21661_ (.A(_01660_),
    .B(_01671_),
    .Y(_01672_));
 sky130_fd_sc_hd__nand2_2 _21662_ (.A(net5783),
    .B(net5484),
    .Y(_01673_));
 sky130_fd_sc_hd__nand2_1 _21663_ (.A(net5768),
    .B(net5502),
    .Y(_01674_));
 sky130_fd_sc_hd__nand2_1 _21664_ (.A(net5798),
    .B(net5460),
    .Y(_01675_));
 sky130_fd_sc_hd__xnor2_1 _21665_ (.A(_01674_),
    .B(_01675_),
    .Y(_01676_));
 sky130_fd_sc_hd__xnor2_2 _21666_ (.A(_01673_),
    .B(_01676_),
    .Y(_01677_));
 sky130_fd_sc_hd__nand2_1 _21667_ (.A(_01562_),
    .B(_01564_),
    .Y(_01678_));
 sky130_fd_sc_hd__nor2_1 _21668_ (.A(_01562_),
    .B(_01564_),
    .Y(_01679_));
 sky130_fd_sc_hd__a31o_1 _21669_ (.A1(net5701),
    .A2(net5572),
    .A3(_01678_),
    .B1(_01679_),
    .X(_01680_));
 sky130_fd_sc_hd__nand2_1 _21670_ (.A(_01571_),
    .B(_01573_),
    .Y(_01681_));
 sky130_fd_sc_hd__nor2_1 _21671_ (.A(_01571_),
    .B(_01573_),
    .Y(_01682_));
 sky130_fd_sc_hd__a31o_1 _21672_ (.A1(net5769),
    .A2(net5505),
    .A3(_01681_),
    .B1(_01682_),
    .X(_01683_));
 sky130_fd_sc_hd__xnor2_1 _21673_ (.A(_01680_),
    .B(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__xnor2_2 _21674_ (.A(_01677_),
    .B(_01684_),
    .Y(_01685_));
 sky130_fd_sc_hd__xnor2_1 _21675_ (.A(_01672_),
    .B(_01685_),
    .Y(_01686_));
 sky130_fd_sc_hd__xnor2_1 _21676_ (.A(_01658_),
    .B(_01686_),
    .Y(_01687_));
 sky130_fd_sc_hd__o21ai_1 _21677_ (.A1(_01586_),
    .A2(_01587_),
    .B1(_01585_),
    .Y(_01688_));
 sky130_fd_sc_hd__a21bo_1 _21678_ (.A1(_01586_),
    .A2(_01587_),
    .B1_N(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__nand2_1 _21679_ (.A(net5859),
    .B(net5401),
    .Y(_01690_));
 sky130_fd_sc_hd__nand2_1 _21680_ (.A(net5842),
    .B(net5413),
    .Y(_01691_));
 sky130_fd_sc_hd__nand2_1 _21681_ (.A(net5813),
    .B(net5440),
    .Y(_01692_));
 sky130_fd_sc_hd__xnor2_1 _21682_ (.A(_01691_),
    .B(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__xnor2_1 _21683_ (.A(_01690_),
    .B(_01693_),
    .Y(_01694_));
 sky130_fd_sc_hd__nor2_1 _21684_ (.A(_01689_),
    .B(_01694_),
    .Y(_01695_));
 sky130_fd_sc_hd__nand2_1 _21685_ (.A(_01689_),
    .B(_01694_),
    .Y(_01696_));
 sky130_fd_sc_hd__or2b_1 _21686_ (.A(_01695_),
    .B_N(_01696_),
    .X(_01697_));
 sky130_fd_sc_hd__xnor2_2 _21687_ (.A(_01593_),
    .B(_01697_),
    .Y(_01698_));
 sky130_fd_sc_hd__a21bo_1 _21688_ (.A1(_01577_),
    .A2(_01579_),
    .B1_N(_01575_),
    .X(_01699_));
 sky130_fd_sc_hd__o21a_1 _21689_ (.A1(_01577_),
    .A2(_01579_),
    .B1(_01699_),
    .X(_01700_));
 sky130_fd_sc_hd__o21a_1 _21690_ (.A1(_01591_),
    .A2(_01593_),
    .B1(_01589_),
    .X(_01701_));
 sky130_fd_sc_hd__a21oi_1 _21691_ (.A1(_01591_),
    .A2(_01593_),
    .B1(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__nor2_1 _21692_ (.A(net1720),
    .B(_01702_),
    .Y(_01703_));
 sky130_fd_sc_hd__nand2_1 _21693_ (.A(net1720),
    .B(_01702_),
    .Y(_01704_));
 sky130_fd_sc_hd__and2b_1 _21694_ (.A_N(_01703_),
    .B(_01704_),
    .X(_01705_));
 sky130_fd_sc_hd__xnor2_2 _21695_ (.A(_01698_),
    .B(_01705_),
    .Y(_01706_));
 sky130_fd_sc_hd__xor2_1 _21696_ (.A(net1173),
    .B(_01706_),
    .X(_01707_));
 sky130_fd_sc_hd__xnor2_1 _21697_ (.A(net1174),
    .B(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hd__inv_2 _21698_ (.A(net5396),
    .Y(_01709_));
 sky130_fd_sc_hd__o21ai_1 _21699_ (.A1(net5891),
    .A2(net3107),
    .B1(net5384),
    .Y(_01710_));
 sky130_fd_sc_hd__a31o_1 _21700_ (.A1(net5896),
    .A2(net3785),
    .A3(net3107),
    .B1(_01710_),
    .X(_01711_));
 sky130_fd_sc_hd__o21ba_1 _21701_ (.A1(net1721),
    .A2(_01599_),
    .B1_N(_01595_),
    .X(_01712_));
 sky130_fd_sc_hd__a21oi_1 _21702_ (.A1(net1721),
    .A2(_01599_),
    .B1(_01712_),
    .Y(_01713_));
 sky130_fd_sc_hd__nor2_1 _21703_ (.A(net2069),
    .B(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__and2_1 _21704_ (.A(net2069),
    .B(_01713_),
    .X(_01715_));
 sky130_fd_sc_hd__or2_1 _21705_ (.A(_01714_),
    .B(_01715_),
    .X(_01716_));
 sky130_fd_sc_hd__xor2_1 _21706_ (.A(_01708_),
    .B(_01716_),
    .X(_01717_));
 sky130_fd_sc_hd__xnor2_2 _21707_ (.A(_01654_),
    .B(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__a21bo_1 _21708_ (.A1(_01612_),
    .A2(_01613_),
    .B1_N(_01605_),
    .X(_01719_));
 sky130_fd_sc_hd__o21a_1 _21709_ (.A1(_01612_),
    .A2(_01613_),
    .B1(_01719_),
    .X(_01720_));
 sky130_fd_sc_hd__xnor2_1 _21710_ (.A(_01718_),
    .B(_01720_),
    .Y(_01721_));
 sky130_fd_sc_hd__xnor2_1 _21711_ (.A(_01652_),
    .B(_01721_),
    .Y(_01722_));
 sky130_fd_sc_hd__nand2_1 _21712_ (.A(_01617_),
    .B(_01625_),
    .Y(_01723_));
 sky130_fd_sc_hd__and3_1 _21713_ (.A(_01626_),
    .B(_01722_),
    .C(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__a21o_1 _21714_ (.A1(_01626_),
    .A2(_01723_),
    .B1(_01722_),
    .X(_01725_));
 sky130_fd_sc_hd__and2b_1 _21715_ (.A_N(_01724_),
    .B(_01725_),
    .X(_01726_));
 sky130_fd_sc_hd__xor2_1 _21716_ (.A(_01649_),
    .B(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__inv_2 _21717_ (.A(\pid_d.curr_error[4] ),
    .Y(_01728_));
 sky130_fd_sc_hd__o21ba_1 _21718_ (.A1(_01728_),
    .A2(_01638_),
    .B1_N(\pid_d.prev_error[4] ),
    .X(_01729_));
 sky130_fd_sc_hd__a21o_1 _21719_ (.A1(_01728_),
    .A2(_01638_),
    .B1(_01729_),
    .X(_01730_));
 sky130_fd_sc_hd__xnor2_1 _21720_ (.A(\pid_d.prev_error[5] ),
    .B(net5969),
    .Y(_01731_));
 sky130_fd_sc_hd__nand2_1 _21721_ (.A(_01730_),
    .B(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__or2_1 _21722_ (.A(_01730_),
    .B(_01731_),
    .X(_01733_));
 sky130_fd_sc_hd__and3_1 _21723_ (.A(net4358),
    .B(_01732_),
    .C(_01733_),
    .X(_01734_));
 sky130_fd_sc_hd__a221o_1 _21724_ (.A1(net4385),
    .A2(_01648_),
    .B1(net524),
    .B2(net4318),
    .C1(net946),
    .X(_01735_));
 sky130_fd_sc_hd__a22o_1 _21725_ (.A1(\pid_d.curr_int[5] ),
    .A2(net3123),
    .B1(net2078),
    .B2(_01735_),
    .X(_00524_));
 sky130_fd_sc_hd__inv_2 _21726_ (.A(\pid_d.prev_int[5] ),
    .Y(_01736_));
 sky130_fd_sc_hd__o21ba_1 _21727_ (.A1(_01736_),
    .A2(_01646_),
    .B1_N(\pid_d.curr_int[5] ),
    .X(_01737_));
 sky130_fd_sc_hd__a21o_1 _21728_ (.A1(_01736_),
    .A2(_01646_),
    .B1(_01737_),
    .X(_01738_));
 sky130_fd_sc_hd__xor2_1 _21729_ (.A(\pid_d.curr_int[6] ),
    .B(\pid_d.prev_int[6] ),
    .X(_01739_));
 sky130_fd_sc_hd__xnor2_1 _21730_ (.A(_01738_),
    .B(_01739_),
    .Y(_01740_));
 sky130_fd_sc_hd__a21o_1 _21731_ (.A1(_01654_),
    .A2(_01716_),
    .B1(_01708_),
    .X(_01741_));
 sky130_fd_sc_hd__o21a_2 _21732_ (.A1(_01654_),
    .A2(_01716_),
    .B1(_01741_),
    .X(_01742_));
 sky130_fd_sc_hd__a21o_1 _21733_ (.A1(net1173),
    .A2(_01706_),
    .B1(net1174),
    .X(_01743_));
 sky130_fd_sc_hd__o21a_2 _21734_ (.A1(net1173),
    .A2(_01706_),
    .B1(_01743_),
    .X(_01744_));
 sky130_fd_sc_hd__o21ba_1 _21735_ (.A1(_01658_),
    .A2(_01685_),
    .B1_N(_01672_),
    .X(_01745_));
 sky130_fd_sc_hd__a21o_1 _21736_ (.A1(_01658_),
    .A2(_01685_),
    .B1(_01745_),
    .X(_01746_));
 sky130_fd_sc_hd__a21bo_1 _21737_ (.A1(_01660_),
    .A2(_01670_),
    .B1_N(_01665_),
    .X(_01747_));
 sky130_fd_sc_hd__o21a_1 _21738_ (.A1(_01660_),
    .A2(_01670_),
    .B1(_01747_),
    .X(_01748_));
 sky130_fd_sc_hd__nand2_1 _21739_ (.A(_01135_),
    .B(net5645),
    .Y(_01749_));
 sky130_fd_sc_hd__nand2_1 _21740_ (.A(net5686),
    .B(net5551),
    .Y(_01750_));
 sky130_fd_sc_hd__nand2_1 _21741_ (.A(net5567),
    .B(net5679),
    .Y(_01751_));
 sky130_fd_sc_hd__xnor2_1 _21742_ (.A(_01750_),
    .B(_01751_),
    .Y(_01752_));
 sky130_fd_sc_hd__xnor2_1 _21743_ (.A(_01749_),
    .B(_01752_),
    .Y(_01753_));
 sky130_fd_sc_hd__o21a_1 _21744_ (.A1(_01661_),
    .A2(_01663_),
    .B1(_01662_),
    .X(_01754_));
 sky130_fd_sc_hd__a21oi_2 _21745_ (.A1(_01661_),
    .A2(_01663_),
    .B1(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hd__nand2_1 _21746_ (.A(net5742),
    .B(net5500),
    .Y(_01756_));
 sky130_fd_sc_hd__nand2_1 _21747_ (.A(net5703),
    .B(net5538),
    .Y(_01757_));
 sky130_fd_sc_hd__nand2_1 _21748_ (.A(net5725),
    .B(net5515),
    .Y(_01758_));
 sky130_fd_sc_hd__xor2_1 _21749_ (.A(_01757_),
    .B(_01758_),
    .X(_01759_));
 sky130_fd_sc_hd__xnor2_2 _21750_ (.A(_01756_),
    .B(_01759_),
    .Y(_01760_));
 sky130_fd_sc_hd__xnor2_1 _21751_ (.A(_01755_),
    .B(_01760_),
    .Y(_01761_));
 sky130_fd_sc_hd__xnor2_1 _21752_ (.A(_01753_),
    .B(_01761_),
    .Y(_01762_));
 sky130_fd_sc_hd__and2_1 _21753_ (.A(net5765),
    .B(net5485),
    .X(_01763_));
 sky130_fd_sc_hd__nand2_1 _21754_ (.A(net5801),
    .B(net5431),
    .Y(_01764_));
 sky130_fd_sc_hd__nand2_1 _21755_ (.A(net5785),
    .B(net5461),
    .Y(_01765_));
 sky130_fd_sc_hd__xor2_1 _21756_ (.A(_01764_),
    .B(_01765_),
    .X(_01766_));
 sky130_fd_sc_hd__xnor2_2 _21757_ (.A(_01763_),
    .B(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__nand2_1 _21758_ (.A(_01666_),
    .B(_01668_),
    .Y(_01768_));
 sky130_fd_sc_hd__nor2_1 _21759_ (.A(_01666_),
    .B(_01668_),
    .Y(_01769_));
 sky130_fd_sc_hd__a31o_1 _21760_ (.A1(net5706),
    .A2(net5549),
    .A3(_01768_),
    .B1(_01769_),
    .X(_01770_));
 sky130_fd_sc_hd__nand2_1 _21761_ (.A(_01673_),
    .B(_01675_),
    .Y(_01771_));
 sky130_fd_sc_hd__nor2_1 _21762_ (.A(_01673_),
    .B(_01675_),
    .Y(_01772_));
 sky130_fd_sc_hd__a31o_1 _21763_ (.A1(net5768),
    .A2(net5502),
    .A3(_01771_),
    .B1(_01772_),
    .X(_01773_));
 sky130_fd_sc_hd__xor2_1 _21764_ (.A(_01770_),
    .B(_01773_),
    .X(_01774_));
 sky130_fd_sc_hd__xnor2_2 _21765_ (.A(_01767_),
    .B(_01774_),
    .Y(_01775_));
 sky130_fd_sc_hd__xnor2_1 _21766_ (.A(_01762_),
    .B(_01775_),
    .Y(_01776_));
 sky130_fd_sc_hd__xnor2_1 _21767_ (.A(_01748_),
    .B(_01776_),
    .Y(_01777_));
 sky130_fd_sc_hd__and2_1 _21768_ (.A(net5384),
    .B(_01592_),
    .X(_01778_));
 sky130_fd_sc_hd__buf_1 _21769_ (.A(_01778_),
    .X(_01779_));
 sky130_fd_sc_hd__o21ai_2 _21770_ (.A1(_01779_),
    .A2(_01695_),
    .B1(_01696_),
    .Y(_01780_));
 sky130_fd_sc_hd__nand2_1 _21771_ (.A(net5857),
    .B(net5376),
    .Y(_01781_));
 sky130_fd_sc_hd__nand2_1 _21772_ (.A(net5812),
    .B(net5406),
    .Y(_01782_));
 sky130_fd_sc_hd__nand2_1 _21773_ (.A(net5839),
    .B(net5394),
    .Y(_01783_));
 sky130_fd_sc_hd__xnor2_1 _21774_ (.A(_01782_),
    .B(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__xnor2_1 _21775_ (.A(_01781_),
    .B(_01784_),
    .Y(_01785_));
 sky130_fd_sc_hd__o21a_1 _21776_ (.A1(_01690_),
    .A2(_01691_),
    .B1(_01692_),
    .X(_01786_));
 sky130_fd_sc_hd__a21o_1 _21777_ (.A1(_01690_),
    .A2(_01691_),
    .B1(_01786_),
    .X(_01787_));
 sky130_fd_sc_hd__xor2_1 _21778_ (.A(net2475),
    .B(_01787_),
    .X(_01788_));
 sky130_fd_sc_hd__o21ba_1 _21779_ (.A1(_01680_),
    .A2(_01683_),
    .B1_N(_01677_),
    .X(_01789_));
 sky130_fd_sc_hd__a21oi_2 _21780_ (.A1(_01680_),
    .A2(_01683_),
    .B1(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__xnor2_1 _21781_ (.A(_01788_),
    .B(_01790_),
    .Y(_01791_));
 sky130_fd_sc_hd__xnor2_1 _21782_ (.A(_01780_),
    .B(_01791_),
    .Y(_01792_));
 sky130_fd_sc_hd__xnor2_1 _21783_ (.A(net1172),
    .B(_01792_),
    .Y(_01793_));
 sky130_fd_sc_hd__xnor2_2 _21784_ (.A(net1048),
    .B(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__a21o_1 _21785_ (.A1(_01698_),
    .A2(_01704_),
    .B1(_01703_),
    .X(_01795_));
 sky130_fd_sc_hd__buf_1 _21786_ (.A(_01593_),
    .X(_01796_));
 sky130_fd_sc_hd__o21a_1 _21787_ (.A1(net5896),
    .A2(net3108),
    .B1(net5385),
    .X(_01797_));
 sky130_fd_sc_hd__clkbuf_1 _21788_ (.A(_01797_),
    .X(_01798_));
 sky130_fd_sc_hd__xnor2_2 _21789_ (.A(_01796_),
    .B(net2063),
    .Y(_01799_));
 sky130_fd_sc_hd__xor2_1 _21790_ (.A(_01795_),
    .B(_01799_),
    .X(_01800_));
 sky130_fd_sc_hd__xnor2_1 _21791_ (.A(_01794_),
    .B(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hd__xnor2_2 _21792_ (.A(_01744_),
    .B(_01801_),
    .Y(_01802_));
 sky130_fd_sc_hd__xnor2_1 _21793_ (.A(_01714_),
    .B(_01802_),
    .Y(_01803_));
 sky130_fd_sc_hd__xnor2_2 _21794_ (.A(_01742_),
    .B(_01803_),
    .Y(_01804_));
 sky130_fd_sc_hd__a21o_1 _21795_ (.A1(_01718_),
    .A2(_01720_),
    .B1(_01652_),
    .X(_01805_));
 sky130_fd_sc_hd__o21a_1 _21796_ (.A1(_01718_),
    .A2(_01720_),
    .B1(_01805_),
    .X(_01806_));
 sky130_fd_sc_hd__xor2_1 _21797_ (.A(_01804_),
    .B(_01806_),
    .X(_01807_));
 sky130_fd_sc_hd__a21oi_1 _21798_ (.A1(_01649_),
    .A2(_01725_),
    .B1(_01724_),
    .Y(_01808_));
 sky130_fd_sc_hd__xnor2_1 _21799_ (.A(_01807_),
    .B(_01808_),
    .Y(_01809_));
 sky130_fd_sc_hd__inv_2 _21800_ (.A(net5969),
    .Y(_01810_));
 sky130_fd_sc_hd__o21ba_1 _21801_ (.A1(_01810_),
    .A2(_01730_),
    .B1_N(\pid_d.prev_error[5] ),
    .X(_01811_));
 sky130_fd_sc_hd__a21o_1 _21802_ (.A1(_01810_),
    .A2(_01730_),
    .B1(_01811_),
    .X(_01812_));
 sky130_fd_sc_hd__xnor2_1 _21803_ (.A(\pid_d.prev_error[6] ),
    .B(net5968),
    .Y(_01813_));
 sky130_fd_sc_hd__nand2_1 _21804_ (.A(_01812_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__or2_1 _21805_ (.A(_01812_),
    .B(_01813_),
    .X(_01815_));
 sky130_fd_sc_hd__and3_1 _21806_ (.A(net4358),
    .B(_01814_),
    .C(_01815_),
    .X(_01816_));
 sky130_fd_sc_hd__a221o_1 _21807_ (.A1(net4385),
    .A2(_01740_),
    .B1(net473),
    .B2(net4319),
    .C1(net804),
    .X(_01817_));
 sky130_fd_sc_hd__a22o_1 _21808_ (.A1(net9243),
    .A2(net3123),
    .B1(net2078),
    .B2(_01817_),
    .X(_00525_));
 sky130_fd_sc_hd__inv_2 _21809_ (.A(\pid_d.prev_int[6] ),
    .Y(_01818_));
 sky130_fd_sc_hd__inv_2 _21810_ (.A(net5979),
    .Y(_01819_));
 sky130_fd_sc_hd__o21a_1 _21811_ (.A1(_01818_),
    .A2(_01738_),
    .B1(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__a21o_1 _21812_ (.A1(_01818_),
    .A2(_01738_),
    .B1(_01820_),
    .X(_01821_));
 sky130_fd_sc_hd__xor2_1 _21813_ (.A(net5978),
    .B(\pid_d.prev_int[7] ),
    .X(_01822_));
 sky130_fd_sc_hd__xnor2_1 _21814_ (.A(_01821_),
    .B(_01822_),
    .Y(_01823_));
 sky130_fd_sc_hd__a211o_1 _21815_ (.A1(net600),
    .A2(_01631_),
    .B1(_01632_),
    .C1(_01724_),
    .X(_01824_));
 sky130_fd_sc_hd__a22o_1 _21816_ (.A1(_01804_),
    .A2(_01806_),
    .B1(_01824_),
    .B2(_01725_),
    .X(_01825_));
 sky130_fd_sc_hd__or2_1 _21817_ (.A(_01804_),
    .B(_01806_),
    .X(_01826_));
 sky130_fd_sc_hd__nand2_1 _21818_ (.A(_01825_),
    .B(_01826_),
    .Y(_01827_));
 sky130_fd_sc_hd__a21bo_1 _21819_ (.A1(_01748_),
    .A2(_01775_),
    .B1_N(_01762_),
    .X(_01828_));
 sky130_fd_sc_hd__o21ai_1 _21820_ (.A1(_01748_),
    .A2(_01775_),
    .B1(_01828_),
    .Y(_01829_));
 sky130_fd_sc_hd__o21a_1 _21821_ (.A1(_01749_),
    .A2(_01751_),
    .B1(_01750_),
    .X(_01830_));
 sky130_fd_sc_hd__a21oi_1 _21822_ (.A1(_01749_),
    .A2(_01751_),
    .B1(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__nand2_2 _21823_ (.A(_01066_),
    .B(net5645),
    .Y(_01832_));
 sky130_fd_sc_hd__nand2_1 _21824_ (.A(net5686),
    .B(net5539),
    .Y(_01833_));
 sky130_fd_sc_hd__nand2_1 _21825_ (.A(net5548),
    .B(net5679),
    .Y(_01834_));
 sky130_fd_sc_hd__xnor2_1 _21826_ (.A(_01833_),
    .B(_01834_),
    .Y(_01835_));
 sky130_fd_sc_hd__xnor2_2 _21827_ (.A(_01832_),
    .B(_01835_),
    .Y(_01836_));
 sky130_fd_sc_hd__nand2_2 _21828_ (.A(net5750),
    .B(net5479),
    .Y(_01837_));
 sky130_fd_sc_hd__nand2_1 _21829_ (.A(net5703),
    .B(net5515),
    .Y(_01838_));
 sky130_fd_sc_hd__nand2_1 _21830_ (.A(net5719),
    .B(net5499),
    .Y(_01839_));
 sky130_fd_sc_hd__xnor2_1 _21831_ (.A(_01838_),
    .B(_01839_),
    .Y(_01840_));
 sky130_fd_sc_hd__xnor2_2 _21832_ (.A(_01837_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__xor2_1 _21833_ (.A(_01836_),
    .B(_01841_),
    .X(_01842_));
 sky130_fd_sc_hd__xnor2_1 _21834_ (.A(_01831_),
    .B(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__a21bo_1 _21835_ (.A1(_01755_),
    .A2(_01760_),
    .B1_N(_01753_),
    .X(_01844_));
 sky130_fd_sc_hd__o21a_1 _21836_ (.A1(_01755_),
    .A2(_01760_),
    .B1(_01844_),
    .X(_01845_));
 sky130_fd_sc_hd__and2_1 _21837_ (.A(net5764),
    .B(net5461),
    .X(_01846_));
 sky130_fd_sc_hd__nand2_1 _21838_ (.A(net5801),
    .B(net5408),
    .Y(_01847_));
 sky130_fd_sc_hd__nand2_1 _21839_ (.A(net5784),
    .B(net5431),
    .Y(_01848_));
 sky130_fd_sc_hd__xor2_1 _21840_ (.A(_01847_),
    .B(_01848_),
    .X(_01849_));
 sky130_fd_sc_hd__xnor2_2 _21841_ (.A(_01846_),
    .B(_01849_),
    .Y(_01850_));
 sky130_fd_sc_hd__o21a_1 _21842_ (.A1(_01756_),
    .A2(_01758_),
    .B1(_01757_),
    .X(_01851_));
 sky130_fd_sc_hd__a21oi_1 _21843_ (.A1(_01756_),
    .A2(_01758_),
    .B1(_01851_),
    .Y(_01852_));
 sky130_fd_sc_hd__o21ba_1 _21844_ (.A1(_01764_),
    .A2(_01765_),
    .B1_N(_01763_),
    .X(_01853_));
 sky130_fd_sc_hd__a21oi_1 _21845_ (.A1(_01764_),
    .A2(_01765_),
    .B1(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__xor2_1 _21846_ (.A(net2474),
    .B(_01854_),
    .X(_01855_));
 sky130_fd_sc_hd__xnor2_2 _21847_ (.A(_01850_),
    .B(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__xnor2_1 _21848_ (.A(_01845_),
    .B(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__xnor2_1 _21849_ (.A(net1719),
    .B(_01857_),
    .Y(_01858_));
 sky130_fd_sc_hd__o21a_1 _21850_ (.A1(net2475),
    .A2(_01787_),
    .B1(net2064),
    .X(_01859_));
 sky130_fd_sc_hd__a21o_1 _21851_ (.A1(net2475),
    .A2(_01787_),
    .B1(_01859_),
    .X(_01860_));
 sky130_fd_sc_hd__o21ba_1 _21852_ (.A1(_01770_),
    .A2(_01773_),
    .B1_N(_01767_),
    .X(_01861_));
 sky130_fd_sc_hd__a21oi_2 _21853_ (.A1(_01770_),
    .A2(_01773_),
    .B1(_01861_),
    .Y(_01862_));
 sky130_fd_sc_hd__inv_2 _21854_ (.A(net5809),
    .Y(_01863_));
 sky130_fd_sc_hd__and2b_1 _21855_ (.A_N(net5406),
    .B(net5857),
    .X(_01864_));
 sky130_fd_sc_hd__o22a_1 _21856_ (.A1(net5406),
    .A2(net5376),
    .B1(_01864_),
    .B2(net5839),
    .X(_01865_));
 sky130_fd_sc_hd__inv_2 _21857_ (.A(net5839),
    .Y(_01866_));
 sky130_fd_sc_hd__a21bo_1 _21858_ (.A1(_01866_),
    .A2(net5857),
    .B1_N(_01783_),
    .X(_01867_));
 sky130_fd_sc_hd__inv_2 _21859_ (.A(_01867_),
    .Y(_01868_));
 sky130_fd_sc_hd__nor2_1 _21860_ (.A(net5406),
    .B(net3786),
    .Y(_01869_));
 sky130_fd_sc_hd__o22a_1 _21861_ (.A1(net5394),
    .A2(_01782_),
    .B1(_01869_),
    .B2(net5857),
    .X(_01870_));
 sky130_fd_sc_hd__or3b_1 _21862_ (.A(net5839),
    .B(net5394),
    .C_N(_01864_),
    .X(_01871_));
 sky130_fd_sc_hd__o221a_1 _21863_ (.A1(net5812),
    .A2(_01868_),
    .B1(_01870_),
    .B2(_01866_),
    .C1(_01871_),
    .X(_01872_));
 sky130_fd_sc_hd__inv_2 _21864_ (.A(net5375),
    .Y(_01873_));
 sky130_fd_sc_hd__o32a_1 _21865_ (.A1(net3780),
    .A2(net3788),
    .A3(_01865_),
    .B1(_01872_),
    .B2(net3776),
    .X(_01874_));
 sky130_fd_sc_hd__xor2_1 _21866_ (.A(_01862_),
    .B(net1718),
    .X(_01875_));
 sky130_fd_sc_hd__xnor2_2 _21867_ (.A(_01860_),
    .B(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__xnor2_1 _21868_ (.A(net1171),
    .B(_01876_),
    .Y(_01877_));
 sky130_fd_sc_hd__xnor2_2 _21869_ (.A(net1047),
    .B(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__and2_1 _21870_ (.A(net1048),
    .B(net1172),
    .X(_01879_));
 sky130_fd_sc_hd__or2_1 _21871_ (.A(net2066),
    .B(_01792_),
    .X(_01880_));
 sky130_fd_sc_hd__nand2_1 _21872_ (.A(net2066),
    .B(_01792_),
    .Y(_01881_));
 sky130_fd_sc_hd__and2_1 _21873_ (.A(_01880_),
    .B(_01881_),
    .X(_01882_));
 sky130_fd_sc_hd__nor2_1 _21874_ (.A(net1048),
    .B(net1172),
    .Y(_01883_));
 sky130_fd_sc_hd__o21ba_1 _21875_ (.A1(_01879_),
    .A2(_01882_),
    .B1_N(_01883_),
    .X(_01884_));
 sky130_fd_sc_hd__xnor2_1 _21876_ (.A(_01878_),
    .B(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__or2_1 _21877_ (.A(net2066),
    .B(_01788_),
    .X(_01886_));
 sky130_fd_sc_hd__buf_1 _21878_ (.A(net2064),
    .X(_01887_));
 sky130_fd_sc_hd__nand2_1 _21879_ (.A(_01887_),
    .B(_01788_),
    .Y(_01888_));
 sky130_fd_sc_hd__a22o_1 _21880_ (.A1(_01780_),
    .A2(_01790_),
    .B1(_01886_),
    .B2(_01888_),
    .X(_01889_));
 sky130_fd_sc_hd__o21a_1 _21881_ (.A1(_01780_),
    .A2(_01790_),
    .B1(_01889_),
    .X(_01890_));
 sky130_fd_sc_hd__xnor2_1 _21882_ (.A(_01799_),
    .B(net1046),
    .Y(_01891_));
 sky130_fd_sc_hd__xnor2_1 _21883_ (.A(_01885_),
    .B(_01891_),
    .Y(_01892_));
 sky130_fd_sc_hd__inv_2 _21884_ (.A(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hd__buf_1 _21885_ (.A(net2477),
    .X(_01894_));
 sky130_fd_sc_hd__xnor2_1 _21886_ (.A(net2068),
    .B(_01794_),
    .Y(_01895_));
 sky130_fd_sc_hd__and2_1 _21887_ (.A(_01795_),
    .B(_01895_),
    .X(_01896_));
 sky130_fd_sc_hd__nor2_1 _21888_ (.A(_01795_),
    .B(_01895_),
    .Y(_01897_));
 sky130_fd_sc_hd__nor2_1 _21889_ (.A(_01744_),
    .B(_01897_),
    .Y(_01898_));
 sky130_fd_sc_hd__or2_1 _21890_ (.A(_01896_),
    .B(_01898_),
    .X(_01899_));
 sky130_fd_sc_hd__and2_1 _21891_ (.A(net2063),
    .B(_01897_),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_1 _21892_ (.A0(_01896_),
    .A1(_01900_),
    .S(_01744_),
    .X(_01901_));
 sky130_fd_sc_hd__a21oi_1 _21893_ (.A1(_01894_),
    .A2(_01899_),
    .B1(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__xnor2_1 _21894_ (.A(_01893_),
    .B(_01902_),
    .Y(_01903_));
 sky130_fd_sc_hd__a21bo_1 _21895_ (.A1(_01742_),
    .A2(_01802_),
    .B1_N(_01714_),
    .X(_01904_));
 sky130_fd_sc_hd__o21ai_2 _21896_ (.A1(_01742_),
    .A2(_01802_),
    .B1(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__xnor2_1 _21897_ (.A(net599),
    .B(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hd__xnor2_1 _21898_ (.A(_01827_),
    .B(_01906_),
    .Y(_01907_));
 sky130_fd_sc_hd__inv_2 _21899_ (.A(net5968),
    .Y(_01908_));
 sky130_fd_sc_hd__o21ba_1 _21900_ (.A1(_01908_),
    .A2(_01812_),
    .B1_N(\pid_d.prev_error[6] ),
    .X(_01909_));
 sky130_fd_sc_hd__a21o_1 _21901_ (.A1(_01908_),
    .A2(_01812_),
    .B1(_01909_),
    .X(_01910_));
 sky130_fd_sc_hd__xnor2_1 _21902_ (.A(\pid_d.prev_error[7] ),
    .B(\pid_d.curr_error[7] ),
    .Y(_01911_));
 sky130_fd_sc_hd__nand2_1 _21903_ (.A(_01910_),
    .B(_01911_),
    .Y(_01912_));
 sky130_fd_sc_hd__or2_1 _21904_ (.A(_01910_),
    .B(_01911_),
    .X(_01913_));
 sky130_fd_sc_hd__and3_1 _21905_ (.A(net4352),
    .B(_01912_),
    .C(_01913_),
    .X(_01914_));
 sky130_fd_sc_hd__a221o_1 _21906_ (.A1(net4385),
    .A2(net803),
    .B1(net413),
    .B2(net4319),
    .C1(net699),
    .X(_01915_));
 sky130_fd_sc_hd__a22o_1 _21907_ (.A1(net9022),
    .A2(net3123),
    .B1(net2078),
    .B2(_01915_),
    .X(_00526_));
 sky130_fd_sc_hd__inv_2 _21908_ (.A(\pid_d.prev_int[7] ),
    .Y(_01916_));
 sky130_fd_sc_hd__inv_2 _21909_ (.A(net5978),
    .Y(_01917_));
 sky130_fd_sc_hd__o21a_1 _21910_ (.A1(_01916_),
    .A2(_01821_),
    .B1(_01917_),
    .X(_01918_));
 sky130_fd_sc_hd__a21o_1 _21911_ (.A1(_01916_),
    .A2(_01821_),
    .B1(_01918_),
    .X(_01919_));
 sky130_fd_sc_hd__xor2_1 _21912_ (.A(net5977),
    .B(\pid_d.prev_int[8] ),
    .X(_01920_));
 sky130_fd_sc_hd__xnor2_1 _21913_ (.A(_01919_),
    .B(_01920_),
    .Y(_01921_));
 sky130_fd_sc_hd__inv_2 _21914_ (.A(_01905_),
    .Y(_01922_));
 sky130_fd_sc_hd__nand2_1 _21915_ (.A(net599),
    .B(_01922_),
    .Y(_01923_));
 sky130_fd_sc_hd__nor2_1 _21916_ (.A(net599),
    .B(_01922_),
    .Y(_01924_));
 sky130_fd_sc_hd__a31o_1 _21917_ (.A1(_01825_),
    .A2(_01826_),
    .A3(_01923_),
    .B1(_01924_),
    .X(_01925_));
 sky130_fd_sc_hd__o21a_1 _21918_ (.A1(_01832_),
    .A2(_01834_),
    .B1(_01833_),
    .X(_01926_));
 sky130_fd_sc_hd__a21oi_1 _21919_ (.A1(_01832_),
    .A2(_01834_),
    .B1(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__nand2_1 _21920_ (.A(_00977_),
    .B(net5649),
    .Y(_01928_));
 sky130_fd_sc_hd__nand2_1 _21921_ (.A(net5693),
    .B(net5514),
    .Y(_01929_));
 sky130_fd_sc_hd__nand2_1 _21922_ (.A(net5540),
    .B(net5669),
    .Y(_01930_));
 sky130_fd_sc_hd__xnor2_1 _21923_ (.A(_01929_),
    .B(_01930_),
    .Y(_01931_));
 sky130_fd_sc_hd__xnor2_1 _21924_ (.A(_01928_),
    .B(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__nand2_2 _21925_ (.A(net5719),
    .B(net5479),
    .Y(_01933_));
 sky130_fd_sc_hd__nand2_1 _21926_ (.A(net5710),
    .B(net5499),
    .Y(_01934_));
 sky130_fd_sc_hd__nand2_1 _21927_ (.A(net5750),
    .B(net5463),
    .Y(_01935_));
 sky130_fd_sc_hd__xnor2_1 _21928_ (.A(_01934_),
    .B(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__xnor2_2 _21929_ (.A(_01933_),
    .B(_01936_),
    .Y(_01937_));
 sky130_fd_sc_hd__xor2_1 _21930_ (.A(_01932_),
    .B(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__xnor2_1 _21931_ (.A(_01927_),
    .B(_01938_),
    .Y(_01939_));
 sky130_fd_sc_hd__o21ba_1 _21932_ (.A1(_01836_),
    .A2(_01841_),
    .B1_N(_01831_),
    .X(_01940_));
 sky130_fd_sc_hd__a21o_1 _21933_ (.A1(_01836_),
    .A2(_01841_),
    .B1(_01940_),
    .X(_01941_));
 sky130_fd_sc_hd__nand2_2 _21934_ (.A(net5799),
    .B(net5393),
    .Y(_01942_));
 sky130_fd_sc_hd__nand2_1 _21935_ (.A(net5784),
    .B(net5408),
    .Y(_01943_));
 sky130_fd_sc_hd__nand2_1 _21936_ (.A(net5763),
    .B(net5432),
    .Y(_01944_));
 sky130_fd_sc_hd__xnor2_1 _21937_ (.A(_01943_),
    .B(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__xnor2_2 _21938_ (.A(_01942_),
    .B(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hd__o21a_1 _21939_ (.A1(_01837_),
    .A2(_01839_),
    .B1(_01838_),
    .X(_01947_));
 sky130_fd_sc_hd__a21oi_2 _21940_ (.A1(_01837_),
    .A2(_01839_),
    .B1(_01947_),
    .Y(_01948_));
 sky130_fd_sc_hd__o21ba_1 _21941_ (.A1(_01847_),
    .A2(_01848_),
    .B1_N(_01846_),
    .X(_01949_));
 sky130_fd_sc_hd__a21oi_2 _21942_ (.A1(_01847_),
    .A2(_01848_),
    .B1(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__xnor2_1 _21943_ (.A(_01948_),
    .B(_01950_),
    .Y(_01951_));
 sky130_fd_sc_hd__xnor2_2 _21944_ (.A(_01946_),
    .B(_01951_),
    .Y(_01952_));
 sky130_fd_sc_hd__xor2_1 _21945_ (.A(_01941_),
    .B(_01952_),
    .X(_01953_));
 sky130_fd_sc_hd__xnor2_1 _21946_ (.A(net1714),
    .B(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__or3b_1 _21947_ (.A(net5839),
    .B(net5394),
    .C_N(net5406),
    .X(_01955_));
 sky130_fd_sc_hd__a21oi_1 _21948_ (.A1(_01783_),
    .A2(_01955_),
    .B1(_01781_),
    .Y(_01956_));
 sky130_fd_sc_hd__a41o_1 _21949_ (.A1(net5839),
    .A2(net5420),
    .A3(net5395),
    .A4(net3776),
    .B1(_01956_),
    .X(_01957_));
 sky130_fd_sc_hd__nor2_1 _21950_ (.A(net2064),
    .B(net1718),
    .Y(_01958_));
 sky130_fd_sc_hd__a21oi_2 _21951_ (.A1(net5812),
    .A2(_01957_),
    .B1(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__a21bo_1 _21952_ (.A1(net2474),
    .A2(_01854_),
    .B1_N(_01850_),
    .X(_01960_));
 sky130_fd_sc_hd__o21ai_1 _21953_ (.A1(net2474),
    .A2(_01854_),
    .B1(_01960_),
    .Y(_01961_));
 sky130_fd_sc_hd__o21a_1 _21954_ (.A1(net5858),
    .A2(net3787),
    .B1(net5841),
    .X(_01962_));
 sky130_fd_sc_hd__a21o_1 _21955_ (.A1(net5858),
    .A2(net3787),
    .B1(_01962_),
    .X(_01963_));
 sky130_fd_sc_hd__nor2_1 _21956_ (.A(net5841),
    .B(net5862),
    .Y(_01964_));
 sky130_fd_sc_hd__nand2_1 _21957_ (.A(net3780),
    .B(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__nand2_1 _21958_ (.A(net5380),
    .B(_01965_),
    .Y(_01966_));
 sky130_fd_sc_hd__a21o_1 _21959_ (.A1(net5817),
    .A2(_01963_),
    .B1(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__xnor2_1 _21960_ (.A(net1713),
    .B(_01967_),
    .Y(_01968_));
 sky130_fd_sc_hd__xnor2_2 _21961_ (.A(_01959_),
    .B(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__a21bo_1 _21962_ (.A1(_01845_),
    .A2(_01856_),
    .B1_N(net1719),
    .X(_01970_));
 sky130_fd_sc_hd__o21a_1 _21963_ (.A1(_01845_),
    .A2(_01856_),
    .B1(_01970_),
    .X(_01971_));
 sky130_fd_sc_hd__xor2_2 _21964_ (.A(_01969_),
    .B(net1170),
    .X(_01972_));
 sky130_fd_sc_hd__xnor2_4 _21965_ (.A(net1045),
    .B(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__and2_1 _21966_ (.A(net1047),
    .B(net1171),
    .X(_01974_));
 sky130_fd_sc_hd__or2_1 _21967_ (.A(net2065),
    .B(_01876_),
    .X(_01975_));
 sky130_fd_sc_hd__nand2_1 _21968_ (.A(net2065),
    .B(_01876_),
    .Y(_01976_));
 sky130_fd_sc_hd__and2_1 _21969_ (.A(_01975_),
    .B(_01976_),
    .X(_01977_));
 sky130_fd_sc_hd__or2_1 _21970_ (.A(net1047),
    .B(net1171),
    .X(_01978_));
 sky130_fd_sc_hd__o21ai_1 _21971_ (.A1(_01974_),
    .A2(_01977_),
    .B1(_01978_),
    .Y(_01979_));
 sky130_fd_sc_hd__xnor2_2 _21972_ (.A(_01973_),
    .B(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__and2_1 _21973_ (.A(net1716),
    .B(net1718),
    .X(_01981_));
 sky130_fd_sc_hd__a211o_1 _21974_ (.A1(_01860_),
    .A2(_01862_),
    .B1(_01958_),
    .C1(_01981_),
    .X(_01982_));
 sky130_fd_sc_hd__o21a_1 _21975_ (.A1(_01860_),
    .A2(_01862_),
    .B1(_01982_),
    .X(_01983_));
 sky130_fd_sc_hd__xor2_1 _21976_ (.A(_01799_),
    .B(net1044),
    .X(_01984_));
 sky130_fd_sc_hd__xnor2_1 _21977_ (.A(_01980_),
    .B(_01984_),
    .Y(_01985_));
 sky130_fd_sc_hd__inv_2 _21978_ (.A(_01985_),
    .Y(_01986_));
 sky130_fd_sc_hd__mux2_1 _21979_ (.A0(_01880_),
    .A1(_01881_),
    .S(_01878_),
    .X(_01987_));
 sky130_fd_sc_hd__xnor2_1 _21980_ (.A(net1717),
    .B(_01878_),
    .Y(_01988_));
 sky130_fd_sc_hd__a2bb2o_1 _21981_ (.A1_N(_01879_),
    .A2_N(_01987_),
    .B1(_01988_),
    .B2(_01883_),
    .X(_01989_));
 sky130_fd_sc_hd__nor2_1 _21982_ (.A(net2477),
    .B(net1046),
    .Y(_01990_));
 sky130_fd_sc_hd__and2_1 _21983_ (.A(_01989_),
    .B(_01990_),
    .X(_01991_));
 sky130_fd_sc_hd__or2_1 _21984_ (.A(net2068),
    .B(_01885_),
    .X(_01992_));
 sky130_fd_sc_hd__nand2_1 _21985_ (.A(net2068),
    .B(_01885_),
    .Y(_01993_));
 sky130_fd_sc_hd__a21oi_1 _21986_ (.A1(_01992_),
    .A2(_01993_),
    .B1(_01990_),
    .Y(_01994_));
 sky130_fd_sc_hd__a21oi_1 _21987_ (.A1(net2477),
    .A2(net1046),
    .B1(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__or2_1 _21988_ (.A(_01989_),
    .B(_01995_),
    .X(_01996_));
 sky130_fd_sc_hd__and2b_1 _21989_ (.A_N(_01991_),
    .B(_01996_),
    .X(_01997_));
 sky130_fd_sc_hd__xnor2_1 _21990_ (.A(_01986_),
    .B(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__or2_1 _21991_ (.A(_01892_),
    .B(_01899_),
    .X(_01999_));
 sky130_fd_sc_hd__o21ai_1 _21992_ (.A1(_01893_),
    .A2(_01897_),
    .B1(_01744_),
    .Y(_02000_));
 sky130_fd_sc_hd__or2_1 _21993_ (.A(_01892_),
    .B(_01896_),
    .X(_02001_));
 sky130_fd_sc_hd__a21o_1 _21994_ (.A1(_02000_),
    .A2(_02001_),
    .B1(_01894_),
    .X(_02002_));
 sky130_fd_sc_hd__nand3_1 _21995_ (.A(_01998_),
    .B(_01999_),
    .C(_02002_),
    .Y(_02003_));
 sky130_fd_sc_hd__a21oi_2 _21996_ (.A1(_01999_),
    .A2(_02002_),
    .B1(_01998_),
    .Y(_02004_));
 sky130_fd_sc_hd__inv_2 _21997_ (.A(_02004_),
    .Y(_02005_));
 sky130_fd_sc_hd__nand2_1 _21998_ (.A(_02003_),
    .B(_02005_),
    .Y(_02006_));
 sky130_fd_sc_hd__xnor2_1 _21999_ (.A(net471),
    .B(_02006_),
    .Y(_02007_));
 sky130_fd_sc_hd__inv_2 _22000_ (.A(\pid_d.curr_error[7] ),
    .Y(_02008_));
 sky130_fd_sc_hd__o21ba_1 _22001_ (.A1(_02008_),
    .A2(_01910_),
    .B1_N(\pid_d.prev_error[7] ),
    .X(_02009_));
 sky130_fd_sc_hd__a21o_1 _22002_ (.A1(_02008_),
    .A2(_01910_),
    .B1(_02009_),
    .X(_02010_));
 sky130_fd_sc_hd__xnor2_1 _22003_ (.A(\pid_d.prev_error[8] ),
    .B(\pid_d.curr_error[8] ),
    .Y(_02011_));
 sky130_fd_sc_hd__nand2_1 _22004_ (.A(_02010_),
    .B(_02011_),
    .Y(_02012_));
 sky130_fd_sc_hd__or2_1 _22005_ (.A(_02010_),
    .B(_02011_),
    .X(_02013_));
 sky130_fd_sc_hd__and3_1 _22006_ (.A(net4353),
    .B(_02012_),
    .C(_02013_),
    .X(_02014_));
 sky130_fd_sc_hd__a221o_1 _22007_ (.A1(net4383),
    .A2(net698),
    .B1(net347),
    .B2(net4319),
    .C1(_02014_),
    .X(_02015_));
 sky130_fd_sc_hd__a22o_1 _22008_ (.A1(net9035),
    .A2(net3123),
    .B1(net2078),
    .B2(_02015_),
    .X(_00527_));
 sky130_fd_sc_hd__inv_2 _22009_ (.A(\pid_d.prev_int[8] ),
    .Y(_02016_));
 sky130_fd_sc_hd__inv_2 _22010_ (.A(net5977),
    .Y(_02017_));
 sky130_fd_sc_hd__a21o_1 _22011_ (.A1(_02016_),
    .A2(_01919_),
    .B1(_02017_),
    .X(_02018_));
 sky130_fd_sc_hd__o21a_1 _22012_ (.A1(_02016_),
    .A2(_01919_),
    .B1(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__xor2_1 _22013_ (.A(net5976),
    .B(\pid_d.prev_int[9] ),
    .X(_02020_));
 sky130_fd_sc_hd__xnor2_1 _22014_ (.A(_02019_),
    .B(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__a21oi_1 _22015_ (.A1(net471),
    .A2(_02003_),
    .B1(_02004_),
    .Y(_02022_));
 sky130_fd_sc_hd__o21a_1 _22016_ (.A1(_01928_),
    .A2(_01930_),
    .B1(_01929_),
    .X(_02023_));
 sky130_fd_sc_hd__a21oi_2 _22017_ (.A1(_01928_),
    .A2(_01930_),
    .B1(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__nand2b_1 _22018_ (.A_N(net5540),
    .B(net5649),
    .Y(_02025_));
 sky130_fd_sc_hd__nand2_1 _22019_ (.A(net5693),
    .B(net5498),
    .Y(_02026_));
 sky130_fd_sc_hd__nand2_1 _22020_ (.A(net5513),
    .B(net5669),
    .Y(_02027_));
 sky130_fd_sc_hd__xnor2_1 _22021_ (.A(_02026_),
    .B(_02027_),
    .Y(_02028_));
 sky130_fd_sc_hd__xnor2_1 _22022_ (.A(_02025_),
    .B(_02028_),
    .Y(_02029_));
 sky130_fd_sc_hd__nand2_1 _22023_ (.A(net5709),
    .B(net5480),
    .Y(_02030_));
 sky130_fd_sc_hd__nand2_1 _22024_ (.A(net5746),
    .B(net5433),
    .Y(_02031_));
 sky130_fd_sc_hd__nand2_1 _22025_ (.A(net5721),
    .B(net5464),
    .Y(_02032_));
 sky130_fd_sc_hd__xor2_1 _22026_ (.A(_02031_),
    .B(_02032_),
    .X(_02033_));
 sky130_fd_sc_hd__xnor2_2 _22027_ (.A(_02030_),
    .B(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__xnor2_1 _22028_ (.A(_02029_),
    .B(_02034_),
    .Y(_02035_));
 sky130_fd_sc_hd__xnor2_1 _22029_ (.A(_02024_),
    .B(_02035_),
    .Y(_02036_));
 sky130_fd_sc_hd__o21ba_1 _22030_ (.A1(_01932_),
    .A2(_01937_),
    .B1_N(_01927_),
    .X(_02037_));
 sky130_fd_sc_hd__a21o_1 _22031_ (.A1(_01932_),
    .A2(_01937_),
    .B1(_02037_),
    .X(_02038_));
 sky130_fd_sc_hd__nand2_2 _22032_ (.A(net5799),
    .B(net5375),
    .Y(_02039_));
 sky130_fd_sc_hd__nand2_1 _22033_ (.A(net5763),
    .B(net5410),
    .Y(_02040_));
 sky130_fd_sc_hd__nand2_1 _22034_ (.A(net5779),
    .B(net5389),
    .Y(_02041_));
 sky130_fd_sc_hd__xnor2_1 _22035_ (.A(_02040_),
    .B(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__xnor2_2 _22036_ (.A(_02039_),
    .B(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__o21a_1 _22037_ (.A1(_01933_),
    .A2(_01935_),
    .B1(_01934_),
    .X(_02044_));
 sky130_fd_sc_hd__a21oi_2 _22038_ (.A1(_01933_),
    .A2(_01935_),
    .B1(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__o21a_1 _22039_ (.A1(_01942_),
    .A2(_01943_),
    .B1(_01944_),
    .X(_02046_));
 sky130_fd_sc_hd__a21oi_2 _22040_ (.A1(_01942_),
    .A2(_01943_),
    .B1(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__xnor2_1 _22041_ (.A(_02045_),
    .B(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__xnor2_2 _22042_ (.A(_02043_),
    .B(_02048_),
    .Y(_02049_));
 sky130_fd_sc_hd__xnor2_1 _22043_ (.A(_02038_),
    .B(_02049_),
    .Y(_02050_));
 sky130_fd_sc_hd__xnor2_1 _22044_ (.A(_02036_),
    .B(_02050_),
    .Y(_02051_));
 sky130_fd_sc_hd__o21a_1 _22045_ (.A1(_01941_),
    .A2(_01952_),
    .B1(net1714),
    .X(_02052_));
 sky130_fd_sc_hd__a21oi_1 _22046_ (.A1(_01941_),
    .A2(_01952_),
    .B1(_02052_),
    .Y(_02053_));
 sky130_fd_sc_hd__or3_1 _22047_ (.A(net3780),
    .B(net5395),
    .C(_01964_),
    .X(_02054_));
 sky130_fd_sc_hd__and3_1 _22048_ (.A(net5817),
    .B(net5841),
    .C(net5858),
    .X(_02055_));
 sky130_fd_sc_hd__a31o_1 _22049_ (.A1(net2067),
    .A2(_01965_),
    .A3(_02054_),
    .B1(_02055_),
    .X(_02056_));
 sky130_fd_sc_hd__nand2_1 _22050_ (.A(net5380),
    .B(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__nor2_1 _22051_ (.A(_01966_),
    .B(_02055_),
    .Y(_02058_));
 sky130_fd_sc_hd__xnor2_2 _22052_ (.A(net2067),
    .B(_02058_),
    .Y(_02059_));
 sky130_fd_sc_hd__and2_1 _22053_ (.A(_02057_),
    .B(_02059_),
    .X(_02060_));
 sky130_fd_sc_hd__nor2_1 _22054_ (.A(_02057_),
    .B(_02059_),
    .Y(_02061_));
 sky130_fd_sc_hd__a21bo_1 _22055_ (.A1(_01948_),
    .A2(_01950_),
    .B1_N(_01946_),
    .X(_02062_));
 sky130_fd_sc_hd__o21ai_1 _22056_ (.A1(_01948_),
    .A2(_01950_),
    .B1(_02062_),
    .Y(_02063_));
 sky130_fd_sc_hd__o21ai_1 _22057_ (.A1(_02060_),
    .A2(_02061_),
    .B1(net1710),
    .Y(_02064_));
 sky130_fd_sc_hd__or3_1 _22058_ (.A(net1710),
    .B(_02060_),
    .C(_02061_),
    .X(_02065_));
 sky130_fd_sc_hd__and2_1 _22059_ (.A(_02064_),
    .B(_02065_),
    .X(_02066_));
 sky130_fd_sc_hd__nor2_1 _22060_ (.A(net1038),
    .B(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__nand2_1 _22061_ (.A(net1038),
    .B(_02066_),
    .Y(_02068_));
 sky130_fd_sc_hd__or2b_1 _22062_ (.A(_02067_),
    .B_N(_02068_),
    .X(_02069_));
 sky130_fd_sc_hd__xnor2_1 _22063_ (.A(net1041),
    .B(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__nand2_1 _22064_ (.A(net1715),
    .B(_01969_),
    .Y(_02071_));
 sky130_fd_sc_hd__or2_1 _22065_ (.A(net1715),
    .B(_01969_),
    .X(_02072_));
 sky130_fd_sc_hd__o211a_1 _22066_ (.A1(net1045),
    .A2(net1170),
    .B1(_02071_),
    .C1(_02072_),
    .X(_02073_));
 sky130_fd_sc_hd__a21oi_1 _22067_ (.A1(net1045),
    .A2(net1170),
    .B1(_02073_),
    .Y(_02074_));
 sky130_fd_sc_hd__nor2_1 _22068_ (.A(net1716),
    .B(_01967_),
    .Y(_02075_));
 sky130_fd_sc_hd__and2_1 _22069_ (.A(net1716),
    .B(_01967_),
    .X(_02076_));
 sky130_fd_sc_hd__o22a_1 _22070_ (.A1(_01959_),
    .A2(net1713),
    .B1(_02075_),
    .B2(_02076_),
    .X(_02077_));
 sky130_fd_sc_hd__a21oi_1 _22071_ (.A1(_01959_),
    .A2(net1713),
    .B1(_02077_),
    .Y(_02078_));
 sky130_fd_sc_hd__xnor2_2 _22072_ (.A(net2062),
    .B(net945),
    .Y(_02079_));
 sky130_fd_sc_hd__xnor2_1 _22073_ (.A(net802),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__xnor2_1 _22074_ (.A(_02070_),
    .B(_02080_),
    .Y(_02081_));
 sky130_fd_sc_hd__mux2_1 _22075_ (.A0(_01975_),
    .A1(_01976_),
    .S(_01973_),
    .X(_02082_));
 sky130_fd_sc_hd__xnor2_1 _22076_ (.A(net2067),
    .B(_01973_),
    .Y(_02083_));
 sky130_fd_sc_hd__o22ai_2 _22077_ (.A1(_01974_),
    .A2(_02082_),
    .B1(_02083_),
    .B2(_01978_),
    .Y(_02084_));
 sky130_fd_sc_hd__or2_1 _22078_ (.A(net1717),
    .B(_01980_),
    .X(_02085_));
 sky130_fd_sc_hd__nand2_1 _22079_ (.A(net1717),
    .B(_01980_),
    .Y(_02086_));
 sky130_fd_sc_hd__nor2_1 _22080_ (.A(net2477),
    .B(net1044),
    .Y(_02087_));
 sky130_fd_sc_hd__a21oi_1 _22081_ (.A1(_02085_),
    .A2(_02086_),
    .B1(_02087_),
    .Y(_02088_));
 sky130_fd_sc_hd__a21oi_1 _22082_ (.A1(net2059),
    .A2(net1044),
    .B1(_02088_),
    .Y(_02089_));
 sky130_fd_sc_hd__nor2_1 _22083_ (.A(_02084_),
    .B(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__nand2_1 _22084_ (.A(_02084_),
    .B(_02087_),
    .Y(_02091_));
 sky130_fd_sc_hd__and2b_1 _22085_ (.A_N(_02090_),
    .B(_02091_),
    .X(_02092_));
 sky130_fd_sc_hd__xnor2_1 _22086_ (.A(_02081_),
    .B(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__a21o_1 _22087_ (.A1(_01986_),
    .A2(_01996_),
    .B1(_01991_),
    .X(_02094_));
 sky130_fd_sc_hd__or2_1 _22088_ (.A(_02093_),
    .B(_02094_),
    .X(_02095_));
 sky130_fd_sc_hd__inv_2 _22089_ (.A(_02095_),
    .Y(_02096_));
 sky130_fd_sc_hd__and2_1 _22090_ (.A(_02093_),
    .B(_02094_),
    .X(_02097_));
 sky130_fd_sc_hd__nor2_1 _22091_ (.A(_02096_),
    .B(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__xnor2_1 _22092_ (.A(_02022_),
    .B(_02098_),
    .Y(_02099_));
 sky130_fd_sc_hd__inv_2 _22093_ (.A(\pid_d.curr_error[8] ),
    .Y(_02100_));
 sky130_fd_sc_hd__o21ba_1 _22094_ (.A1(_02100_),
    .A2(_02010_),
    .B1_N(\pid_d.prev_error[8] ),
    .X(_02101_));
 sky130_fd_sc_hd__a21o_1 _22095_ (.A1(_02100_),
    .A2(_02010_),
    .B1(_02101_),
    .X(_02102_));
 sky130_fd_sc_hd__xnor2_1 _22096_ (.A(\pid_d.prev_error[9] ),
    .B(net5967),
    .Y(_02103_));
 sky130_fd_sc_hd__nand2_1 _22097_ (.A(_02102_),
    .B(_02103_),
    .Y(_02104_));
 sky130_fd_sc_hd__or2_1 _22098_ (.A(_02102_),
    .B(_02103_),
    .X(_02105_));
 sky130_fd_sc_hd__and3_1 _22099_ (.A(net4353),
    .B(_02104_),
    .C(_02105_),
    .X(_02106_));
 sky130_fd_sc_hd__a221o_1 _22100_ (.A1(net4383),
    .A2(_02021_),
    .B1(net343),
    .B2(net4319),
    .C1(net522),
    .X(_02107_));
 sky130_fd_sc_hd__a22o_1 _22101_ (.A1(net9018),
    .A2(_12500_),
    .B1(_12503_),
    .B2(_02107_),
    .X(_00528_));
 sky130_fd_sc_hd__inv_2 _22102_ (.A(\pid_d.prev_int[9] ),
    .Y(_02108_));
 sky130_fd_sc_hd__inv_2 _22103_ (.A(net5976),
    .Y(_02109_));
 sky130_fd_sc_hd__o21a_1 _22104_ (.A1(_02108_),
    .A2(_02019_),
    .B1(_02109_),
    .X(_02110_));
 sky130_fd_sc_hd__a21o_1 _22105_ (.A1(_02108_),
    .A2(_02019_),
    .B1(_02110_),
    .X(_02111_));
 sky130_fd_sc_hd__xor2_1 _22106_ (.A(\pid_d.curr_int[10] ),
    .B(\pid_d.prev_int[10] ),
    .X(_02112_));
 sky130_fd_sc_hd__xnor2_1 _22107_ (.A(_02111_),
    .B(_02112_),
    .Y(_02113_));
 sky130_fd_sc_hd__a211o_1 _22108_ (.A1(net471),
    .A2(_02003_),
    .B1(_02004_),
    .C1(_02097_),
    .X(_02114_));
 sky130_fd_sc_hd__nand2_1 _22109_ (.A(_02095_),
    .B(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__o21ai_1 _22110_ (.A1(_02081_),
    .A2(_02090_),
    .B1(_02091_),
    .Y(_02116_));
 sky130_fd_sc_hd__a21o_1 _22111_ (.A1(net802),
    .A2(_02079_),
    .B1(_02070_),
    .X(_02117_));
 sky130_fd_sc_hd__o21ai_2 _22112_ (.A1(net802),
    .A2(_02079_),
    .B1(_02117_),
    .Y(_02118_));
 sky130_fd_sc_hd__and2_1 _22113_ (.A(net2062),
    .B(net945),
    .X(_02119_));
 sky130_fd_sc_hd__a21bo_1 _22114_ (.A1(_02024_),
    .A2(_02034_),
    .B1_N(_02029_),
    .X(_02120_));
 sky130_fd_sc_hd__o21a_1 _22115_ (.A1(_02024_),
    .A2(_02034_),
    .B1(_02120_),
    .X(_02121_));
 sky130_fd_sc_hd__nand2_1 _22116_ (.A(_00917_),
    .B(net5661),
    .Y(_02122_));
 sky130_fd_sc_hd__nand2_1 _22117_ (.A(net5692),
    .B(net5481),
    .Y(_02123_));
 sky130_fd_sc_hd__nand2_1 _22118_ (.A(net5497),
    .B(net5672),
    .Y(_02124_));
 sky130_fd_sc_hd__xnor2_1 _22119_ (.A(_02123_),
    .B(_02124_),
    .Y(_02125_));
 sky130_fd_sc_hd__xnor2_1 _22120_ (.A(_02122_),
    .B(_02125_),
    .Y(_02126_));
 sky130_fd_sc_hd__o21a_1 _22121_ (.A1(_02025_),
    .A2(_02027_),
    .B1(_02026_),
    .X(_02127_));
 sky130_fd_sc_hd__a21oi_2 _22122_ (.A1(_02025_),
    .A2(_02027_),
    .B1(_02127_),
    .Y(_02128_));
 sky130_fd_sc_hd__nand2_1 _22123_ (.A(net5708),
    .B(net5464),
    .Y(_02129_));
 sky130_fd_sc_hd__nand2_1 _22124_ (.A(net5745),
    .B(net5411),
    .Y(_02130_));
 sky130_fd_sc_hd__nand2_1 _22125_ (.A(net5720),
    .B(net5437),
    .Y(_02131_));
 sky130_fd_sc_hd__xor2_1 _22126_ (.A(_02130_),
    .B(_02131_),
    .X(_02132_));
 sky130_fd_sc_hd__xnor2_2 _22127_ (.A(_02129_),
    .B(_02132_),
    .Y(_02133_));
 sky130_fd_sc_hd__xnor2_1 _22128_ (.A(_02128_),
    .B(_02133_),
    .Y(_02134_));
 sky130_fd_sc_hd__xnor2_1 _22129_ (.A(_02126_),
    .B(_02134_),
    .Y(_02135_));
 sky130_fd_sc_hd__xnor2_1 _22130_ (.A(net5779),
    .B(net5799),
    .Y(_02136_));
 sky130_fd_sc_hd__o211a_1 _22131_ (.A1(net3779),
    .A2(_02136_),
    .B1(net5764),
    .C1(net5389),
    .X(_02137_));
 sky130_fd_sc_hd__a211o_1 _22132_ (.A1(net5764),
    .A2(net5389),
    .B1(net3779),
    .C1(_02136_),
    .X(_02138_));
 sky130_fd_sc_hd__or2b_1 _22133_ (.A(_02137_),
    .B_N(_02138_),
    .X(_02139_));
 sky130_fd_sc_hd__o21ai_1 _22134_ (.A1(_02031_),
    .A2(_02032_),
    .B1(_02030_),
    .Y(_02140_));
 sky130_fd_sc_hd__a21bo_1 _22135_ (.A1(_02031_),
    .A2(_02032_),
    .B1_N(_02140_),
    .X(_02141_));
 sky130_fd_sc_hd__o21a_1 _22136_ (.A1(_02039_),
    .A2(_02041_),
    .B1(_02040_),
    .X(_02142_));
 sky130_fd_sc_hd__a21o_1 _22137_ (.A1(_02039_),
    .A2(_02041_),
    .B1(_02142_),
    .X(_02143_));
 sky130_fd_sc_hd__xnor2_1 _22138_ (.A(_02141_),
    .B(_02143_),
    .Y(_02144_));
 sky130_fd_sc_hd__xnor2_2 _22139_ (.A(_02139_),
    .B(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__xnor2_1 _22140_ (.A(_02135_),
    .B(_02145_),
    .Y(_02146_));
 sky130_fd_sc_hd__xnor2_1 _22141_ (.A(net1389),
    .B(_02146_),
    .Y(_02147_));
 sky130_fd_sc_hd__o21a_1 _22142_ (.A1(_02038_),
    .A2(_02049_),
    .B1(_02036_),
    .X(_02148_));
 sky130_fd_sc_hd__a21oi_1 _22143_ (.A1(_02038_),
    .A2(_02049_),
    .B1(_02148_),
    .Y(_02149_));
 sky130_fd_sc_hd__a21o_1 _22144_ (.A1(net5841),
    .A2(net5858),
    .B1(net2067),
    .X(_02150_));
 sky130_fd_sc_hd__a2bb2o_1 _22145_ (.A1_N(net2065),
    .A2_N(_01964_),
    .B1(_02150_),
    .B2(net5817),
    .X(_02151_));
 sky130_fd_sc_hd__nand2_2 _22146_ (.A(net5380),
    .B(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__a21bo_1 _22147_ (.A1(_02045_),
    .A2(_02047_),
    .B1_N(_02043_),
    .X(_02153_));
 sky130_fd_sc_hd__o21a_1 _22148_ (.A1(_02045_),
    .A2(_02047_),
    .B1(_02153_),
    .X(_02154_));
 sky130_fd_sc_hd__inv_2 _22149_ (.A(net1708),
    .Y(_02155_));
 sky130_fd_sc_hd__xnor2_1 _22150_ (.A(_02152_),
    .B(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hd__xnor2_1 _22151_ (.A(net1036),
    .B(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__xnor2_1 _22152_ (.A(net1168),
    .B(_02157_),
    .Y(_02158_));
 sky130_fd_sc_hd__a21oi_4 _22153_ (.A1(net1041),
    .A2(_02068_),
    .B1(_02067_),
    .Y(_02159_));
 sky130_fd_sc_hd__nor2_1 _22154_ (.A(net1710),
    .B(_02057_),
    .Y(_02160_));
 sky130_fd_sc_hd__and2_1 _22155_ (.A(net1710),
    .B(_02057_),
    .X(_02161_));
 sky130_fd_sc_hd__inv_2 _22156_ (.A(_02059_),
    .Y(_02162_));
 sky130_fd_sc_hd__mux2_1 _22157_ (.A0(_02160_),
    .A1(_02161_),
    .S(_02162_),
    .X(_02163_));
 sky130_fd_sc_hd__xnor2_1 _22158_ (.A(net2476),
    .B(_02163_),
    .Y(_02164_));
 sky130_fd_sc_hd__xnor2_1 _22159_ (.A(_02159_),
    .B(_02164_),
    .Y(_02165_));
 sky130_fd_sc_hd__xnor2_2 _22160_ (.A(net859),
    .B(_02165_),
    .Y(_02166_));
 sky130_fd_sc_hd__xnor2_1 _22161_ (.A(_02119_),
    .B(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__xnor2_1 _22162_ (.A(_02118_),
    .B(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__nand2_1 _22163_ (.A(_02116_),
    .B(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__or2_1 _22164_ (.A(_02116_),
    .B(_02168_),
    .X(_02170_));
 sky130_fd_sc_hd__nand2_1 _22165_ (.A(_02169_),
    .B(_02170_),
    .Y(_02171_));
 sky130_fd_sc_hd__xnor2_1 _22166_ (.A(_02115_),
    .B(_02171_),
    .Y(_02172_));
 sky130_fd_sc_hd__inv_2 _22167_ (.A(net339),
    .Y(_02173_));
 sky130_fd_sc_hd__inv_2 _22168_ (.A(net5967),
    .Y(_02174_));
 sky130_fd_sc_hd__o21ba_1 _22169_ (.A1(_02174_),
    .A2(_02102_),
    .B1_N(\pid_d.prev_error[9] ),
    .X(_02175_));
 sky130_fd_sc_hd__a21o_1 _22170_ (.A1(_02174_),
    .A2(_02102_),
    .B1(_02175_),
    .X(_02176_));
 sky130_fd_sc_hd__xnor2_1 _22171_ (.A(\pid_d.prev_error[10] ),
    .B(\pid_d.curr_error[10] ),
    .Y(_02177_));
 sky130_fd_sc_hd__nand2_1 _22172_ (.A(_02176_),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__or2_1 _22173_ (.A(_02176_),
    .B(_02177_),
    .X(_02179_));
 sky130_fd_sc_hd__and3_1 _22174_ (.A(net4367),
    .B(_02178_),
    .C(_02179_),
    .X(_02180_));
 sky130_fd_sc_hd__a221o_1 _22175_ (.A1(net4381),
    .A2(_02113_),
    .B1(_02173_),
    .B2(net4314),
    .C1(net410),
    .X(_02181_));
 sky130_fd_sc_hd__a22o_1 _22176_ (.A1(\pid_d.curr_int[10] ),
    .A2(net3843),
    .B1(net2487),
    .B2(_02181_),
    .X(_00529_));
 sky130_fd_sc_hd__inv_2 _22177_ (.A(\pid_d.prev_int[10] ),
    .Y(_02182_));
 sky130_fd_sc_hd__inv_2 _22178_ (.A(\pid_d.curr_int[10] ),
    .Y(_02183_));
 sky130_fd_sc_hd__o21a_1 _22179_ (.A1(_02182_),
    .A2(_02111_),
    .B1(_02183_),
    .X(_02184_));
 sky130_fd_sc_hd__a21o_1 _22180_ (.A1(_02182_),
    .A2(_02111_),
    .B1(_02184_),
    .X(_02185_));
 sky130_fd_sc_hd__xor2_1 _22181_ (.A(\pid_d.curr_int[11] ),
    .B(\pid_d.prev_int[11] ),
    .X(_02186_));
 sky130_fd_sc_hd__xnor2_1 _22182_ (.A(_02185_),
    .B(_02186_),
    .Y(_02187_));
 sky130_fd_sc_hd__or2_1 _22183_ (.A(_02162_),
    .B(net859),
    .X(_02188_));
 sky130_fd_sc_hd__nand2_1 _22184_ (.A(_02159_),
    .B(_02188_),
    .Y(_02189_));
 sky130_fd_sc_hd__nor2_1 _22185_ (.A(_02059_),
    .B(_02161_),
    .Y(_02190_));
 sky130_fd_sc_hd__or2b_1 _22186_ (.A(net859),
    .B_N(_02159_),
    .X(_02191_));
 sky130_fd_sc_hd__a22o_1 _22187_ (.A1(_02160_),
    .A2(_02189_),
    .B1(_02190_),
    .B2(_02191_),
    .X(_02192_));
 sky130_fd_sc_hd__nand2_1 _22188_ (.A(net1710),
    .B(_02057_),
    .Y(_02193_));
 sky130_fd_sc_hd__a211o_1 _22189_ (.A1(_02159_),
    .A2(net859),
    .B1(_02160_),
    .C1(_02162_),
    .X(_02194_));
 sky130_fd_sc_hd__o21a_1 _22190_ (.A1(_02159_),
    .A2(_02193_),
    .B1(_02194_),
    .X(_02195_));
 sky130_fd_sc_hd__o21a_1 _22191_ (.A1(net2062),
    .A2(_02193_),
    .B1(_02159_),
    .X(_02196_));
 sky130_fd_sc_hd__or3b_1 _22192_ (.A(_02059_),
    .B(_02196_),
    .C_N(net859),
    .X(_02197_));
 sky130_fd_sc_hd__o221a_1 _22193_ (.A1(_02159_),
    .A2(_02188_),
    .B1(_02195_),
    .B2(net2062),
    .C1(_02197_),
    .X(_02198_));
 sky130_fd_sc_hd__a21bo_1 _22194_ (.A1(net2062),
    .A2(_02192_),
    .B1_N(_02198_),
    .X(_02199_));
 sky130_fd_sc_hd__a21o_1 _22195_ (.A1(net1712),
    .A2(_02152_),
    .B1(net1169),
    .X(_02200_));
 sky130_fd_sc_hd__buf_1 _22196_ (.A(_02200_),
    .X(_02201_));
 sky130_fd_sc_hd__xnor2_1 _22197_ (.A(net1708),
    .B(_02201_),
    .Y(_02202_));
 sky130_fd_sc_hd__a21bo_1 _22198_ (.A1(net1036),
    .A2(_02202_),
    .B1_N(net1168),
    .X(_02203_));
 sky130_fd_sc_hd__o21a_1 _22199_ (.A1(net1036),
    .A2(_02202_),
    .B1(_02203_),
    .X(_02204_));
 sky130_fd_sc_hd__o21ba_1 _22200_ (.A1(_02141_),
    .A2(_02143_),
    .B1_N(_02139_),
    .X(_02205_));
 sky130_fd_sc_hd__a21o_1 _22201_ (.A1(_02141_),
    .A2(_02143_),
    .B1(_02205_),
    .X(_02206_));
 sky130_fd_sc_hd__xor2_2 _22202_ (.A(net944),
    .B(net1706),
    .X(_02207_));
 sky130_fd_sc_hd__o21a_1 _22203_ (.A1(_02122_),
    .A2(_02124_),
    .B1(_02123_),
    .X(_02208_));
 sky130_fd_sc_hd__a21oi_1 _22204_ (.A1(_02122_),
    .A2(_02124_),
    .B1(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__nand2b_1 _22205_ (.A_N(\pid_d.mult0.a[9] ),
    .B(net5658),
    .Y(_02210_));
 sky130_fd_sc_hd__nand2_1 _22206_ (.A(net5489),
    .B(net5675),
    .Y(_02211_));
 sky130_fd_sc_hd__nand2_1 _22207_ (.A(net5690),
    .B(net5466),
    .Y(_02212_));
 sky130_fd_sc_hd__xnor2_1 _22208_ (.A(_02211_),
    .B(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__xnor2_1 _22209_ (.A(_02210_),
    .B(_02213_),
    .Y(_02214_));
 sky130_fd_sc_hd__nand2_2 _22210_ (.A(net5747),
    .B(net5404),
    .Y(_02215_));
 sky130_fd_sc_hd__nand2_1 _22211_ (.A(net5726),
    .B(net5409),
    .Y(_02216_));
 sky130_fd_sc_hd__nand2_1 _22212_ (.A(net5707),
    .B(net5430),
    .Y(_02217_));
 sky130_fd_sc_hd__xor2_1 _22213_ (.A(_02216_),
    .B(_02217_),
    .X(_02218_));
 sky130_fd_sc_hd__xnor2_2 _22214_ (.A(_02215_),
    .B(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__xnor2_1 _22215_ (.A(_02214_),
    .B(_02219_),
    .Y(_02220_));
 sky130_fd_sc_hd__xnor2_2 _22216_ (.A(net2052),
    .B(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__a21bo_1 _22217_ (.A1(_02128_),
    .A2(_02133_),
    .B1_N(_02126_),
    .X(_02222_));
 sky130_fd_sc_hd__o21a_1 _22218_ (.A1(_02128_),
    .A2(_02133_),
    .B1(_02222_),
    .X(_02223_));
 sky130_fd_sc_hd__o21ai_1 _22219_ (.A1(_02130_),
    .A2(_02131_),
    .B1(_02129_),
    .Y(_02224_));
 sky130_fd_sc_hd__a21boi_1 _22220_ (.A1(_02130_),
    .A2(_02131_),
    .B1_N(_02224_),
    .Y(_02225_));
 sky130_fd_sc_hd__o21a_1 _22221_ (.A1(net5800),
    .A2(net3786),
    .B1(net5780),
    .X(_02226_));
 sky130_fd_sc_hd__a21o_1 _22222_ (.A1(net5800),
    .A2(net3786),
    .B1(_02226_),
    .X(_02227_));
 sky130_fd_sc_hd__or2_2 _22223_ (.A(net5785),
    .B(net5800),
    .X(_02228_));
 sky130_fd_sc_hd__nor2_1 _22224_ (.A(net5762),
    .B(_02228_),
    .Y(_02229_));
 sky130_fd_sc_hd__a211o_1 _22225_ (.A1(net5762),
    .A2(_02227_),
    .B1(_02229_),
    .C1(net3778),
    .X(_02230_));
 sky130_fd_sc_hd__xnor2_1 _22226_ (.A(net2473),
    .B(_02230_),
    .Y(_02231_));
 sky130_fd_sc_hd__xor2_1 _22227_ (.A(net1704),
    .B(net1703),
    .X(_02232_));
 sky130_fd_sc_hd__xnor2_2 _22228_ (.A(_02221_),
    .B(_02232_),
    .Y(_02233_));
 sky130_fd_sc_hd__a21bo_1 _22229_ (.A1(net1389),
    .A2(_02145_),
    .B1_N(_02135_),
    .X(_02234_));
 sky130_fd_sc_hd__o21a_1 _22230_ (.A1(net1389),
    .A2(_02145_),
    .B1(_02234_),
    .X(_02235_));
 sky130_fd_sc_hd__xor2_1 _22231_ (.A(_02233_),
    .B(net1033),
    .X(_02236_));
 sky130_fd_sc_hd__xnor2_2 _22232_ (.A(_02207_),
    .B(_02236_),
    .Y(_02237_));
 sky130_fd_sc_hd__o21a_1 _22233_ (.A1(_02152_),
    .A2(_02155_),
    .B1(net1712),
    .X(_02238_));
 sky130_fd_sc_hd__a21o_1 _22234_ (.A1(_02152_),
    .A2(_02155_),
    .B1(_02238_),
    .X(_02239_));
 sky130_fd_sc_hd__xnor2_2 _22235_ (.A(net2058),
    .B(net943),
    .Y(_02240_));
 sky130_fd_sc_hd__xnor2_1 _22236_ (.A(_02237_),
    .B(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__xnor2_2 _22237_ (.A(net756),
    .B(_02241_),
    .Y(_02242_));
 sky130_fd_sc_hd__o21a_1 _22238_ (.A1(_02160_),
    .A2(_02190_),
    .B1(net2062),
    .X(_02243_));
 sky130_fd_sc_hd__xnor2_1 _22239_ (.A(_02242_),
    .B(_02243_),
    .Y(_02244_));
 sky130_fd_sc_hd__xnor2_1 _22240_ (.A(_02199_),
    .B(_02244_),
    .Y(_02245_));
 sky130_fd_sc_hd__a21o_1 _22241_ (.A1(_02118_),
    .A2(_02166_),
    .B1(_02119_),
    .X(_02246_));
 sky130_fd_sc_hd__o21ai_1 _22242_ (.A1(_02118_),
    .A2(_02166_),
    .B1(_02246_),
    .Y(_02247_));
 sky130_fd_sc_hd__nand2_1 _22243_ (.A(_02245_),
    .B(_02247_),
    .Y(_02248_));
 sky130_fd_sc_hd__nor2_1 _22244_ (.A(_02245_),
    .B(_02247_),
    .Y(_02249_));
 sky130_fd_sc_hd__inv_2 _22245_ (.A(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__nand2_1 _22246_ (.A(_02248_),
    .B(_02250_),
    .Y(_02251_));
 sky130_fd_sc_hd__a21bo_1 _22247_ (.A1(_02115_),
    .A2(_02169_),
    .B1_N(_02170_),
    .X(_02252_));
 sky130_fd_sc_hd__xor2_1 _22248_ (.A(_02251_),
    .B(_02252_),
    .X(_02253_));
 sky130_fd_sc_hd__inv_2 _22249_ (.A(\pid_d.curr_error[10] ),
    .Y(_02254_));
 sky130_fd_sc_hd__o21ba_1 _22250_ (.A1(_02254_),
    .A2(_02176_),
    .B1_N(\pid_d.prev_error[10] ),
    .X(_02255_));
 sky130_fd_sc_hd__a21o_1 _22251_ (.A1(_02254_),
    .A2(_02176_),
    .B1(_02255_),
    .X(_02256_));
 sky130_fd_sc_hd__xnor2_1 _22252_ (.A(\pid_d.prev_error[11] ),
    .B(net5966),
    .Y(_02257_));
 sky130_fd_sc_hd__nand2_1 _22253_ (.A(_02256_),
    .B(_02257_),
    .Y(_02258_));
 sky130_fd_sc_hd__or2_1 _22254_ (.A(_02256_),
    .B(_02257_),
    .X(_02259_));
 sky130_fd_sc_hd__and3_1 _22255_ (.A(net4364),
    .B(_02258_),
    .C(_02259_),
    .X(_02260_));
 sky130_fd_sc_hd__a221o_1 _22256_ (.A1(net4381),
    .A2(_02187_),
    .B1(net299),
    .B2(net4317),
    .C1(net337),
    .X(_02261_));
 sky130_fd_sc_hd__a22o_1 _22257_ (.A1(\pid_d.curr_int[11] ),
    .A2(net3843),
    .B1(net2487),
    .B2(_02261_),
    .X(_00530_));
 sky130_fd_sc_hd__nand2_1 _22258_ (.A(\pid_d.prev_error[12] ),
    .B(\pid_d.curr_error[12] ),
    .Y(_02262_));
 sky130_fd_sc_hd__or2_1 _22259_ (.A(\pid_d.prev_error[12] ),
    .B(\pid_d.curr_error[12] ),
    .X(_02263_));
 sky130_fd_sc_hd__nand2_1 _22260_ (.A(_02262_),
    .B(_02263_),
    .Y(_02264_));
 sky130_fd_sc_hd__nor2_1 _22261_ (.A(\pid_d.prev_error[11] ),
    .B(net5966),
    .Y(_02265_));
 sky130_fd_sc_hd__nand2_1 _22262_ (.A(\pid_d.prev_error[11] ),
    .B(net5966),
    .Y(_02266_));
 sky130_fd_sc_hd__o21ai_1 _22263_ (.A1(_02256_),
    .A2(_02265_),
    .B1(_02266_),
    .Y(_02267_));
 sky130_fd_sc_hd__xnor2_1 _22264_ (.A(_02264_),
    .B(_02267_),
    .Y(_02268_));
 sky130_fd_sc_hd__inv_2 _22265_ (.A(\pid_d.prev_int[11] ),
    .Y(_02269_));
 sky130_fd_sc_hd__inv_2 _22266_ (.A(\pid_d.curr_int[11] ),
    .Y(_02270_));
 sky130_fd_sc_hd__o21a_1 _22267_ (.A1(_02269_),
    .A2(_02185_),
    .B1(_02270_),
    .X(_02271_));
 sky130_fd_sc_hd__a21o_1 _22268_ (.A1(_02269_),
    .A2(_02185_),
    .B1(_02271_),
    .X(_02272_));
 sky130_fd_sc_hd__xor2_1 _22269_ (.A(\pid_d.curr_int[12] ),
    .B(net4391),
    .X(_02273_));
 sky130_fd_sc_hd__xnor2_1 _22270_ (.A(net381),
    .B(_02273_),
    .Y(_02274_));
 sky130_fd_sc_hd__inv_2 _22271_ (.A(_02169_),
    .Y(_02275_));
 sky130_fd_sc_hd__a31o_1 _22272_ (.A1(_02095_),
    .A2(_02114_),
    .A3(_02170_),
    .B1(_02275_),
    .X(_02276_));
 sky130_fd_sc_hd__a21oi_1 _22273_ (.A1(_02248_),
    .A2(_02276_),
    .B1(_02249_),
    .Y(_02277_));
 sky130_fd_sc_hd__o21ba_1 _22274_ (.A1(_02242_),
    .A2(_02243_),
    .B1_N(_02199_),
    .X(_02278_));
 sky130_fd_sc_hd__a21oi_1 _22275_ (.A1(_02242_),
    .A2(_02243_),
    .B1(_02278_),
    .Y(_02279_));
 sky130_fd_sc_hd__a21o_1 _22276_ (.A1(_02233_),
    .A2(net1033),
    .B1(_02207_),
    .X(_02280_));
 sky130_fd_sc_hd__o21ai_2 _22277_ (.A1(_02233_),
    .A2(net1033),
    .B1(_02280_),
    .Y(_02281_));
 sky130_fd_sc_hd__a21bo_1 _22278_ (.A1(net2052),
    .A2(_02219_),
    .B1_N(_02214_),
    .X(_02282_));
 sky130_fd_sc_hd__o21a_1 _22279_ (.A1(net2052),
    .A2(_02219_),
    .B1(_02282_),
    .X(_02283_));
 sky130_fd_sc_hd__nand2_1 _22280_ (.A(net5752),
    .B(net5378),
    .Y(_02284_));
 sky130_fd_sc_hd__nand2_1 _22281_ (.A(net5707),
    .B(net5409),
    .Y(_02285_));
 sky130_fd_sc_hd__nand2_1 _22282_ (.A(net5722),
    .B(net5388),
    .Y(_02286_));
 sky130_fd_sc_hd__xnor2_1 _22283_ (.A(_02285_),
    .B(_02286_),
    .Y(_02287_));
 sky130_fd_sc_hd__xnor2_1 _22284_ (.A(_02284_),
    .B(_02287_),
    .Y(_02288_));
 sky130_fd_sc_hd__o21a_1 _22285_ (.A1(_02210_),
    .A2(_02211_),
    .B1(_02212_),
    .X(_02289_));
 sky130_fd_sc_hd__a21oi_2 _22286_ (.A1(_02210_),
    .A2(_02211_),
    .B1(_02289_),
    .Y(_02290_));
 sky130_fd_sc_hd__nand2_2 _22287_ (.A(_01317_),
    .B(net5646),
    .Y(_02291_));
 sky130_fd_sc_hd__nand2_1 _22288_ (.A(net5465),
    .B(net5670),
    .Y(_02292_));
 sky130_fd_sc_hd__nand2_1 _22289_ (.A(net5691),
    .B(net5435),
    .Y(_02293_));
 sky130_fd_sc_hd__xor2_1 _22290_ (.A(_02292_),
    .B(_02293_),
    .X(_02294_));
 sky130_fd_sc_hd__xnor2_2 _22291_ (.A(_02291_),
    .B(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__xnor2_1 _22292_ (.A(_02290_),
    .B(_02295_),
    .Y(_02296_));
 sky130_fd_sc_hd__xnor2_1 _22293_ (.A(_02288_),
    .B(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__o21a_1 _22294_ (.A1(_02215_),
    .A2(_02216_),
    .B1(_02217_),
    .X(_02298_));
 sky130_fd_sc_hd__a21oi_2 _22295_ (.A1(_02215_),
    .A2(_02216_),
    .B1(_02298_),
    .Y(_02299_));
 sky130_fd_sc_hd__and3_1 _22296_ (.A(net5765),
    .B(net5780),
    .C(net5800),
    .X(_02300_));
 sky130_fd_sc_hd__or3_1 _22297_ (.A(net3778),
    .B(_02229_),
    .C(_02300_),
    .X(_02301_));
 sky130_fd_sc_hd__xnor2_2 _22298_ (.A(_02299_),
    .B(net2471),
    .Y(_02302_));
 sky130_fd_sc_hd__xor2_1 _22299_ (.A(net1702),
    .B(_02302_),
    .X(_02303_));
 sky130_fd_sc_hd__xnor2_2 _22300_ (.A(_02283_),
    .B(_02303_),
    .Y(_02304_));
 sky130_fd_sc_hd__or2_1 _22301_ (.A(net5762),
    .B(_02228_),
    .X(_02305_));
 sky130_fd_sc_hd__nand3_1 _22302_ (.A(net5762),
    .B(net3786),
    .C(_02228_),
    .Y(_02306_));
 sky130_fd_sc_hd__a31o_1 _22303_ (.A1(net2473),
    .A2(_02305_),
    .A3(_02306_),
    .B1(_02300_),
    .X(_02307_));
 sky130_fd_sc_hd__nand2_1 _22304_ (.A(net5380),
    .B(net2051),
    .Y(_02308_));
 sky130_fd_sc_hd__xor2_2 _22305_ (.A(net944),
    .B(_02308_),
    .X(_02309_));
 sky130_fd_sc_hd__a21bo_1 _22306_ (.A1(net1704),
    .A2(net1703),
    .B1_N(_02221_),
    .X(_02310_));
 sky130_fd_sc_hd__o21a_1 _22307_ (.A1(net1704),
    .A2(net1703),
    .B1(_02310_),
    .X(_02311_));
 sky130_fd_sc_hd__xor2_1 _22308_ (.A(_02309_),
    .B(_02311_),
    .X(_02312_));
 sky130_fd_sc_hd__xnor2_2 _22309_ (.A(_02304_),
    .B(_02312_),
    .Y(_02313_));
 sky130_fd_sc_hd__o21a_1 _22310_ (.A1(_02152_),
    .A2(net1706),
    .B1(net1712),
    .X(_02314_));
 sky130_fd_sc_hd__a21o_1 _22311_ (.A1(_02152_),
    .A2(net1706),
    .B1(_02314_),
    .X(_02315_));
 sky130_fd_sc_hd__xnor2_2 _22312_ (.A(net2057),
    .B(_02315_),
    .Y(_02316_));
 sky130_fd_sc_hd__xnor2_1 _22313_ (.A(_02313_),
    .B(_02316_),
    .Y(_02317_));
 sky130_fd_sc_hd__xnor2_2 _22314_ (.A(_02281_),
    .B(_02317_),
    .Y(_02318_));
 sky130_fd_sc_hd__o21ba_1 _22315_ (.A1(_02237_),
    .A2(_02240_),
    .B1_N(net756),
    .X(_02319_));
 sky130_fd_sc_hd__a21o_1 _22316_ (.A1(_02237_),
    .A2(_02240_),
    .B1(_02319_),
    .X(_02320_));
 sky130_fd_sc_hd__nor2_1 _22317_ (.A(net2058),
    .B(net943),
    .Y(_02321_));
 sky130_fd_sc_hd__xor2_1 _22318_ (.A(_02320_),
    .B(_02321_),
    .X(_02322_));
 sky130_fd_sc_hd__xnor2_1 _22319_ (.A(_02318_),
    .B(_02322_),
    .Y(_02323_));
 sky130_fd_sc_hd__or2_1 _22320_ (.A(_02279_),
    .B(net552),
    .X(_02324_));
 sky130_fd_sc_hd__nand2_1 _22321_ (.A(_02279_),
    .B(net552),
    .Y(_02325_));
 sky130_fd_sc_hd__nand2_1 _22322_ (.A(_02324_),
    .B(_02325_),
    .Y(_02326_));
 sky130_fd_sc_hd__xnor2_1 _22323_ (.A(net336),
    .B(_02326_),
    .Y(_02327_));
 sky130_fd_sc_hd__nor2_1 _22324_ (.A(_04887_),
    .B(net297),
    .Y(_02328_));
 sky130_fd_sc_hd__a221o_1 _22325_ (.A1(net4363),
    .A2(_02268_),
    .B1(_02274_),
    .B2(net4380),
    .C1(_02328_),
    .X(_02329_));
 sky130_fd_sc_hd__a22o_1 _22326_ (.A1(\pid_d.curr_int[12] ),
    .A2(net3844),
    .B1(net2489),
    .B2(_02329_),
    .X(_00531_));
 sky130_fd_sc_hd__and2_1 _22327_ (.A(\pid_d.curr_int[13] ),
    .B(\pid_d.prev_int[13] ),
    .X(_02330_));
 sky130_fd_sc_hd__or2_1 _22328_ (.A(\pid_d.curr_int[13] ),
    .B(\pid_d.prev_int[13] ),
    .X(_02331_));
 sky130_fd_sc_hd__or2b_1 _22329_ (.A(_02330_),
    .B_N(_02331_),
    .X(_02332_));
 sky130_fd_sc_hd__o21ba_1 _22330_ (.A1(\pid_d.curr_int[12] ),
    .A2(net4391),
    .B1_N(net381),
    .X(_02333_));
 sky130_fd_sc_hd__and2_1 _22331_ (.A(\pid_d.curr_int[12] ),
    .B(net4391),
    .X(_02334_));
 sky130_fd_sc_hd__or2_1 _22332_ (.A(_02333_),
    .B(_02334_),
    .X(_02335_));
 sky130_fd_sc_hd__xnor2_1 _22333_ (.A(_02332_),
    .B(_02335_),
    .Y(_02336_));
 sky130_fd_sc_hd__a21bo_1 _22334_ (.A1(net336),
    .A2(_02324_),
    .B1_N(_02325_),
    .X(_02337_));
 sky130_fd_sc_hd__o21ba_1 _22335_ (.A1(_02320_),
    .A2(_02318_),
    .B1_N(_02321_),
    .X(_02338_));
 sky130_fd_sc_hd__a21oi_1 _22336_ (.A1(_02320_),
    .A2(_02318_),
    .B1(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hd__a21o_1 _22337_ (.A1(_02304_),
    .A2(_02309_),
    .B1(_02311_),
    .X(_02340_));
 sky130_fd_sc_hd__o21ai_2 _22338_ (.A1(_02304_),
    .A2(_02309_),
    .B1(_02340_),
    .Y(_02341_));
 sky130_fd_sc_hd__o21a_1 _22339_ (.A1(net3829),
    .A2(net2472),
    .B1(net5762),
    .X(_02342_));
 sky130_fd_sc_hd__a21oi_1 _22340_ (.A1(_02228_),
    .A2(net2472),
    .B1(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__nor2_2 _22341_ (.A(net3778),
    .B(_02343_),
    .Y(_02344_));
 sky130_fd_sc_hd__xnor2_2 _22342_ (.A(net944),
    .B(_02344_),
    .Y(_02345_));
 sky130_fd_sc_hd__o21a_1 _22343_ (.A1(_02291_),
    .A2(_02292_),
    .B1(_02293_),
    .X(_02346_));
 sky130_fd_sc_hd__a21oi_2 _22344_ (.A1(_02291_),
    .A2(_02292_),
    .B1(_02346_),
    .Y(_02347_));
 sky130_fd_sc_hd__nand2_1 _22345_ (.A(net5708),
    .B(net5388),
    .Y(_02348_));
 sky130_fd_sc_hd__xor2_1 _22346_ (.A(net5720),
    .B(net5745),
    .X(_02349_));
 sky130_fd_sc_hd__nand2_1 _22347_ (.A(net5378),
    .B(_02349_),
    .Y(_02350_));
 sky130_fd_sc_hd__xor2_2 _22348_ (.A(_02348_),
    .B(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__nand2_2 _22349_ (.A(_01405_),
    .B(net5647),
    .Y(_02352_));
 sky130_fd_sc_hd__nand2_1 _22350_ (.A(net5438),
    .B(net5670),
    .Y(_02353_));
 sky130_fd_sc_hd__nand2_1 _22351_ (.A(net5694),
    .B(net5411),
    .Y(_02354_));
 sky130_fd_sc_hd__xor2_1 _22352_ (.A(_02353_),
    .B(_02354_),
    .X(_02355_));
 sky130_fd_sc_hd__xnor2_2 _22353_ (.A(_02352_),
    .B(_02355_),
    .Y(_02356_));
 sky130_fd_sc_hd__xor2_1 _22354_ (.A(_02351_),
    .B(_02356_),
    .X(_02357_));
 sky130_fd_sc_hd__xnor2_2 _22355_ (.A(_02347_),
    .B(_02357_),
    .Y(_02358_));
 sky130_fd_sc_hd__a21bo_1 _22356_ (.A1(_02290_),
    .A2(_02295_),
    .B1_N(_02288_),
    .X(_02359_));
 sky130_fd_sc_hd__o21a_1 _22357_ (.A1(_02290_),
    .A2(_02295_),
    .B1(_02359_),
    .X(_02360_));
 sky130_fd_sc_hd__o21a_1 _22358_ (.A1(_02284_),
    .A2(_02286_),
    .B1(_02285_),
    .X(_02361_));
 sky130_fd_sc_hd__a21oi_1 _22359_ (.A1(_02284_),
    .A2(_02286_),
    .B1(_02361_),
    .Y(_02362_));
 sky130_fd_sc_hd__xnor2_1 _22360_ (.A(net2471),
    .B(_02362_),
    .Y(_02363_));
 sky130_fd_sc_hd__nor2_1 _22361_ (.A(_02360_),
    .B(_02363_),
    .Y(_02364_));
 sky130_fd_sc_hd__nand2_1 _22362_ (.A(_02360_),
    .B(_02363_),
    .Y(_02365_));
 sky130_fd_sc_hd__and2b_1 _22363_ (.A_N(_02364_),
    .B(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__xnor2_2 _22364_ (.A(_02358_),
    .B(_02366_),
    .Y(_02367_));
 sky130_fd_sc_hd__a21bo_1 _22365_ (.A1(_02283_),
    .A2(_02302_),
    .B1_N(net1702),
    .X(_02368_));
 sky130_fd_sc_hd__o21a_1 _22366_ (.A1(_02283_),
    .A2(_02302_),
    .B1(_02368_),
    .X(_02369_));
 sky130_fd_sc_hd__xor2_1 _22367_ (.A(_02367_),
    .B(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__xnor2_1 _22368_ (.A(_02345_),
    .B(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__a31o_1 _22369_ (.A1(net5841),
    .A2(net5862),
    .A3(net2067),
    .B1(net2051),
    .X(_02372_));
 sky130_fd_sc_hd__nand2_1 _22370_ (.A(net1715),
    .B(_01964_),
    .Y(_02373_));
 sky130_fd_sc_hd__a22o_1 _22371_ (.A1(net5817),
    .A2(_02372_),
    .B1(_02373_),
    .B2(net2051),
    .X(_02374_));
 sky130_fd_sc_hd__nand2_1 _22372_ (.A(net5380),
    .B(_02374_),
    .Y(_02375_));
 sky130_fd_sc_hd__xnor2_1 _22373_ (.A(net2476),
    .B(_02375_),
    .Y(_02376_));
 sky130_fd_sc_hd__and2_1 _22374_ (.A(_02371_),
    .B(_02376_),
    .X(_02377_));
 sky130_fd_sc_hd__or2_1 _22375_ (.A(_02371_),
    .B(_02376_),
    .X(_02378_));
 sky130_fd_sc_hd__and2b_1 _22376_ (.A_N(_02377_),
    .B(_02378_),
    .X(_02379_));
 sky130_fd_sc_hd__xnor2_2 _22377_ (.A(_02341_),
    .B(_02379_),
    .Y(_02380_));
 sky130_fd_sc_hd__o21a_1 _22378_ (.A1(_02313_),
    .A2(_02316_),
    .B1(_02281_),
    .X(_02381_));
 sky130_fd_sc_hd__a21o_1 _22379_ (.A1(_02313_),
    .A2(_02316_),
    .B1(_02381_),
    .X(_02382_));
 sky130_fd_sc_hd__nor2_1 _22380_ (.A(net2057),
    .B(_02315_),
    .Y(_02383_));
 sky130_fd_sc_hd__xor2_1 _22381_ (.A(_02382_),
    .B(_02383_),
    .X(_02384_));
 sky130_fd_sc_hd__xnor2_1 _22382_ (.A(_02380_),
    .B(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__or2_1 _22383_ (.A(net551),
    .B(net549),
    .X(_02386_));
 sky130_fd_sc_hd__inv_2 _22384_ (.A(_02386_),
    .Y(_02387_));
 sky130_fd_sc_hd__and2_1 _22385_ (.A(net551),
    .B(net549),
    .X(_02388_));
 sky130_fd_sc_hd__nor2_1 _22386_ (.A(_02387_),
    .B(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__xnor2_1 _22387_ (.A(_02337_),
    .B(_02389_),
    .Y(_02390_));
 sky130_fd_sc_hd__nand2_1 _22388_ (.A(_02263_),
    .B(_02267_),
    .Y(_02391_));
 sky130_fd_sc_hd__xor2_1 _22389_ (.A(\pid_d.prev_error[13] ),
    .B(net5965),
    .X(_02392_));
 sky130_fd_sc_hd__and3_1 _22390_ (.A(_02262_),
    .B(_02391_),
    .C(_02392_),
    .X(_02393_));
 sky130_fd_sc_hd__a21oi_1 _22391_ (.A1(_02262_),
    .A2(_02391_),
    .B1(_02392_),
    .Y(_02394_));
 sky130_fd_sc_hd__o21a_1 _22392_ (.A1(_02393_),
    .A2(_02394_),
    .B1(net4364),
    .X(_02395_));
 sky130_fd_sc_hd__a221o_1 _22393_ (.A1(net4382),
    .A2(_02336_),
    .B1(net272),
    .B2(net4316),
    .C1(_02395_),
    .X(_02396_));
 sky130_fd_sc_hd__a22o_1 _22394_ (.A1(\pid_d.curr_int[13] ),
    .A2(net3844),
    .B1(net2488),
    .B2(_02396_),
    .X(_00532_));
 sky130_fd_sc_hd__o31a_1 _22395_ (.A1(_02330_),
    .A2(_02333_),
    .A3(_02334_),
    .B1(_02331_),
    .X(_02397_));
 sky130_fd_sc_hd__xor2_1 _22396_ (.A(\pid_d.curr_int[14] ),
    .B(\pid_d.prev_int[14] ),
    .X(_02398_));
 sky130_fd_sc_hd__or2_1 _22397_ (.A(_02397_),
    .B(_02398_),
    .X(_02399_));
 sky130_fd_sc_hd__nand2_1 _22398_ (.A(_02397_),
    .B(_02398_),
    .Y(_02400_));
 sky130_fd_sc_hd__a2bb2o_1 _22399_ (.A1_N(\pid_d.prev_error[13] ),
    .A2_N(net5965),
    .B1(_02262_),
    .B2(_02391_),
    .X(_02401_));
 sky130_fd_sc_hd__a21bo_1 _22400_ (.A1(\pid_d.prev_error[13] ),
    .A2(net5965),
    .B1_N(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__and2_1 _22401_ (.A(\pid_d.prev_error[14] ),
    .B(\pid_d.curr_error[14] ),
    .X(_02403_));
 sky130_fd_sc_hd__or2_1 _22402_ (.A(\pid_d.prev_error[14] ),
    .B(\pid_d.curr_error[14] ),
    .X(_02404_));
 sky130_fd_sc_hd__or2b_1 _22403_ (.A(_02403_),
    .B_N(_02404_),
    .X(_02405_));
 sky130_fd_sc_hd__xor2_1 _22404_ (.A(_02402_),
    .B(_02405_),
    .X(_02406_));
 sky130_fd_sc_hd__nor2_1 _22405_ (.A(_04872_),
    .B(_02406_),
    .Y(_02407_));
 sky130_fd_sc_hd__a31o_1 _22406_ (.A1(net4382),
    .A2(_02399_),
    .A3(_02400_),
    .B1(net206),
    .X(_02408_));
 sky130_fd_sc_hd__inv_2 _22407_ (.A(net549),
    .Y(_02409_));
 sky130_fd_sc_hd__o21ba_1 _22408_ (.A1(_02337_),
    .A2(_02409_),
    .B1_N(net551),
    .X(_02410_));
 sky130_fd_sc_hd__a21o_1 _22409_ (.A1(_02337_),
    .A2(_02409_),
    .B1(_02410_),
    .X(_02411_));
 sky130_fd_sc_hd__inv_2 _22410_ (.A(_02380_),
    .Y(_02412_));
 sky130_fd_sc_hd__nand2_1 _22411_ (.A(_02382_),
    .B(_02412_),
    .Y(_02413_));
 sky130_fd_sc_hd__nor2_1 _22412_ (.A(_02382_),
    .B(_02412_),
    .Y(_02414_));
 sky130_fd_sc_hd__a21o_1 _22413_ (.A1(_02383_),
    .A2(_02413_),
    .B1(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__a21o_1 _22414_ (.A1(_02367_),
    .A2(_02345_),
    .B1(_02369_),
    .X(_02416_));
 sky130_fd_sc_hd__o21ai_2 _22415_ (.A1(_02367_),
    .A2(_02345_),
    .B1(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__a21o_1 _22416_ (.A1(_02352_),
    .A2(_02353_),
    .B1(_02354_),
    .X(_02418_));
 sky130_fd_sc_hd__o21ai_2 _22417_ (.A1(_02352_),
    .A2(_02353_),
    .B1(_02418_),
    .Y(_02419_));
 sky130_fd_sc_hd__and2b_1 _22418_ (.A_N(net5434),
    .B(net5646),
    .X(_02420_));
 sky130_fd_sc_hd__nand2_1 _22419_ (.A(net5691),
    .B(net5390),
    .Y(_02421_));
 sky130_fd_sc_hd__nand2_1 _22420_ (.A(net5412),
    .B(net5676),
    .Y(_02422_));
 sky130_fd_sc_hd__xnor2_1 _22421_ (.A(_02421_),
    .B(_02422_),
    .Y(_02423_));
 sky130_fd_sc_hd__xnor2_2 _22422_ (.A(_02420_),
    .B(_02423_),
    .Y(_02424_));
 sky130_fd_sc_hd__nor2_1 _22423_ (.A(net5708),
    .B(_02349_),
    .Y(_02425_));
 sky130_fd_sc_hd__and2_1 _22424_ (.A(net5708),
    .B(_02349_),
    .X(_02426_));
 sky130_fd_sc_hd__or3_1 _22425_ (.A(net3777),
    .B(_02425_),
    .C(_02426_),
    .X(_02427_));
 sky130_fd_sc_hd__xor2_1 _22426_ (.A(_02424_),
    .B(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__xnor2_2 _22427_ (.A(_02419_),
    .B(_02428_),
    .Y(_02429_));
 sky130_fd_sc_hd__a21o_1 _22428_ (.A1(_02351_),
    .A2(_02356_),
    .B1(_02347_),
    .X(_02430_));
 sky130_fd_sc_hd__o21a_1 _22429_ (.A1(_02351_),
    .A2(_02356_),
    .B1(_02430_),
    .X(_02431_));
 sky130_fd_sc_hd__a22o_1 _22430_ (.A1(net5723),
    .A2(net5749),
    .B1(net5389),
    .B2(net5711),
    .X(_02432_));
 sky130_fd_sc_hd__o21ai_2 _22431_ (.A1(net5723),
    .A2(net5749),
    .B1(_02432_),
    .Y(_02433_));
 sky130_fd_sc_hd__or3_1 _22432_ (.A(_02229_),
    .B(_02300_),
    .C(_02433_),
    .X(_02434_));
 sky130_fd_sc_hd__o21ai_1 _22433_ (.A1(_02229_),
    .A2(_02300_),
    .B1(_02433_),
    .Y(_02435_));
 sky130_fd_sc_hd__and3_1 _22434_ (.A(net5377),
    .B(_02434_),
    .C(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__xnor2_1 _22435_ (.A(_02431_),
    .B(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__xnor2_2 _22436_ (.A(_02429_),
    .B(_02437_),
    .Y(_02438_));
 sky130_fd_sc_hd__a21o_1 _22437_ (.A1(_02358_),
    .A2(_02365_),
    .B1(_02364_),
    .X(_02439_));
 sky130_fd_sc_hd__xor2_1 _22438_ (.A(_02438_),
    .B(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__nand2_1 _22439_ (.A(net1712),
    .B(_02152_),
    .Y(_02441_));
 sky130_fd_sc_hd__o21a_1 _22440_ (.A1(net1169),
    .A2(_02344_),
    .B1(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__xnor2_2 _22441_ (.A(net2060),
    .B(_02442_),
    .Y(_02443_));
 sky130_fd_sc_hd__or2_1 _22442_ (.A(net3829),
    .B(net2470),
    .X(_02444_));
 sky130_fd_sc_hd__a22o_1 _22443_ (.A1(_02228_),
    .A2(net2470),
    .B1(_02444_),
    .B2(net5765),
    .X(_02445_));
 sky130_fd_sc_hd__nand2_1 _22444_ (.A(net5377),
    .B(_02445_),
    .Y(_02446_));
 sky130_fd_sc_hd__xnor2_2 _22445_ (.A(net944),
    .B(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__xor2_1 _22446_ (.A(_02443_),
    .B(_02447_),
    .X(_02448_));
 sky130_fd_sc_hd__xnor2_1 _22447_ (.A(_02440_),
    .B(_02448_),
    .Y(_02449_));
 sky130_fd_sc_hd__xnor2_2 _22448_ (.A(_02417_),
    .B(_02449_),
    .Y(_02450_));
 sky130_fd_sc_hd__o21ai_2 _22449_ (.A1(_02341_),
    .A2(_02377_),
    .B1(_02378_),
    .Y(_02451_));
 sky130_fd_sc_hd__nor2_1 _22450_ (.A(net2057),
    .B(_02375_),
    .Y(_02452_));
 sky130_fd_sc_hd__xnor2_1 _22451_ (.A(_02451_),
    .B(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__xnor2_1 _22452_ (.A(_02450_),
    .B(_02453_),
    .Y(_02454_));
 sky130_fd_sc_hd__or2_1 _22453_ (.A(net520),
    .B(net597),
    .X(_02455_));
 sky130_fd_sc_hd__inv_2 _22454_ (.A(_02455_),
    .Y(_02456_));
 sky130_fd_sc_hd__and2_1 _22455_ (.A(net520),
    .B(net597),
    .X(_02457_));
 sky130_fd_sc_hd__nor2_1 _22456_ (.A(_02456_),
    .B(_02457_),
    .Y(_02458_));
 sky130_fd_sc_hd__xnor2_1 _22457_ (.A(_02411_),
    .B(_02458_),
    .Y(_02459_));
 sky130_fd_sc_hd__and3_1 _22458_ (.A(net4316),
    .B(net2488),
    .C(net205),
    .X(_02460_));
 sky130_fd_sc_hd__a221o_1 _22459_ (.A1(\pid_d.curr_int[14] ),
    .A2(_12499_),
    .B1(net2488),
    .B2(_02408_),
    .C1(_02460_),
    .X(_00533_));
 sky130_fd_sc_hd__o21ai_1 _22460_ (.A1(_02402_),
    .A2(_02403_),
    .B1(_02404_),
    .Y(_02461_));
 sky130_fd_sc_hd__xnor2_1 _22461_ (.A(\pid_d.prev_error[15] ),
    .B(net5964),
    .Y(_02462_));
 sky130_fd_sc_hd__xnor2_1 _22462_ (.A(_02461_),
    .B(_02462_),
    .Y(_02463_));
 sky130_fd_sc_hd__xnor2_1 _22463_ (.A(\pid_d.curr_int[15] ),
    .B(\pid_d.prev_int[15] ),
    .Y(_02464_));
 sky130_fd_sc_hd__a21o_1 _22464_ (.A1(\pid_d.prev_int[14] ),
    .A2(_02397_),
    .B1(\pid_d.curr_int[14] ),
    .X(_02465_));
 sky130_fd_sc_hd__o21a_1 _22465_ (.A1(\pid_d.prev_int[14] ),
    .A2(_02397_),
    .B1(_02465_),
    .X(_02466_));
 sky130_fd_sc_hd__xnor2_1 _22466_ (.A(_02464_),
    .B(_02466_),
    .Y(_02467_));
 sky130_fd_sc_hd__a2bb2o_1 _22467_ (.A1_N(net4297),
    .A2_N(_02463_),
    .B1(_02467_),
    .B2(net4379),
    .X(_02468_));
 sky130_fd_sc_hd__a21oi_1 _22468_ (.A1(_02344_),
    .A2(_02446_),
    .B1(net1169),
    .Y(_02469_));
 sky130_fd_sc_hd__mux2_1 _22469_ (.A0(net1169),
    .A1(_02344_),
    .S(net2060),
    .X(_02470_));
 sky130_fd_sc_hd__o221a_1 _22470_ (.A1(net2056),
    .A2(_02469_),
    .B1(_02470_),
    .B2(_02446_),
    .C1(_02441_),
    .X(_02471_));
 sky130_fd_sc_hd__nand3_1 _22471_ (.A(net5713),
    .B(net5721),
    .C(net5746),
    .Y(_02472_));
 sky130_fd_sc_hd__or3_1 _22472_ (.A(net5713),
    .B(net5732),
    .C(net5753),
    .X(_02473_));
 sky130_fd_sc_hd__and3_1 _22473_ (.A(net5689),
    .B(_02472_),
    .C(_02473_),
    .X(_02474_));
 sky130_fd_sc_hd__a21oi_1 _22474_ (.A1(_02472_),
    .A2(_02473_),
    .B1(net5689),
    .Y(_02475_));
 sky130_fd_sc_hd__or3_1 _22475_ (.A(net3778),
    .B(_02474_),
    .C(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__xnor2_1 _22476_ (.A(net2055),
    .B(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__or2_1 _22477_ (.A(net3829),
    .B(_02433_),
    .X(_02478_));
 sky130_fd_sc_hd__a22o_1 _22478_ (.A1(_02228_),
    .A2(_02433_),
    .B1(_02478_),
    .B2(net5765),
    .X(_02479_));
 sky130_fd_sc_hd__nand2_1 _22479_ (.A(net5377),
    .B(_02479_),
    .Y(_02480_));
 sky130_fd_sc_hd__xnor2_1 _22480_ (.A(_02477_),
    .B(_02480_),
    .Y(_02481_));
 sky130_fd_sc_hd__a21bo_1 _22481_ (.A1(net5407),
    .A2(net5434),
    .B1_N(net5647),
    .X(_02482_));
 sky130_fd_sc_hd__and2b_1 _22482_ (.A_N(net5433),
    .B(net5692),
    .X(_02483_));
 sky130_fd_sc_hd__and2b_1 _22483_ (.A_N(net5671),
    .B(net5647),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _22484_ (.A0(net5671),
    .A1(_02484_),
    .S(net5407),
    .X(_02485_));
 sky130_fd_sc_hd__a32o_1 _22485_ (.A1(net5671),
    .A2(_02354_),
    .A3(_02482_),
    .B1(_02483_),
    .B2(_02485_),
    .X(_02486_));
 sky130_fd_sc_hd__o21a_1 _22486_ (.A1(net5671),
    .A2(_02483_),
    .B1(net5390),
    .X(_02487_));
 sky130_fd_sc_hd__or3b_1 _22487_ (.A(net5434),
    .B(net5390),
    .C_N(net5671),
    .X(_02488_));
 sky130_fd_sc_hd__o21ai_1 _22488_ (.A1(net5407),
    .A2(_02487_),
    .B1(_02488_),
    .Y(_02489_));
 sky130_fd_sc_hd__a22o_1 _22489_ (.A1(net5390),
    .A2(_02486_),
    .B1(_02489_),
    .B2(net5647),
    .X(_02490_));
 sky130_fd_sc_hd__a21bo_1 _22490_ (.A1(_02419_),
    .A2(_02424_),
    .B1_N(_02427_),
    .X(_02491_));
 sky130_fd_sc_hd__o21ai_1 _22491_ (.A1(_02419_),
    .A2(_02424_),
    .B1(_02491_),
    .Y(_02492_));
 sky130_fd_sc_hd__xnor2_1 _22492_ (.A(_02490_),
    .B(_02492_),
    .Y(_02493_));
 sky130_fd_sc_hd__xnor2_1 _22493_ (.A(_02481_),
    .B(_02493_),
    .Y(_02494_));
 sky130_fd_sc_hd__a21o_1 _22494_ (.A1(_02429_),
    .A2(_02436_),
    .B1(_02431_),
    .X(_02495_));
 sky130_fd_sc_hd__o21a_1 _22495_ (.A1(_02429_),
    .A2(_02436_),
    .B1(_02495_),
    .X(_02496_));
 sky130_fd_sc_hd__xnor2_1 _22496_ (.A(_02494_),
    .B(_02496_),
    .Y(_02497_));
 sky130_fd_sc_hd__xnor2_1 _22497_ (.A(_02471_),
    .B(_02497_),
    .Y(_02498_));
 sky130_fd_sc_hd__nand2_1 _22498_ (.A(_02443_),
    .B(_02439_),
    .Y(_02499_));
 sky130_fd_sc_hd__nor2_1 _22499_ (.A(_02438_),
    .B(_02499_),
    .Y(_02500_));
 sky130_fd_sc_hd__nor2_1 _22500_ (.A(_02443_),
    .B(_02439_),
    .Y(_02501_));
 sky130_fd_sc_hd__nand2_1 _22501_ (.A(_02438_),
    .B(_02501_),
    .Y(_02502_));
 sky130_fd_sc_hd__nor2_1 _22502_ (.A(_02447_),
    .B(_02502_),
    .Y(_02503_));
 sky130_fd_sc_hd__o21ai_1 _22503_ (.A1(_02438_),
    .A2(_02501_),
    .B1(_02499_),
    .Y(_02504_));
 sky130_fd_sc_hd__o21ai_1 _22504_ (.A1(_02447_),
    .A2(_02504_),
    .B1(_02502_),
    .Y(_02505_));
 sky130_fd_sc_hd__a21o_1 _22505_ (.A1(_02447_),
    .A2(_02504_),
    .B1(_02500_),
    .X(_02506_));
 sky130_fd_sc_hd__mux2_1 _22506_ (.A0(_02505_),
    .A1(_02506_),
    .S(_02417_),
    .X(_02507_));
 sky130_fd_sc_hd__a211o_1 _22507_ (.A1(_02447_),
    .A2(_02500_),
    .B1(_02503_),
    .C1(_02507_),
    .X(_02508_));
 sky130_fd_sc_hd__xnor2_1 _22508_ (.A(_02498_),
    .B(_02508_),
    .Y(_02509_));
 sky130_fd_sc_hd__a21o_1 _22509_ (.A1(_02451_),
    .A2(_02450_),
    .B1(_02452_),
    .X(_02510_));
 sky130_fd_sc_hd__o21a_1 _22510_ (.A1(_02451_),
    .A2(_02450_),
    .B1(_02510_),
    .X(_02511_));
 sky130_fd_sc_hd__xnor2_1 _22511_ (.A(_02509_),
    .B(_02511_),
    .Y(_02512_));
 sky130_fd_sc_hd__mux2_1 _22512_ (.A0(_02456_),
    .A1(_02457_),
    .S(net517),
    .X(_02513_));
 sky130_fd_sc_hd__and2_1 _22513_ (.A(_02455_),
    .B(net517),
    .X(_02514_));
 sky130_fd_sc_hd__nor2_1 _22514_ (.A(_02457_),
    .B(net517),
    .Y(_02515_));
 sky130_fd_sc_hd__mux2_1 _22515_ (.A0(_02514_),
    .A1(_02515_),
    .S(_02411_),
    .X(_02516_));
 sky130_fd_sc_hd__o211a_1 _22516_ (.A1(net380),
    .A2(net204),
    .B1(net4315),
    .C1(net2489),
    .X(_02517_));
 sky130_fd_sc_hd__a221o_1 _22517_ (.A1(net9195),
    .A2(_12499_),
    .B1(net2489),
    .B2(_02468_),
    .C1(_02517_),
    .X(_00534_));
 sky130_fd_sc_hd__or4_1 _22518_ (.A(net4390),
    .B(net4380),
    .C(net4316),
    .D(net4346),
    .X(_02518_));
 sky130_fd_sc_hd__clkbuf_1 _22519_ (.A(_02518_),
    .X(_02519_));
 sky130_fd_sc_hd__buf_1 _22520_ (.A(net3105),
    .X(_02520_));
 sky130_fd_sc_hd__o21a_1 _22521_ (.A1(net4325),
    .A2(net2462),
    .B1(net8887),
    .X(_02521_));
 sky130_fd_sc_hd__clkbuf_1 _22522_ (.A(net2050),
    .X(_02522_));
 sky130_fd_sc_hd__o21ai_1 _22523_ (.A1(net4325),
    .A2(net3101),
    .B1(net8887),
    .Y(_02523_));
 sky130_fd_sc_hd__clkbuf_1 _22524_ (.A(_02523_),
    .X(_02524_));
 sky130_fd_sc_hd__and3_1 _22525_ (.A(net5973),
    .B(net2379),
    .C(net2046),
    .X(_02525_));
 sky130_fd_sc_hd__a21o_1 _22526_ (.A1(\pid_d.prev_error[0] ),
    .A2(net1699),
    .B1(_02525_),
    .X(_00535_));
 sky130_fd_sc_hd__and3_1 _22527_ (.A(net5972),
    .B(net2379),
    .C(net2046),
    .X(_02526_));
 sky130_fd_sc_hd__a21o_1 _22528_ (.A1(net9182),
    .A2(net1699),
    .B1(_02526_),
    .X(_00536_));
 sky130_fd_sc_hd__and3_1 _22529_ (.A(net5971),
    .B(net2379),
    .C(net2046),
    .X(_02527_));
 sky130_fd_sc_hd__a21o_1 _22530_ (.A1(net9135),
    .A2(net1699),
    .B1(_02527_),
    .X(_00537_));
 sky130_fd_sc_hd__and3_1 _22531_ (.A(net5970),
    .B(net2380),
    .C(net2046),
    .X(_02528_));
 sky130_fd_sc_hd__a21o_1 _22532_ (.A1(net9106),
    .A2(net1699),
    .B1(_02528_),
    .X(_00538_));
 sky130_fd_sc_hd__and3_1 _22533_ (.A(\pid_d.curr_error[4] ),
    .B(net2380),
    .C(net2047),
    .X(_02529_));
 sky130_fd_sc_hd__a21o_1 _22534_ (.A1(net9138),
    .A2(net1700),
    .B1(_02529_),
    .X(_00539_));
 sky130_fd_sc_hd__and3_1 _22535_ (.A(net5969),
    .B(net2379),
    .C(net2047),
    .X(_02530_));
 sky130_fd_sc_hd__a21o_1 _22536_ (.A1(net9124),
    .A2(net1700),
    .B1(_02530_),
    .X(_00540_));
 sky130_fd_sc_hd__and3_1 _22537_ (.A(net5968),
    .B(net2381),
    .C(net2047),
    .X(_02531_));
 sky130_fd_sc_hd__a21o_1 _22538_ (.A1(net9117),
    .A2(net1700),
    .B1(_02531_),
    .X(_00541_));
 sky130_fd_sc_hd__and3_1 _22539_ (.A(\pid_d.curr_error[7] ),
    .B(net2381),
    .C(net2048),
    .X(_02532_));
 sky130_fd_sc_hd__a21o_1 _22540_ (.A1(net9114),
    .A2(net1701),
    .B1(_02532_),
    .X(_00542_));
 sky130_fd_sc_hd__and3_1 _22541_ (.A(\pid_d.curr_error[8] ),
    .B(net2381),
    .C(net2048),
    .X(_02533_));
 sky130_fd_sc_hd__a21o_1 _22542_ (.A1(net9119),
    .A2(net1701),
    .B1(_02533_),
    .X(_00543_));
 sky130_fd_sc_hd__and3_1 _22543_ (.A(net5967),
    .B(net3016),
    .C(net2048),
    .X(_02534_));
 sky130_fd_sc_hd__a21o_1 _22544_ (.A1(net9105),
    .A2(net1701),
    .B1(_02534_),
    .X(_00544_));
 sky130_fd_sc_hd__and3_1 _22545_ (.A(\pid_d.curr_error[10] ),
    .B(net3016),
    .C(net2461),
    .X(_02535_));
 sky130_fd_sc_hd__a21o_1 _22546_ (.A1(net9121),
    .A2(net2050),
    .B1(_02535_),
    .X(_00545_));
 sky130_fd_sc_hd__and3_1 _22547_ (.A(net5966),
    .B(net3017),
    .C(net2461),
    .X(_02536_));
 sky130_fd_sc_hd__a21o_1 _22548_ (.A1(net9181),
    .A2(_02521_),
    .B1(_02536_),
    .X(_00546_));
 sky130_fd_sc_hd__and3_1 _22549_ (.A(\pid_d.curr_error[12] ),
    .B(net3017),
    .C(net2460),
    .X(_02537_));
 sky130_fd_sc_hd__a21o_1 _22550_ (.A1(net9012),
    .A2(net2049),
    .B1(_02537_),
    .X(_00547_));
 sky130_fd_sc_hd__and3_1 _22551_ (.A(net5965),
    .B(net3018),
    .C(net2460),
    .X(_02538_));
 sky130_fd_sc_hd__a21o_1 _22552_ (.A1(net9159),
    .A2(net2049),
    .B1(_02538_),
    .X(_00548_));
 sky130_fd_sc_hd__and3_1 _22553_ (.A(\pid_d.curr_error[14] ),
    .B(net3018),
    .C(net2460),
    .X(_02539_));
 sky130_fd_sc_hd__a21o_1 _22554_ (.A1(net8988),
    .A2(net2049),
    .B1(_02539_),
    .X(_00549_));
 sky130_fd_sc_hd__and3_1 _22555_ (.A(net5964),
    .B(net3017),
    .C(net2461),
    .X(_02540_));
 sky130_fd_sc_hd__a21o_1 _22556_ (.A1(net9083),
    .A2(_02521_),
    .B1(_02540_),
    .X(_00550_));
 sky130_fd_sc_hd__nor4_1 _22557_ (.A(net4390),
    .B(net4380),
    .C(net4315),
    .D(net4327),
    .Y(_02541_));
 sky130_fd_sc_hd__nor2_1 _22558_ (.A(_04865_),
    .B(net3775),
    .Y(_02542_));
 sky130_fd_sc_hd__or2_1 _22559_ (.A(_04873_),
    .B(_02542_),
    .X(_02543_));
 sky130_fd_sc_hd__buf_1 _22560_ (.A(net2459),
    .X(_02544_));
 sky130_fd_sc_hd__and3_1 _22561_ (.A(net6754),
    .B(net6603),
    .C(net4347),
    .X(_02545_));
 sky130_fd_sc_hd__and3_1 _22562_ (.A(net8887),
    .B(net4301),
    .C(net3774),
    .X(_02546_));
 sky130_fd_sc_hd__and2_1 _22563_ (.A(net3768),
    .B(net3093),
    .X(_02547_));
 sky130_fd_sc_hd__clkbuf_2 _22564_ (.A(_02547_),
    .X(_02548_));
 sky130_fd_sc_hd__a22o_1 _22565_ (.A1(net8987),
    .A2(net2043),
    .B1(_02548_),
    .B2(net7368),
    .X(_00551_));
 sky130_fd_sc_hd__xor2_1 _22566_ (.A(net7368),
    .B(net7353),
    .X(_02549_));
 sky130_fd_sc_hd__a22o_1 _22567_ (.A1(net9037),
    .A2(net2043),
    .B1(_02548_),
    .B2(_02549_),
    .X(_00552_));
 sky130_fd_sc_hd__o21ai_1 _22568_ (.A1(net7369),
    .A2(net7352),
    .B1(net7343),
    .Y(_02550_));
 sky130_fd_sc_hd__or3_1 _22569_ (.A(net7369),
    .B(net7352),
    .C(net7343),
    .X(_02551_));
 sky130_fd_sc_hd__and3_1 _22570_ (.A(net3769),
    .B(_02550_),
    .C(_02551_),
    .X(_02552_));
 sky130_fd_sc_hd__a22o_1 _22571_ (.A1(net9050),
    .A2(net2043),
    .B1(net3093),
    .B2(net3092),
    .X(_00553_));
 sky130_fd_sc_hd__buf_1 _22572_ (.A(net3768),
    .X(_02553_));
 sky130_fd_sc_hd__or2_1 _22573_ (.A(net7329),
    .B(_02551_),
    .X(_02554_));
 sky130_fd_sc_hd__nand2_1 _22574_ (.A(net7329),
    .B(_02551_),
    .Y(_02555_));
 sky130_fd_sc_hd__and3_1 _22575_ (.A(net3091),
    .B(_02554_),
    .C(_02555_),
    .X(_02556_));
 sky130_fd_sc_hd__a22o_1 _22576_ (.A1(net9028),
    .A2(net2043),
    .B1(net3093),
    .B2(net2458),
    .X(_00554_));
 sky130_fd_sc_hd__or2_1 _22577_ (.A(net7317),
    .B(_02554_),
    .X(_02557_));
 sky130_fd_sc_hd__nand2_1 _22578_ (.A(net7317),
    .B(_02554_),
    .Y(_02558_));
 sky130_fd_sc_hd__and3_1 _22579_ (.A(net3769),
    .B(_02557_),
    .C(_02558_),
    .X(_02559_));
 sky130_fd_sc_hd__or4_1 _22580_ (.A(net4390),
    .B(\pid_d.state[1] ),
    .C(net4315),
    .D(net4326),
    .X(_02560_));
 sky130_fd_sc_hd__nor2_1 _22581_ (.A(net4367),
    .B(net3767),
    .Y(_02561_));
 sky130_fd_sc_hd__mux2_1 _22582_ (.A0(\pid_d.curr_error[4] ),
    .A1(net2040),
    .S(net3087),
    .X(_02562_));
 sky130_fd_sc_hd__and2_1 _22583_ (.A(net8891),
    .B(_02562_),
    .X(_02563_));
 sky130_fd_sc_hd__clkbuf_1 _22584_ (.A(_02563_),
    .X(_00555_));
 sky130_fd_sc_hd__or3_1 _22585_ (.A(net7317),
    .B(net7306),
    .C(_02554_),
    .X(_02564_));
 sky130_fd_sc_hd__o21ai_1 _22586_ (.A1(net7317),
    .A2(_02554_),
    .B1(net7306),
    .Y(_02565_));
 sky130_fd_sc_hd__a32o_1 _22587_ (.A1(_02548_),
    .A2(_02564_),
    .A3(_02565_),
    .B1(net2044),
    .B2(net8957),
    .X(_00556_));
 sky130_fd_sc_hd__or2_1 _22588_ (.A(net7294),
    .B(_02564_),
    .X(_02566_));
 sky130_fd_sc_hd__nand2_1 _22589_ (.A(net7294),
    .B(_02564_),
    .Y(_02567_));
 sky130_fd_sc_hd__and3_1 _22590_ (.A(net3091),
    .B(_02566_),
    .C(_02567_),
    .X(_02568_));
 sky130_fd_sc_hd__a22o_1 _22591_ (.A1(net5968),
    .A2(net2044),
    .B1(net3093),
    .B2(net1698),
    .X(_00557_));
 sky130_fd_sc_hd__nor2_1 _22592_ (.A(net7287),
    .B(_02566_),
    .Y(_02569_));
 sky130_fd_sc_hd__nand2_1 _22593_ (.A(net7287),
    .B(_02566_),
    .Y(_02570_));
 sky130_fd_sc_hd__and3b_1 _22594_ (.A_N(_02569_),
    .B(_02570_),
    .C(net3768),
    .X(_02571_));
 sky130_fd_sc_hd__mux2_1 _22595_ (.A0(\pid_d.curr_error[7] ),
    .A1(net1388),
    .S(net3087),
    .X(_02572_));
 sky130_fd_sc_hd__and2_1 _22596_ (.A(net8889),
    .B(_02572_),
    .X(_02573_));
 sky130_fd_sc_hd__clkbuf_1 _22597_ (.A(_02573_),
    .X(_00558_));
 sky130_fd_sc_hd__nand2_1 _22598_ (.A(net4226),
    .B(_02569_),
    .Y(_02574_));
 sky130_fd_sc_hd__or2_1 _22599_ (.A(net4226),
    .B(_02569_),
    .X(_02575_));
 sky130_fd_sc_hd__a32o_1 _22600_ (.A1(net2042),
    .A2(_02574_),
    .A3(_02575_),
    .B1(net2459),
    .B2(\pid_d.curr_error[8] ),
    .X(_00559_));
 sky130_fd_sc_hd__or2_2 _22601_ (.A(net7265),
    .B(_02574_),
    .X(_02576_));
 sky130_fd_sc_hd__nand2_1 _22602_ (.A(net7265),
    .B(_02574_),
    .Y(_02577_));
 sky130_fd_sc_hd__and2_1 _22603_ (.A(_02576_),
    .B(_02577_),
    .X(_02578_));
 sky130_fd_sc_hd__a22o_1 _22604_ (.A1(net9013),
    .A2(net2045),
    .B1(net2042),
    .B2(_02578_),
    .X(_00560_));
 sky130_fd_sc_hd__nor2_1 _22605_ (.A(net7250),
    .B(_02576_),
    .Y(_02579_));
 sky130_fd_sc_hd__nand2_1 _22606_ (.A(net7250),
    .B(_02576_),
    .Y(_02580_));
 sky130_fd_sc_hd__and3b_1 _22607_ (.A_N(_02579_),
    .B(_02580_),
    .C(net3770),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _22608_ (.A0(\pid_d.curr_error[10] ),
    .A1(net941),
    .S(net3088),
    .X(_02582_));
 sky130_fd_sc_hd__and2_1 _22609_ (.A(net8888),
    .B(_02582_),
    .X(_02583_));
 sky130_fd_sc_hd__clkbuf_1 _22610_ (.A(_02583_),
    .X(_00561_));
 sky130_fd_sc_hd__xnor2_1 _22611_ (.A(net7237),
    .B(_02579_),
    .Y(_02584_));
 sky130_fd_sc_hd__a22o_1 _22612_ (.A1(net9043),
    .A2(_02544_),
    .B1(net2042),
    .B2(_02584_),
    .X(_00562_));
 sky130_fd_sc_hd__o31a_1 _22613_ (.A1(net7250),
    .A2(net7237),
    .A3(_02576_),
    .B1(net7227),
    .X(_02585_));
 sky130_fd_sc_hd__or4_1 _22614_ (.A(net7250),
    .B(net7237),
    .C(net7227),
    .D(_02576_),
    .X(_02586_));
 sky130_fd_sc_hd__and3b_1 _22615_ (.A_N(_02585_),
    .B(net3770),
    .C(_02586_),
    .X(_02587_));
 sky130_fd_sc_hd__mux2_1 _22616_ (.A0(\pid_d.curr_error[12] ),
    .A1(net939),
    .S(net3088),
    .X(_02588_));
 sky130_fd_sc_hd__and2_1 _22617_ (.A(net8888),
    .B(_02588_),
    .X(_02589_));
 sky130_fd_sc_hd__clkbuf_1 _22618_ (.A(_02589_),
    .X(_00563_));
 sky130_fd_sc_hd__or2_1 _22619_ (.A(net7218),
    .B(_02586_),
    .X(_02590_));
 sky130_fd_sc_hd__nand2_1 _22620_ (.A(net7218),
    .B(_02586_),
    .Y(_02591_));
 sky130_fd_sc_hd__and3_1 _22621_ (.A(net3089),
    .B(_02590_),
    .C(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__a22o_1 _22622_ (.A1(net8993),
    .A2(_02544_),
    .B1(_02546_),
    .B2(net858),
    .X(_00564_));
 sky130_fd_sc_hd__or2_1 _22623_ (.A(net7203),
    .B(_02590_),
    .X(_02593_));
 sky130_fd_sc_hd__nand2_1 _22624_ (.A(net7203),
    .B(_02590_),
    .Y(_02594_));
 sky130_fd_sc_hd__and3_1 _22625_ (.A(net3770),
    .B(_02593_),
    .C(_02594_),
    .X(_02595_));
 sky130_fd_sc_hd__mux2_1 _22626_ (.A0(\pid_d.curr_error[14] ),
    .A1(net800),
    .S(_02561_),
    .X(_02596_));
 sky130_fd_sc_hd__and2_1 _22627_ (.A(net8905),
    .B(_02596_),
    .X(_02597_));
 sky130_fd_sc_hd__clkbuf_1 _22628_ (.A(_02597_),
    .X(_00565_));
 sky130_fd_sc_hd__xor2_1 _22629_ (.A(net7192),
    .B(_02593_),
    .X(_02598_));
 sky130_fd_sc_hd__a22o_1 _22630_ (.A1(net9061),
    .A2(_02544_),
    .B1(net2042),
    .B2(_02598_),
    .X(_00566_));
 sky130_fd_sc_hd__buf_1 _22631_ (.A(net3774),
    .X(_02599_));
 sky130_fd_sc_hd__clkbuf_2 _22632_ (.A(_02560_),
    .X(_02600_));
 sky130_fd_sc_hd__a211o_1 _22633_ (.A1(net7368),
    .A2(net3090),
    .B1(net3080),
    .C1(_01245_),
    .X(_02601_));
 sky130_fd_sc_hd__o211a_1 _22634_ (.A1(net5958),
    .A2(net3083),
    .B1(net2456),
    .C1(net8891),
    .X(_00567_));
 sky130_fd_sc_hd__a21o_1 _22635_ (.A1(net3090),
    .A2(_02549_),
    .B1(net3080),
    .X(_02602_));
 sky130_fd_sc_hd__o221a_1 _22636_ (.A1(net5941),
    .A2(net3082),
    .B1(_02602_),
    .B2(_01335_),
    .C1(net8893),
    .X(_00568_));
 sky130_fd_sc_hd__nor2_1 _22637_ (.A(net3081),
    .B(net3092),
    .Y(_02603_));
 sky130_fd_sc_hd__a221oi_1 _22638_ (.A1(net3821),
    .A2(_02600_),
    .B1(net2455),
    .B2(net2070),
    .C1(net3717),
    .Y(_00569_));
 sky130_fd_sc_hd__clkbuf_1 _22639_ (.A(net3767),
    .X(_02604_));
 sky130_fd_sc_hd__nand2_1 _22640_ (.A(net3114),
    .B(net3076),
    .Y(_02605_));
 sky130_fd_sc_hd__o311a_1 _22641_ (.A1(net1724),
    .A2(net3076),
    .A3(net2457),
    .B1(_02605_),
    .C1(net8891),
    .X(_00570_));
 sky130_fd_sc_hd__or2_1 _22642_ (.A(net5860),
    .B(net3083),
    .X(_02606_));
 sky130_fd_sc_hd__o311a_1 _22643_ (.A1(_01642_),
    .A2(net3076),
    .A3(net2040),
    .B1(_02606_),
    .C1(net8891),
    .X(_00571_));
 sky130_fd_sc_hd__a31o_1 _22644_ (.A1(net3090),
    .A2(_02564_),
    .A3(_02565_),
    .B1(net3080),
    .X(_02607_));
 sky130_fd_sc_hd__o221a_1 _22645_ (.A1(net5840),
    .A2(net3082),
    .B1(_02607_),
    .B2(net946),
    .C1(net8893),
    .X(_00572_));
 sky130_fd_sc_hd__nand2_1 _22646_ (.A(_01863_),
    .B(net3077),
    .Y(_02608_));
 sky130_fd_sc_hd__o311a_1 _22647_ (.A1(net805),
    .A2(net3077),
    .A3(net1697),
    .B1(_02608_),
    .C1(net8892),
    .X(_00573_));
 sky130_fd_sc_hd__nand2_1 _22648_ (.A(_00882_),
    .B(net3077),
    .Y(_02609_));
 sky130_fd_sc_hd__o311a_1 _22649_ (.A1(net700),
    .A2(net3077),
    .A3(net1388),
    .B1(_02609_),
    .C1(net8889),
    .X(_00574_));
 sky130_fd_sc_hd__a31o_1 _22650_ (.A1(_02553_),
    .A2(_02574_),
    .A3(_02575_),
    .B1(net3081),
    .X(_02610_));
 sky130_fd_sc_hd__o221a_1 _22651_ (.A1(net9154),
    .A2(net3086),
    .B1(_02610_),
    .B2(_02014_),
    .C1(net8901),
    .X(_00575_));
 sky130_fd_sc_hd__a21o_1 _22652_ (.A1(_02553_),
    .A2(_02578_),
    .B1(net3081),
    .X(_02611_));
 sky130_fd_sc_hd__o221a_1 _22653_ (.A1(net9171),
    .A2(net3086),
    .B1(_02611_),
    .B2(net522),
    .C1(net8894),
    .X(_00576_));
 sky130_fd_sc_hd__or2_1 _22654_ (.A(net5751),
    .B(net3085),
    .X(_02612_));
 sky130_fd_sc_hd__o311a_1 _22655_ (.A1(_02180_),
    .A2(net3078),
    .A3(net941),
    .B1(_02612_),
    .C1(net8889),
    .X(_00577_));
 sky130_fd_sc_hd__a21o_1 _22656_ (.A1(net3089),
    .A2(_02584_),
    .B1(_02600_),
    .X(_02613_));
 sky130_fd_sc_hd__o221a_1 _22657_ (.A1(net9156),
    .A2(_02599_),
    .B1(_02613_),
    .B2(net337),
    .C1(net8890),
    .X(_00578_));
 sky130_fd_sc_hd__a211o_1 _22658_ (.A1(net4364),
    .A2(_02268_),
    .B1(_02600_),
    .C1(net940),
    .X(_02614_));
 sky130_fd_sc_hd__o211a_1 _22659_ (.A1(net5712),
    .A2(net3085),
    .B1(net294),
    .C1(net8888),
    .X(_00579_));
 sky130_fd_sc_hd__or2_1 _22660_ (.A(\pid_d.mult0.b[13] ),
    .B(net3775),
    .X(_02615_));
 sky130_fd_sc_hd__o311a_1 _22661_ (.A1(_02395_),
    .A2(net3079),
    .A3(net856),
    .B1(_02615_),
    .C1(net8905),
    .X(_00580_));
 sky130_fd_sc_hd__or2_1 _22662_ (.A(\pid_d.mult0.b[14] ),
    .B(net3775),
    .X(_02616_));
 sky130_fd_sc_hd__o311a_1 _22663_ (.A1(_02407_),
    .A2(net3079),
    .A3(net800),
    .B1(_02616_),
    .C1(net8905),
    .X(_00581_));
 sky130_fd_sc_hd__a21oi_1 _22664_ (.A1(net3089),
    .A2(_02598_),
    .B1(_02600_),
    .Y(_02617_));
 sky130_fd_sc_hd__o21ai_1 _22665_ (.A1(net4301),
    .A2(_02463_),
    .B1(_02617_),
    .Y(_02618_));
 sky130_fd_sc_hd__o211a_1 _22666_ (.A1(net5650),
    .A2(net3085),
    .B1(net178),
    .C1(net8888),
    .X(_00582_));
 sky130_fd_sc_hd__a22o_1 _22667_ (.A1(\pid_d.ki[0] ),
    .A2(net3010),
    .B1(net2994),
    .B2(\pid_d.kp[0] ),
    .X(_02619_));
 sky130_fd_sc_hd__clkbuf_1 _22668_ (.A(net3098),
    .X(_02620_));
 sky130_fd_sc_hd__mux2_1 _22669_ (.A0(_02619_),
    .A1(net5644),
    .S(net2448),
    .X(_02621_));
 sky130_fd_sc_hd__clkbuf_1 _22670_ (.A(_02621_),
    .X(_00583_));
 sky130_fd_sc_hd__a22o_1 _22671_ (.A1(\pid_d.ki[1] ),
    .A2(net3010),
    .B1(net2994),
    .B2(\pid_d.kp[1] ),
    .X(_02622_));
 sky130_fd_sc_hd__mux2_1 _22672_ (.A0(_02622_),
    .A1(net5630),
    .S(net2448),
    .X(_02623_));
 sky130_fd_sc_hd__clkbuf_1 _22673_ (.A(_02623_),
    .X(_00584_));
 sky130_fd_sc_hd__clkbuf_1 _22674_ (.A(net3705),
    .X(_02624_));
 sky130_fd_sc_hd__a22o_1 _22675_ (.A1(\pid_d.ki[2] ),
    .A2(net2439),
    .B1(net2994),
    .B2(\pid_d.kp[2] ),
    .X(_02625_));
 sky130_fd_sc_hd__mux2_1 _22676_ (.A0(_02625_),
    .A1(net5620),
    .S(net2448),
    .X(_02626_));
 sky130_fd_sc_hd__clkbuf_1 _22677_ (.A(_02626_),
    .X(_00585_));
 sky130_fd_sc_hd__a22o_1 _22678_ (.A1(\pid_d.ki[3] ),
    .A2(net2439),
    .B1(net2994),
    .B2(\pid_d.kp[3] ),
    .X(_02627_));
 sky130_fd_sc_hd__mux2_1 _22679_ (.A0(_02627_),
    .A1(net5606),
    .S(net2448),
    .X(_02628_));
 sky130_fd_sc_hd__clkbuf_1 _22680_ (.A(_02628_),
    .X(_00586_));
 sky130_fd_sc_hd__a22o_1 _22681_ (.A1(\pid_d.ki[4] ),
    .A2(net2439),
    .B1(net2994),
    .B2(\pid_d.kp[4] ),
    .X(_02629_));
 sky130_fd_sc_hd__mux2_1 _22682_ (.A0(_02629_),
    .A1(net5580),
    .S(net2448),
    .X(_02630_));
 sky130_fd_sc_hd__clkbuf_1 _22683_ (.A(_02630_),
    .X(_00587_));
 sky130_fd_sc_hd__a22o_1 _22684_ (.A1(\pid_d.ki[5] ),
    .A2(net2439),
    .B1(net2993),
    .B2(\pid_d.kp[5] ),
    .X(_02631_));
 sky130_fd_sc_hd__mux2_1 _22685_ (.A0(_02631_),
    .A1(net5563),
    .S(net2447),
    .X(_02632_));
 sky130_fd_sc_hd__clkbuf_1 _22686_ (.A(_02632_),
    .X(_00588_));
 sky130_fd_sc_hd__a22o_1 _22687_ (.A1(\pid_d.ki[6] ),
    .A2(net2440),
    .B1(net2993),
    .B2(\pid_d.kp[6] ),
    .X(_02633_));
 sky130_fd_sc_hd__mux2_1 _22688_ (.A0(_02633_),
    .A1(net5548),
    .S(net2447),
    .X(_02634_));
 sky130_fd_sc_hd__clkbuf_1 _22689_ (.A(_02634_),
    .X(_00589_));
 sky130_fd_sc_hd__a22o_1 _22690_ (.A1(\pid_d.ki[7] ),
    .A2(net2440),
    .B1(net2993),
    .B2(\pid_d.kp[7] ),
    .X(_02635_));
 sky130_fd_sc_hd__mux2_1 _22691_ (.A0(_02635_),
    .A1(net5532),
    .S(net2447),
    .X(_02636_));
 sky130_fd_sc_hd__clkbuf_1 _22692_ (.A(_02636_),
    .X(_00590_));
 sky130_fd_sc_hd__a22o_1 _22693_ (.A1(\pid_d.ki[8] ),
    .A2(net2445),
    .B1(net3000),
    .B2(\pid_d.kp[8] ),
    .X(_02637_));
 sky130_fd_sc_hd__mux2_1 _22694_ (.A0(_02637_),
    .A1(net5512),
    .S(net2451),
    .X(_02638_));
 sky130_fd_sc_hd__clkbuf_1 _22695_ (.A(_02638_),
    .X(_00591_));
 sky130_fd_sc_hd__a22o_1 _22696_ (.A1(\pid_d.ki[9] ),
    .A2(net2446),
    .B1(net3696),
    .B2(\pid_d.kp[9] ),
    .X(_02639_));
 sky130_fd_sc_hd__mux2_1 _22697_ (.A0(_02639_),
    .A1(net5496),
    .S(net2451),
    .X(_02640_));
 sky130_fd_sc_hd__clkbuf_1 _22698_ (.A(_02640_),
    .X(_00592_));
 sky130_fd_sc_hd__a22o_1 _22699_ (.A1(\pid_d.ki[10] ),
    .A2(net2446),
    .B1(net3696),
    .B2(\pid_d.kp[10] ),
    .X(_02641_));
 sky130_fd_sc_hd__mux2_1 _22700_ (.A0(_02641_),
    .A1(net5478),
    .S(net3095),
    .X(_02642_));
 sky130_fd_sc_hd__clkbuf_1 _22701_ (.A(_02642_),
    .X(_00593_));
 sky130_fd_sc_hd__a22o_1 _22702_ (.A1(\pid_d.ki[11] ),
    .A2(net2446),
    .B1(net3696),
    .B2(\pid_d.kp[11] ),
    .X(_02643_));
 sky130_fd_sc_hd__mux2_1 _22703_ (.A0(_02643_),
    .A1(net5459),
    .S(net3095),
    .X(_02644_));
 sky130_fd_sc_hd__clkbuf_1 _22704_ (.A(_02644_),
    .X(_00594_));
 sky130_fd_sc_hd__a22o_1 _22705_ (.A1(\pid_d.ki[12] ),
    .A2(net3705),
    .B1(_04886_),
    .B2(\pid_d.kp[12] ),
    .X(_02645_));
 sky130_fd_sc_hd__mux2_1 _22706_ (.A0(_02645_),
    .A1(net5436),
    .S(net3094),
    .X(_02646_));
 sky130_fd_sc_hd__clkbuf_1 _22707_ (.A(_02646_),
    .X(_00595_));
 sky130_fd_sc_hd__a22o_1 _22708_ (.A1(\pid_d.ki[13] ),
    .A2(net3705),
    .B1(_04886_),
    .B2(\pid_d.kp[13] ),
    .X(_02647_));
 sky130_fd_sc_hd__mux2_1 _22709_ (.A0(_02647_),
    .A1(\pid_d.mult0.a[13] ),
    .S(net3094),
    .X(_02648_));
 sky130_fd_sc_hd__clkbuf_1 _22710_ (.A(_02648_),
    .X(_00596_));
 sky130_fd_sc_hd__a22o_1 _22711_ (.A1(\pid_d.ki[14] ),
    .A2(net3705),
    .B1(_04886_),
    .B2(\pid_d.kp[14] ),
    .X(_02649_));
 sky130_fd_sc_hd__mux2_1 _22712_ (.A0(_02649_),
    .A1(net5391),
    .S(net3094),
    .X(_02650_));
 sky130_fd_sc_hd__clkbuf_1 _22713_ (.A(_02650_),
    .X(_00597_));
 sky130_fd_sc_hd__a22o_1 _22714_ (.A1(net5373),
    .A2(net3705),
    .B1(_04886_),
    .B2(net5372),
    .X(_02651_));
 sky130_fd_sc_hd__mux2_1 _22715_ (.A0(_02651_),
    .A1(net5374),
    .S(net3094),
    .X(_02652_));
 sky130_fd_sc_hd__clkbuf_1 _22716_ (.A(_02652_),
    .X(_00598_));
 sky130_fd_sc_hd__and2_1 _22717_ (.A(net3718),
    .B(net97),
    .X(_02653_));
 sky130_fd_sc_hd__inv_2 _22718_ (.A(net8108),
    .Y(_02654_));
 sky130_fd_sc_hd__or4_1 _22719_ (.A(net8096),
    .B(net8098),
    .C(net8106),
    .D(net86),
    .X(_02655_));
 sky130_fd_sc_hd__or4_1 _22720_ (.A(net8107),
    .B(net8105),
    .C(net84),
    .D(net8103),
    .X(_02656_));
 sky130_fd_sc_hd__or4_1 _22721_ (.A(net8921),
    .B(net8102),
    .C(net90),
    .D(net93),
    .X(_02657_));
 sky130_fd_sc_hd__or4_1 _22722_ (.A(net8101),
    .B(net92),
    .C(net8099),
    .D(net94),
    .X(_02658_));
 sky130_fd_sc_hd__or4_1 _22723_ (.A(_02655_),
    .B(_02656_),
    .C(net8084),
    .D(_02658_),
    .X(_02659_));
 sky130_fd_sc_hd__or4_1 _22724_ (.A(_04865_),
    .B(net4366),
    .C(net4327),
    .D(net3102),
    .X(_02660_));
 sky130_fd_sc_hd__o21ai_1 _22725_ (.A1(_02654_),
    .A2(net3764),
    .B1(net2434),
    .Y(_02661_));
 sky130_fd_sc_hd__clkbuf_1 _22726_ (.A(net2037),
    .X(_02662_));
 sky130_fd_sc_hd__mux2_1 _22727_ (.A0(\pid_d.ki[0] ),
    .A1(_02653_),
    .S(net1688),
    .X(_02663_));
 sky130_fd_sc_hd__clkbuf_1 _22728_ (.A(_02663_),
    .X(_00599_));
 sky130_fd_sc_hd__and2_1 _22729_ (.A(net3718),
    .B(net104),
    .X(_02664_));
 sky130_fd_sc_hd__mux2_1 _22730_ (.A0(\pid_d.ki[1] ),
    .A1(_02664_),
    .S(net1688),
    .X(_02665_));
 sky130_fd_sc_hd__clkbuf_1 _22731_ (.A(_02665_),
    .X(_00600_));
 sky130_fd_sc_hd__and2_1 _22732_ (.A(net3718),
    .B(net105),
    .X(_02666_));
 sky130_fd_sc_hd__mux2_1 _22733_ (.A0(\pid_d.ki[2] ),
    .A1(_02666_),
    .S(net1688),
    .X(_02667_));
 sky130_fd_sc_hd__clkbuf_1 _22734_ (.A(_02667_),
    .X(_00601_));
 sky130_fd_sc_hd__and2_1 _22735_ (.A(net3718),
    .B(net106),
    .X(_02668_));
 sky130_fd_sc_hd__mux2_1 _22736_ (.A0(\pid_d.ki[3] ),
    .A1(_02668_),
    .S(net1688),
    .X(_02669_));
 sky130_fd_sc_hd__clkbuf_1 _22737_ (.A(_02669_),
    .X(_00602_));
 sky130_fd_sc_hd__and2_1 _22738_ (.A(net3718),
    .B(net107),
    .X(_02670_));
 sky130_fd_sc_hd__mux2_1 _22739_ (.A0(\pid_d.ki[4] ),
    .A1(_02670_),
    .S(net1689),
    .X(_02671_));
 sky130_fd_sc_hd__clkbuf_1 _22740_ (.A(_02671_),
    .X(_00603_));
 sky130_fd_sc_hd__and2_1 _22741_ (.A(net3719),
    .B(net108),
    .X(_02672_));
 sky130_fd_sc_hd__mux2_1 _22742_ (.A0(\pid_d.ki[5] ),
    .A1(_02672_),
    .S(net1689),
    .X(_02673_));
 sky130_fd_sc_hd__clkbuf_1 _22743_ (.A(_02673_),
    .X(_00604_));
 sky130_fd_sc_hd__and2_1 _22744_ (.A(net3719),
    .B(net109),
    .X(_02674_));
 sky130_fd_sc_hd__mux2_1 _22745_ (.A0(\pid_d.ki[6] ),
    .A1(_02674_),
    .S(net1689),
    .X(_02675_));
 sky130_fd_sc_hd__clkbuf_1 _22746_ (.A(_02675_),
    .X(_00605_));
 sky130_fd_sc_hd__and2_1 _22747_ (.A(net3719),
    .B(net110),
    .X(_02676_));
 sky130_fd_sc_hd__mux2_1 _22748_ (.A0(net9234),
    .A1(_02676_),
    .S(net1690),
    .X(_02677_));
 sky130_fd_sc_hd__clkbuf_1 _22749_ (.A(_02677_),
    .X(_00606_));
 sky130_fd_sc_hd__and2_1 _22750_ (.A(net4304),
    .B(net8928),
    .X(_02678_));
 sky130_fd_sc_hd__mux2_1 _22751_ (.A0(\pid_d.ki[8] ),
    .A1(net3072),
    .S(net1696),
    .X(_02679_));
 sky130_fd_sc_hd__clkbuf_1 _22752_ (.A(_02679_),
    .X(_00607_));
 sky130_fd_sc_hd__and2_1 _22753_ (.A(net4303),
    .B(net8924),
    .X(_02680_));
 sky130_fd_sc_hd__mux2_1 _22754_ (.A0(\pid_d.ki[9] ),
    .A1(net3070),
    .S(net1696),
    .X(_02681_));
 sky130_fd_sc_hd__clkbuf_1 _22755_ (.A(_02681_),
    .X(_00608_));
 sky130_fd_sc_hd__and2_1 _22756_ (.A(net4303),
    .B(net8092),
    .X(_02682_));
 sky130_fd_sc_hd__mux2_1 _22757_ (.A0(\pid_d.ki[10] ),
    .A1(net3069),
    .S(net2037),
    .X(_02683_));
 sky130_fd_sc_hd__clkbuf_1 _22758_ (.A(_02683_),
    .X(_00609_));
 sky130_fd_sc_hd__and2_1 _22759_ (.A(net4302),
    .B(net8086),
    .X(_02684_));
 sky130_fd_sc_hd__mux2_1 _22760_ (.A0(\pid_d.ki[11] ),
    .A1(net3068),
    .S(net2037),
    .X(_02685_));
 sky130_fd_sc_hd__clkbuf_1 _22761_ (.A(_02685_),
    .X(_00610_));
 sky130_fd_sc_hd__and2_1 _22762_ (.A(net4303),
    .B(net8946),
    .X(_02686_));
 sky130_fd_sc_hd__mux2_1 _22763_ (.A0(\pid_d.ki[12] ),
    .A1(_02686_),
    .S(net2038),
    .X(_02687_));
 sky130_fd_sc_hd__clkbuf_1 _22764_ (.A(_02687_),
    .X(_00611_));
 sky130_fd_sc_hd__and2_1 _22765_ (.A(net4302),
    .B(net8940),
    .X(_02688_));
 sky130_fd_sc_hd__mux2_1 _22766_ (.A0(\pid_d.ki[13] ),
    .A1(_02688_),
    .S(net2038),
    .X(_02689_));
 sky130_fd_sc_hd__clkbuf_1 _22767_ (.A(_02689_),
    .X(_00612_));
 sky130_fd_sc_hd__and2_1 _22768_ (.A(net4302),
    .B(net8936),
    .X(_02690_));
 sky130_fd_sc_hd__mux2_1 _22769_ (.A0(\pid_d.ki[14] ),
    .A1(_02690_),
    .S(net2039),
    .X(_02691_));
 sky130_fd_sc_hd__clkbuf_1 _22770_ (.A(_02691_),
    .X(_00613_));
 sky130_fd_sc_hd__and2_1 _22771_ (.A(net4302),
    .B(net8932),
    .X(_02692_));
 sky130_fd_sc_hd__mux2_1 _22772_ (.A0(\pid_d.ki[15] ),
    .A1(_02692_),
    .S(net2039),
    .X(_02693_));
 sky130_fd_sc_hd__clkbuf_1 _22773_ (.A(_02693_),
    .X(_00614_));
 sky130_fd_sc_hd__o21ai_1 _22774_ (.A1(net8108),
    .A2(net3764),
    .B1(net2434),
    .Y(_02694_));
 sky130_fd_sc_hd__clkbuf_1 _22775_ (.A(net2035),
    .X(_02695_));
 sky130_fd_sc_hd__mux2_1 _22776_ (.A0(\pid_d.kp[0] ),
    .A1(_02653_),
    .S(net1679),
    .X(_02696_));
 sky130_fd_sc_hd__clkbuf_1 _22777_ (.A(_02696_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _22778_ (.A0(\pid_d.kp[1] ),
    .A1(_02664_),
    .S(net1679),
    .X(_02697_));
 sky130_fd_sc_hd__clkbuf_1 _22779_ (.A(_02697_),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _22780_ (.A0(\pid_d.kp[2] ),
    .A1(_02666_),
    .S(net1680),
    .X(_02698_));
 sky130_fd_sc_hd__clkbuf_1 _22781_ (.A(_02698_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _22782_ (.A0(\pid_d.kp[3] ),
    .A1(_02668_),
    .S(net1679),
    .X(_02699_));
 sky130_fd_sc_hd__clkbuf_1 _22783_ (.A(_02699_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _22784_ (.A0(\pid_d.kp[4] ),
    .A1(_02670_),
    .S(net1680),
    .X(_02700_));
 sky130_fd_sc_hd__clkbuf_1 _22785_ (.A(_02700_),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _22786_ (.A0(\pid_d.kp[5] ),
    .A1(_02672_),
    .S(net1680),
    .X(_02701_));
 sky130_fd_sc_hd__clkbuf_1 _22787_ (.A(_02701_),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _22788_ (.A0(\pid_d.kp[6] ),
    .A1(_02674_),
    .S(net1681),
    .X(_02702_));
 sky130_fd_sc_hd__clkbuf_1 _22789_ (.A(_02702_),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _22790_ (.A0(\pid_d.kp[7] ),
    .A1(_02676_),
    .S(net1681),
    .X(_02703_));
 sky130_fd_sc_hd__clkbuf_1 _22791_ (.A(_02703_),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _22792_ (.A0(\pid_d.kp[8] ),
    .A1(net3072),
    .S(net1687),
    .X(_02704_));
 sky130_fd_sc_hd__clkbuf_1 _22793_ (.A(_02704_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _22794_ (.A0(\pid_d.kp[9] ),
    .A1(net3070),
    .S(net1687),
    .X(_02705_));
 sky130_fd_sc_hd__clkbuf_1 _22795_ (.A(_02705_),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _22796_ (.A0(\pid_d.kp[10] ),
    .A1(net3069),
    .S(net2035),
    .X(_02706_));
 sky130_fd_sc_hd__clkbuf_1 _22797_ (.A(_02706_),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _22798_ (.A0(\pid_d.kp[11] ),
    .A1(net3068),
    .S(net2035),
    .X(_02707_));
 sky130_fd_sc_hd__clkbuf_1 _22799_ (.A(_02707_),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_1 _22800_ (.A0(\pid_d.kp[12] ),
    .A1(_02686_),
    .S(_02694_),
    .X(_02708_));
 sky130_fd_sc_hd__clkbuf_1 _22801_ (.A(_02708_),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _22802_ (.A0(\pid_d.kp[13] ),
    .A1(_02688_),
    .S(net2036),
    .X(_02709_));
 sky130_fd_sc_hd__clkbuf_1 _22803_ (.A(_02709_),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _22804_ (.A0(\pid_d.kp[14] ),
    .A1(_02690_),
    .S(net2036),
    .X(_02710_));
 sky130_fd_sc_hd__clkbuf_1 _22805_ (.A(_02710_),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _22806_ (.A0(\pid_d.kp[15] ),
    .A1(_02692_),
    .S(net2036),
    .X(_02711_));
 sky130_fd_sc_hd__clkbuf_1 _22807_ (.A(_02711_),
    .X(_00630_));
 sky130_fd_sc_hd__or4_1 _22808_ (.A(net4381),
    .B(net4317),
    .C(net4350),
    .D(net4373),
    .X(_02712_));
 sky130_fd_sc_hd__mux2_1 _22809_ (.A0(net4328),
    .A1(\pid_d.out_valid ),
    .S(net3763),
    .X(_02713_));
 sky130_fd_sc_hd__and2_1 _22810_ (.A(net8895),
    .B(_02713_),
    .X(_02714_));
 sky130_fd_sc_hd__clkbuf_1 _22811_ (.A(_02714_),
    .X(_00631_));
 sky130_fd_sc_hd__nor2_1 _22812_ (.A(net4299),
    .B(net2464),
    .Y(_02715_));
 sky130_fd_sc_hd__nor4_1 _22813_ (.A(net4389),
    .B(net4382),
    .C(net4321),
    .D(net4351),
    .Y(_02716_));
 sky130_fd_sc_hd__nand2_1 _22814_ (.A(net5986),
    .B(net3759),
    .Y(_02717_));
 sky130_fd_sc_hd__mux2_1 _22815_ (.A0(_02717_),
    .A1(net5986),
    .S(\pid_d.out[0] ),
    .X(_02718_));
 sky130_fd_sc_hd__and2b_1 _22816_ (.A_N(_02718_),
    .B(net4336),
    .X(_02719_));
 sky130_fd_sc_hd__a221o_1 _22817_ (.A1(\pid_d.out[0] ),
    .A2(net2463),
    .B1(net2034),
    .B2(net479),
    .C1(_02719_),
    .X(_02720_));
 sky130_fd_sc_hd__and2_1 _22818_ (.A(net8896),
    .B(_02720_),
    .X(_02721_));
 sky130_fd_sc_hd__clkbuf_1 _22819_ (.A(_02721_),
    .X(_00632_));
 sky130_fd_sc_hd__clkbuf_1 _22820_ (.A(net3759),
    .X(_02722_));
 sky130_fd_sc_hd__nand2_1 _22821_ (.A(\pid_d.out[0] ),
    .B(net5986),
    .Y(_02723_));
 sky130_fd_sc_hd__xor2_1 _22822_ (.A(net5366),
    .B(net5984),
    .X(_02724_));
 sky130_fd_sc_hd__xnor2_1 _22823_ (.A(_02723_),
    .B(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__a221o_1 _22824_ (.A1(net4360),
    .A2(net560),
    .B1(_02725_),
    .B2(net4335),
    .C1(net2463),
    .X(_02726_));
 sky130_fd_sc_hd__o211a_1 _22825_ (.A1(net5366),
    .A2(net3065),
    .B1(_02726_),
    .C1(net8897),
    .X(_00633_));
 sky130_fd_sc_hd__nand2_1 _22826_ (.A(net5366),
    .B(net5984),
    .Y(_02727_));
 sky130_fd_sc_hd__o211ai_2 _22827_ (.A1(net5366),
    .A2(net5984),
    .B1(net5986),
    .C1(\pid_d.out[0] ),
    .Y(_02728_));
 sky130_fd_sc_hd__nand2_1 _22828_ (.A(_02727_),
    .B(_02728_),
    .Y(_02729_));
 sky130_fd_sc_hd__xnor2_1 _22829_ (.A(net5365),
    .B(net5983),
    .Y(_02730_));
 sky130_fd_sc_hd__xnor2_1 _22830_ (.A(_02729_),
    .B(_02730_),
    .Y(_02731_));
 sky130_fd_sc_hd__a221o_1 _22831_ (.A1(net4354),
    .A2(net553),
    .B1(_02731_),
    .B2(net4335),
    .C1(net2463),
    .X(_02732_));
 sky130_fd_sc_hd__o211a_1 _22832_ (.A1(net5365),
    .A2(net3065),
    .B1(_02732_),
    .C1(net8897),
    .X(_00634_));
 sky130_fd_sc_hd__inv_2 _22833_ (.A(net5983),
    .Y(_02733_));
 sky130_fd_sc_hd__a21o_1 _22834_ (.A1(_02727_),
    .A2(_02728_),
    .B1(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__inv_2 _22835_ (.A(net5365),
    .Y(_02735_));
 sky130_fd_sc_hd__a31o_1 _22836_ (.A1(_02733_),
    .A2(_02727_),
    .A3(_02728_),
    .B1(_02735_),
    .X(_02736_));
 sky130_fd_sc_hd__and2_1 _22837_ (.A(_02734_),
    .B(_02736_),
    .X(_02737_));
 sky130_fd_sc_hd__xnor2_1 _22838_ (.A(\pid_d.out[3] ),
    .B(net5982),
    .Y(_02738_));
 sky130_fd_sc_hd__nand2_1 _22839_ (.A(_02737_),
    .B(_02738_),
    .Y(_02739_));
 sky130_fd_sc_hd__or2_1 _22840_ (.A(_02737_),
    .B(_02738_),
    .X(_02740_));
 sky130_fd_sc_hd__a32o_1 _22841_ (.A1(net4335),
    .A2(_02739_),
    .A3(_02740_),
    .B1(net415),
    .B2(net4354),
    .X(_02741_));
 sky130_fd_sc_hd__mux2_1 _22842_ (.A0(\pid_d.out[3] ),
    .A1(_02741_),
    .S(net3065),
    .X(_02742_));
 sky130_fd_sc_hd__and2_1 _22843_ (.A(net8897),
    .B(_02742_),
    .X(_02743_));
 sky130_fd_sc_hd__clkbuf_1 _22844_ (.A(_02743_),
    .X(_00635_));
 sky130_fd_sc_hd__inv_2 _22845_ (.A(net5982),
    .Y(_02744_));
 sky130_fd_sc_hd__inv_2 _22846_ (.A(\pid_d.out[3] ),
    .Y(_02745_));
 sky130_fd_sc_hd__a31o_1 _22847_ (.A1(_02744_),
    .A2(_02734_),
    .A3(_02736_),
    .B1(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__o21ai_4 _22848_ (.A1(_02744_),
    .A2(_02737_),
    .B1(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__xnor2_1 _22849_ (.A(\pid_d.out[4] ),
    .B(net5981),
    .Y(_02748_));
 sky130_fd_sc_hd__xnor2_1 _22850_ (.A(_02747_),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__a221o_1 _22851_ (.A1(net4360),
    .A2(net475),
    .B1(_02749_),
    .B2(net4336),
    .C1(net2465),
    .X(_02750_));
 sky130_fd_sc_hd__o211a_1 _22852_ (.A1(\pid_d.out[4] ),
    .A2(net3065),
    .B1(_02750_),
    .C1(net8897),
    .X(_00636_));
 sky130_fd_sc_hd__a21o_1 _22853_ (.A1(net5981),
    .A2(_02747_),
    .B1(\pid_d.out[4] ),
    .X(_02751_));
 sky130_fd_sc_hd__o21a_1 _22854_ (.A1(net5981),
    .A2(_02747_),
    .B1(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__xor2_1 _22855_ (.A(net5364),
    .B(net5980),
    .X(_02753_));
 sky130_fd_sc_hd__or2_1 _22856_ (.A(_02752_),
    .B(_02753_),
    .X(_02754_));
 sky130_fd_sc_hd__nand2_1 _22857_ (.A(_02752_),
    .B(_02753_),
    .Y(_02755_));
 sky130_fd_sc_hd__a32o_1 _22858_ (.A1(net4337),
    .A2(_02754_),
    .A3(_02755_),
    .B1(net523),
    .B2(net4359),
    .X(_02756_));
 sky130_fd_sc_hd__mux2_1 _22859_ (.A0(net5364),
    .A1(_02756_),
    .S(net3066),
    .X(_02757_));
 sky130_fd_sc_hd__and2_1 _22860_ (.A(net8897),
    .B(_02757_),
    .X(_02758_));
 sky130_fd_sc_hd__clkbuf_1 _22861_ (.A(_02758_),
    .X(_00637_));
 sky130_fd_sc_hd__o21a_1 _22862_ (.A1(net5981),
    .A2(_02747_),
    .B1(\pid_d.out[4] ),
    .X(_02759_));
 sky130_fd_sc_hd__a211o_1 _22863_ (.A1(net5981),
    .A2(_02747_),
    .B1(_02759_),
    .C1(net5980),
    .X(_02760_));
 sky130_fd_sc_hd__o211a_1 _22864_ (.A1(net5981),
    .A2(_02747_),
    .B1(_02751_),
    .C1(net5980),
    .X(_02761_));
 sky130_fd_sc_hd__a21oi_2 _22865_ (.A1(net5364),
    .A2(_02760_),
    .B1(_02761_),
    .Y(_02762_));
 sky130_fd_sc_hd__xnor2_1 _22866_ (.A(net5363),
    .B(net5979),
    .Y(_02763_));
 sky130_fd_sc_hd__nand2_1 _22867_ (.A(_02762_),
    .B(_02763_),
    .Y(_02764_));
 sky130_fd_sc_hd__or2_1 _22868_ (.A(_02762_),
    .B(_02763_),
    .X(_02765_));
 sky130_fd_sc_hd__a32o_1 _22869_ (.A1(net4337),
    .A2(_02764_),
    .A3(_02765_),
    .B1(net472),
    .B2(net4359),
    .X(_02766_));
 sky130_fd_sc_hd__mux2_1 _22870_ (.A0(net5363),
    .A1(_02766_),
    .S(net3066),
    .X(_02767_));
 sky130_fd_sc_hd__and2_1 _22871_ (.A(net8898),
    .B(_02767_),
    .X(_02768_));
 sky130_fd_sc_hd__clkbuf_1 _22872_ (.A(_02768_),
    .X(_00638_));
 sky130_fd_sc_hd__o21ba_1 _22873_ (.A1(_01819_),
    .A2(_02762_),
    .B1_N(net5363),
    .X(_02769_));
 sky130_fd_sc_hd__a21o_1 _22874_ (.A1(_01819_),
    .A2(_02762_),
    .B1(_02769_),
    .X(_02770_));
 sky130_fd_sc_hd__xnor2_1 _22875_ (.A(net5360),
    .B(net5978),
    .Y(_02771_));
 sky130_fd_sc_hd__nand2_1 _22876_ (.A(_02770_),
    .B(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__or2_1 _22877_ (.A(_02770_),
    .B(_02771_),
    .X(_02773_));
 sky130_fd_sc_hd__a32o_1 _22878_ (.A1(net4337),
    .A2(_02772_),
    .A3(_02773_),
    .B1(net412),
    .B2(net4359),
    .X(_02774_));
 sky130_fd_sc_hd__mux2_1 _22879_ (.A0(net5360),
    .A1(_02774_),
    .S(net3066),
    .X(_02775_));
 sky130_fd_sc_hd__and2_1 _22880_ (.A(net8898),
    .B(_02775_),
    .X(_02776_));
 sky130_fd_sc_hd__clkbuf_1 _22881_ (.A(_02776_),
    .X(_00639_));
 sky130_fd_sc_hd__nor2_1 _22882_ (.A(net5357),
    .B(net3103),
    .Y(_02777_));
 sky130_fd_sc_hd__o21ba_1 _22883_ (.A1(_01917_),
    .A2(_02770_),
    .B1_N(net5360),
    .X(_02778_));
 sky130_fd_sc_hd__a21o_1 _22884_ (.A1(_01917_),
    .A2(_02770_),
    .B1(_02778_),
    .X(_02779_));
 sky130_fd_sc_hd__xnor2_1 _22885_ (.A(net5977),
    .B(_02779_),
    .Y(_02780_));
 sky130_fd_sc_hd__mux2_1 _22886_ (.A0(net5357),
    .A1(_02777_),
    .S(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__a22o_1 _22887_ (.A1(net5357),
    .A2(net3103),
    .B1(_02781_),
    .B2(net4338),
    .X(_02782_));
 sky130_fd_sc_hd__a21o_1 _22888_ (.A1(net346),
    .A2(net2033),
    .B1(_02782_),
    .X(_02783_));
 sky130_fd_sc_hd__and2_1 _22889_ (.A(net8895),
    .B(_02783_),
    .X(_02784_));
 sky130_fd_sc_hd__clkbuf_1 _22890_ (.A(_02784_),
    .X(_00640_));
 sky130_fd_sc_hd__nor2_1 _22891_ (.A(net5354),
    .B(net3103),
    .Y(_02785_));
 sky130_fd_sc_hd__o21ba_1 _22892_ (.A1(_02017_),
    .A2(_02779_),
    .B1_N(net5357),
    .X(_02786_));
 sky130_fd_sc_hd__a21o_1 _22893_ (.A1(_02017_),
    .A2(_02779_),
    .B1(_02786_),
    .X(_02787_));
 sky130_fd_sc_hd__xnor2_1 _22894_ (.A(net5976),
    .B(_02787_),
    .Y(_02788_));
 sky130_fd_sc_hd__mux2_1 _22895_ (.A0(net5354),
    .A1(_02785_),
    .S(_02788_),
    .X(_02789_));
 sky130_fd_sc_hd__a22o_1 _22896_ (.A1(net5354),
    .A2(net3103),
    .B1(_02789_),
    .B2(net4328),
    .X(_02790_));
 sky130_fd_sc_hd__a21o_1 _22897_ (.A1(net342),
    .A2(net2033),
    .B1(_02790_),
    .X(_02791_));
 sky130_fd_sc_hd__and2_1 _22898_ (.A(net8899),
    .B(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__clkbuf_1 _22899_ (.A(_02792_),
    .X(_00641_));
 sky130_fd_sc_hd__nand2_1 _22900_ (.A(net4370),
    .B(net3761),
    .Y(_02793_));
 sky130_fd_sc_hd__nor2_1 _22901_ (.A(net338),
    .B(_02793_),
    .Y(_02794_));
 sky130_fd_sc_hd__nor2_1 _22902_ (.A(\pid_d.out[10] ),
    .B(net3103),
    .Y(_02795_));
 sky130_fd_sc_hd__o21ba_1 _22903_ (.A1(_02109_),
    .A2(_02787_),
    .B1_N(net5354),
    .X(_02796_));
 sky130_fd_sc_hd__a21o_1 _22904_ (.A1(_02109_),
    .A2(_02787_),
    .B1(_02796_),
    .X(_02797_));
 sky130_fd_sc_hd__xnor2_1 _22905_ (.A(\pid_d.curr_int[10] ),
    .B(_02797_),
    .Y(_02798_));
 sky130_fd_sc_hd__mux2_1 _22906_ (.A0(\pid_d.out[10] ),
    .A1(_02795_),
    .S(_02798_),
    .X(_02799_));
 sky130_fd_sc_hd__a22o_1 _22907_ (.A1(\pid_d.out[10] ),
    .A2(net2466),
    .B1(_02799_),
    .B2(net4329),
    .X(_02800_));
 sky130_fd_sc_hd__o21a_1 _22908_ (.A1(_02794_),
    .A2(_02800_),
    .B1(net8903),
    .X(_00642_));
 sky130_fd_sc_hd__a21bo_1 _22909_ (.A1(_02183_),
    .A2(_02797_),
    .B1_N(\pid_d.out[10] ),
    .X(_02801_));
 sky130_fd_sc_hd__o21a_1 _22910_ (.A1(_02183_),
    .A2(_02797_),
    .B1(_02801_),
    .X(_02802_));
 sky130_fd_sc_hd__xnor2_1 _22911_ (.A(net5340),
    .B(\pid_d.curr_int[11] ),
    .Y(_02803_));
 sky130_fd_sc_hd__nand2_1 _22912_ (.A(_02802_),
    .B(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__or2_1 _22913_ (.A(_02802_),
    .B(_02803_),
    .X(_02805_));
 sky130_fd_sc_hd__a32o_1 _22914_ (.A1(net4333),
    .A2(_02804_),
    .A3(_02805_),
    .B1(net298),
    .B2(net4362),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_1 _22915_ (.A0(net5340),
    .A1(_02806_),
    .S(net3064),
    .X(_02807_));
 sky130_fd_sc_hd__and2_1 _22916_ (.A(net8903),
    .B(_02807_),
    .X(_02808_));
 sky130_fd_sc_hd__clkbuf_1 _22917_ (.A(_02808_),
    .X(_00643_));
 sky130_fd_sc_hd__nor2_1 _22918_ (.A(net5339),
    .B(net3104),
    .Y(_02809_));
 sky130_fd_sc_hd__o21ba_1 _22919_ (.A1(_02270_),
    .A2(_02802_),
    .B1_N(net5340),
    .X(_02810_));
 sky130_fd_sc_hd__a21o_1 _22920_ (.A1(_02270_),
    .A2(_02802_),
    .B1(_02810_),
    .X(_02811_));
 sky130_fd_sc_hd__inv_2 _22921_ (.A(_02811_),
    .Y(_02812_));
 sky130_fd_sc_hd__or2_1 _22922_ (.A(net5975),
    .B(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__nand2_1 _22923_ (.A(net5975),
    .B(_02812_),
    .Y(_02814_));
 sky130_fd_sc_hd__and2_1 _22924_ (.A(_02813_),
    .B(_02814_),
    .X(_02815_));
 sky130_fd_sc_hd__mux2_1 _22925_ (.A0(net5339),
    .A1(_02809_),
    .S(_02815_),
    .X(_02816_));
 sky130_fd_sc_hd__nor2_1 _22926_ (.A(net295),
    .B(_02793_),
    .Y(_02817_));
 sky130_fd_sc_hd__a221o_1 _22927_ (.A1(net5339),
    .A2(net2467),
    .B1(_02816_),
    .B2(net4333),
    .C1(_02817_),
    .X(_02818_));
 sky130_fd_sc_hd__and2_1 _22928_ (.A(net8907),
    .B(_02818_),
    .X(_02819_));
 sky130_fd_sc_hd__clkbuf_1 _22929_ (.A(_02819_),
    .X(_00644_));
 sky130_fd_sc_hd__a21o_1 _22930_ (.A1(net5975),
    .A2(_02812_),
    .B1(net5339),
    .X(_02820_));
 sky130_fd_sc_hd__xor2_1 _22931_ (.A(net5327),
    .B(\pid_d.curr_int[13] ),
    .X(_02821_));
 sky130_fd_sc_hd__a21o_1 _22932_ (.A1(_02813_),
    .A2(_02820_),
    .B1(_02821_),
    .X(_02822_));
 sky130_fd_sc_hd__nand3_1 _22933_ (.A(_02813_),
    .B(_02820_),
    .C(_02821_),
    .Y(_02823_));
 sky130_fd_sc_hd__a32o_1 _22934_ (.A1(net4331),
    .A2(_02822_),
    .A3(_02823_),
    .B1(net271),
    .B2(net4362),
    .X(_02824_));
 sky130_fd_sc_hd__mux2_1 _22935_ (.A0(net5327),
    .A1(_02824_),
    .S(net3064),
    .X(_02825_));
 sky130_fd_sc_hd__and2_1 _22936_ (.A(net8908),
    .B(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__clkbuf_1 _22937_ (.A(_02826_),
    .X(_00645_));
 sky130_fd_sc_hd__and2_1 _22938_ (.A(net205),
    .B(net2030),
    .X(_02827_));
 sky130_fd_sc_hd__nor2_1 _22939_ (.A(\pid_d.out[14] ),
    .B(net3104),
    .Y(_02828_));
 sky130_fd_sc_hd__o211a_1 _22940_ (.A1(net5327),
    .A2(\pid_d.curr_int[13] ),
    .B1(_02813_),
    .C1(_02820_),
    .X(_02829_));
 sky130_fd_sc_hd__a21oi_1 _22941_ (.A1(net5327),
    .A2(\pid_d.curr_int[13] ),
    .B1(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__xnor2_1 _22942_ (.A(\pid_d.curr_int[14] ),
    .B(_02830_),
    .Y(_02831_));
 sky130_fd_sc_hd__mux2_1 _22943_ (.A0(\pid_d.out[14] ),
    .A1(_02828_),
    .S(_02831_),
    .X(_02832_));
 sky130_fd_sc_hd__a22o_1 _22944_ (.A1(\pid_d.out[14] ),
    .A2(net2468),
    .B1(_02832_),
    .B2(net4331),
    .X(_02833_));
 sky130_fd_sc_hd__o21a_1 _22945_ (.A1(_02827_),
    .A2(_02833_),
    .B1(net8904),
    .X(_00646_));
 sky130_fd_sc_hd__o21ba_1 _22946_ (.A1(net551),
    .A2(net549),
    .B1_N(_02324_),
    .X(_02834_));
 sky130_fd_sc_hd__a2bb2o_1 _22947_ (.A1_N(_02388_),
    .A2_N(_02834_),
    .B1(_02455_),
    .B2(net517),
    .X(_02835_));
 sky130_fd_sc_hd__a21o_1 _22948_ (.A1(net551),
    .A2(net549),
    .B1(_02325_),
    .X(_02836_));
 sky130_fd_sc_hd__a21o_1 _22949_ (.A1(_02386_),
    .A2(_02836_),
    .B1(_02515_),
    .X(_02837_));
 sky130_fd_sc_hd__a211o_1 _22950_ (.A1(_02279_),
    .A2(net552),
    .B1(_02514_),
    .C1(net336),
    .X(_02838_));
 sky130_fd_sc_hd__nand2_1 _22951_ (.A(net336),
    .B(_02324_),
    .Y(_02839_));
 sky130_fd_sc_hd__o22a_1 _22952_ (.A1(_02839_),
    .A2(_02515_),
    .B1(_02838_),
    .B2(_02387_),
    .X(_02840_));
 sky130_fd_sc_hd__a21o_1 _22953_ (.A1(_02388_),
    .A2(_02838_),
    .B1(_02840_),
    .X(_02841_));
 sky130_fd_sc_hd__a31o_1 _22954_ (.A1(_02835_),
    .A2(_02837_),
    .A3(_02841_),
    .B1(_02513_),
    .X(_02842_));
 sky130_fd_sc_hd__xnor2_1 _22955_ (.A(net5314),
    .B(net5974),
    .Y(_02843_));
 sky130_fd_sc_hd__nand2_1 _22956_ (.A(\pid_d.out[14] ),
    .B(\pid_d.curr_int[14] ),
    .Y(_02844_));
 sky130_fd_sc_hd__nor2_1 _22957_ (.A(\pid_d.out[14] ),
    .B(\pid_d.curr_int[14] ),
    .Y(_02845_));
 sky130_fd_sc_hd__a21oi_1 _22958_ (.A1(_02830_),
    .A2(_02844_),
    .B1(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__xnor2_1 _22959_ (.A(_02843_),
    .B(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__a221o_1 _22960_ (.A1(net4370),
    .A2(net201),
    .B1(_02847_),
    .B2(net4331),
    .C1(net2467),
    .X(_02848_));
 sky130_fd_sc_hd__o211a_1 _22961_ (.A1(net5314),
    .A2(net3064),
    .B1(_02848_),
    .C1(net8910),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _22962_ (.A0(\matmul0.beta_pass[0] ),
    .A1(net4063),
    .S(net6572),
    .X(_02849_));
 sky130_fd_sc_hd__clkbuf_1 _22963_ (.A(_02849_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _22964_ (.A0(\matmul0.beta_pass[1] ),
    .A1(net3383),
    .S(net6570),
    .X(_02850_));
 sky130_fd_sc_hd__clkbuf_1 _22965_ (.A(_02850_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _22966_ (.A0(\matmul0.beta_pass[2] ),
    .A1(net2613),
    .S(net6569),
    .X(_02851_));
 sky130_fd_sc_hd__clkbuf_1 _22967_ (.A(_02851_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _22968_ (.A0(\matmul0.beta_pass[3] ),
    .A1(net2202),
    .S(net6567),
    .X(_02852_));
 sky130_fd_sc_hd__clkbuf_1 _22969_ (.A(_02852_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _22970_ (.A0(\matmul0.beta_pass[4] ),
    .A1(net1838),
    .S(net6567),
    .X(_02853_));
 sky130_fd_sc_hd__clkbuf_1 _22971_ (.A(_02853_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _22972_ (.A0(net9238),
    .A1(net1240),
    .S(net6570),
    .X(_02854_));
 sky130_fd_sc_hd__clkbuf_1 _22973_ (.A(_02854_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _22974_ (.A0(\matmul0.beta_pass[6] ),
    .A1(net972),
    .S(net6573),
    .X(_02855_));
 sky130_fd_sc_hd__clkbuf_1 _22975_ (.A(_02855_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _22976_ (.A0(\matmul0.beta_pass[7] ),
    .A1(net823),
    .S(net6569),
    .X(_02856_));
 sky130_fd_sc_hd__clkbuf_1 _22977_ (.A(_02856_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _22978_ (.A0(net5243),
    .A1(net720),
    .S(net6571),
    .X(_02857_));
 sky130_fd_sc_hd__clkbuf_1 _22979_ (.A(_02857_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _22980_ (.A0(net5242),
    .A1(net619),
    .S(net6568),
    .X(_02858_));
 sky130_fd_sc_hd__clkbuf_1 _22981_ (.A(_02858_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _22982_ (.A0(net5219),
    .A1(net528),
    .S(net6568),
    .X(_02859_));
 sky130_fd_sc_hd__clkbuf_1 _22983_ (.A(_02859_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _22984_ (.A0(net5218),
    .A1(net423),
    .S(net6568),
    .X(_02860_));
 sky130_fd_sc_hd__clkbuf_1 _22985_ (.A(_02860_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _22986_ (.A0(\matmul0.beta_pass[12] ),
    .A1(net353),
    .S(net6578),
    .X(_02861_));
 sky130_fd_sc_hd__clkbuf_1 _22987_ (.A(_02861_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _22988_ (.A0(net9235),
    .A1(_08738_),
    .S(net6574),
    .X(_02862_));
 sky130_fd_sc_hd__clkbuf_1 _22989_ (.A(_02862_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _22990_ (.A0(\matmul0.beta_pass[14] ),
    .A1(_08744_),
    .S(net6575),
    .X(_02863_));
 sky130_fd_sc_hd__clkbuf_1 _22991_ (.A(_02863_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _22992_ (.A0(\matmul0.beta_pass[15] ),
    .A1(_08750_),
    .S(net6575),
    .X(_02864_));
 sky130_fd_sc_hd__clkbuf_1 _22993_ (.A(_02864_),
    .X(_00663_));
 sky130_fd_sc_hd__nor2_1 _22994_ (.A(net2885),
    .B(_06513_),
    .Y(_02865_));
 sky130_fd_sc_hd__o2bb2a_1 _22995_ (.A1_N(net6447),
    .A2_N(net6445),
    .B1(net9110),
    .B2(_02865_),
    .X(_00664_));
 sky130_fd_sc_hd__o31a_1 _22996_ (.A1(net7470),
    .A2(\pid_q.state[0] ),
    .A3(net7489),
    .B1(net8865),
    .X(_02866_));
 sky130_fd_sc_hd__buf_1 _22997_ (.A(_02866_),
    .X(_02867_));
 sky130_fd_sc_hd__inv_2 _22998_ (.A(net3758),
    .Y(_02868_));
 sky130_fd_sc_hd__o311a_1 _22999_ (.A1(net7524),
    .A2(net7500),
    .A3(net7464),
    .B1(_02868_),
    .C1(net8865),
    .X(_02869_));
 sky130_fd_sc_hd__buf_1 _23000_ (.A(_02869_),
    .X(_02870_));
 sky130_fd_sc_hd__nand2_2 _23001_ (.A(net5016),
    .B(net4685),
    .Y(_02871_));
 sky130_fd_sc_hd__nand2_1 _23002_ (.A(net5069),
    .B(net4629),
    .Y(_02872_));
 sky130_fd_sc_hd__nand2_1 _23003_ (.A(net5044),
    .B(net4654),
    .Y(_02873_));
 sky130_fd_sc_hd__xor2_1 _23004_ (.A(_02872_),
    .B(_02873_),
    .X(_02874_));
 sky130_fd_sc_hd__xnor2_2 _23005_ (.A(_02871_),
    .B(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__nand2_1 _23006_ (.A(net5086),
    .B(net4613),
    .Y(_02876_));
 sky130_fd_sc_hd__nand2_1 _23007_ (.A(net5141),
    .B(net4571),
    .Y(_02877_));
 sky130_fd_sc_hd__nand2_1 _23008_ (.A(net5133),
    .B(net4595),
    .Y(_02878_));
 sky130_fd_sc_hd__xnor2_1 _23009_ (.A(_02877_),
    .B(_02878_),
    .Y(_02879_));
 sky130_fd_sc_hd__xnor2_1 _23010_ (.A(_02876_),
    .B(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__nand2_1 _23011_ (.A(net5087),
    .B(net4623),
    .Y(_02881_));
 sky130_fd_sc_hd__nand2_1 _23012_ (.A(net5132),
    .B(net4610),
    .Y(_02882_));
 sky130_fd_sc_hd__nand2_1 _23013_ (.A(net5141),
    .B(net4595),
    .Y(_02883_));
 sky130_fd_sc_hd__o21a_1 _23014_ (.A1(_02881_),
    .A2(_02882_),
    .B1(_02883_),
    .X(_02884_));
 sky130_fd_sc_hd__a21o_1 _23015_ (.A1(_02881_),
    .A2(_02882_),
    .B1(_02884_),
    .X(_02885_));
 sky130_fd_sc_hd__and2_1 _23016_ (.A(_02880_),
    .B(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__nor2_1 _23017_ (.A(_02880_),
    .B(_02885_),
    .Y(_02887_));
 sky130_fd_sc_hd__nor2_1 _23018_ (.A(_02886_),
    .B(_02887_),
    .Y(_02888_));
 sky130_fd_sc_hd__xnor2_2 _23019_ (.A(_02875_),
    .B(_02888_),
    .Y(_02889_));
 sky130_fd_sc_hd__nand2_2 _23020_ (.A(net4949),
    .B(net4740),
    .Y(_02890_));
 sky130_fd_sc_hd__nand2_1 _23021_ (.A(net4969),
    .B(net4715),
    .Y(_02891_));
 sky130_fd_sc_hd__nand2_1 _23022_ (.A(net4982),
    .B(net4694),
    .Y(_02892_));
 sky130_fd_sc_hd__xnor2_1 _23023_ (.A(_02891_),
    .B(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__xnor2_2 _23024_ (.A(_02890_),
    .B(_02893_),
    .Y(_02894_));
 sky130_fd_sc_hd__nand2_1 _23025_ (.A(net5015),
    .B(net4693),
    .Y(_02895_));
 sky130_fd_sc_hd__nand2_1 _23026_ (.A(net5037),
    .B(net4684),
    .Y(_02896_));
 sky130_fd_sc_hd__nand2_1 _23027_ (.A(net5062),
    .B(net4647),
    .Y(_02897_));
 sky130_fd_sc_hd__o21a_1 _23028_ (.A1(_02895_),
    .A2(_02896_),
    .B1(_02897_),
    .X(_02898_));
 sky130_fd_sc_hd__a21oi_1 _23029_ (.A1(_02895_),
    .A2(_02896_),
    .B1(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__nand2_1 _23030_ (.A(net4968),
    .B(net4740),
    .Y(_02900_));
 sky130_fd_sc_hd__nand2_1 _23031_ (.A(net4948),
    .B(net4753),
    .Y(_02901_));
 sky130_fd_sc_hd__nand2_1 _23032_ (.A(_02900_),
    .B(_02901_),
    .Y(_02902_));
 sky130_fd_sc_hd__nor2_1 _23033_ (.A(_02900_),
    .B(_02901_),
    .Y(_02903_));
 sky130_fd_sc_hd__a31o_1 _23034_ (.A1(net4981),
    .A2(net4715),
    .A3(_02902_),
    .B1(_02903_),
    .X(_02904_));
 sky130_fd_sc_hd__nand2_1 _23035_ (.A(_02899_),
    .B(_02904_),
    .Y(_02905_));
 sky130_fd_sc_hd__or2_1 _23036_ (.A(_02899_),
    .B(_02904_),
    .X(_02906_));
 sky130_fd_sc_hd__nand2_1 _23037_ (.A(_02905_),
    .B(_02906_),
    .Y(_02907_));
 sky130_fd_sc_hd__xnor2_2 _23038_ (.A(_02894_),
    .B(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__nand2_1 _23039_ (.A(net5113),
    .B(net4623),
    .Y(_02909_));
 sky130_fd_sc_hd__nand2_1 _23040_ (.A(net5087),
    .B(net4647),
    .Y(_02910_));
 sky130_fd_sc_hd__nand2_1 _23041_ (.A(net5142),
    .B(net4610),
    .Y(_02911_));
 sky130_fd_sc_hd__o21ai_1 _23042_ (.A1(_02909_),
    .A2(_02910_),
    .B1(_02911_),
    .Y(_02912_));
 sky130_fd_sc_hd__a21bo_1 _23043_ (.A1(_02909_),
    .A2(_02910_),
    .B1_N(_02912_),
    .X(_02913_));
 sky130_fd_sc_hd__xnor2_1 _23044_ (.A(_02882_),
    .B(_02883_),
    .Y(_02914_));
 sky130_fd_sc_hd__xnor2_2 _23045_ (.A(_02881_),
    .B(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__xor2_1 _23046_ (.A(_02897_),
    .B(_02896_),
    .X(_02916_));
 sky130_fd_sc_hd__xnor2_1 _23047_ (.A(_02895_),
    .B(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hd__o21ba_1 _23048_ (.A1(_02913_),
    .A2(_02915_),
    .B1_N(_02917_),
    .X(_02918_));
 sky130_fd_sc_hd__a21oi_1 _23049_ (.A1(_02913_),
    .A2(_02915_),
    .B1(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__a21bo_1 _23050_ (.A1(_02889_),
    .A2(_02908_),
    .B1_N(_02919_),
    .X(_02920_));
 sky130_fd_sc_hd__o21a_1 _23051_ (.A1(_02889_),
    .A2(_02908_),
    .B1(_02920_),
    .X(_02921_));
 sky130_fd_sc_hd__xor2_1 _23052_ (.A(net4865),
    .B(net4742),
    .X(_02922_));
 sky130_fd_sc_hd__a21o_1 _23053_ (.A1(net4865),
    .A2(net4772),
    .B1(net4913),
    .X(_02923_));
 sky130_fd_sc_hd__o21ai_1 _23054_ (.A1(net4742),
    .A2(net4772),
    .B1(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__inv_2 _23055_ (.A(net4911),
    .Y(_02925_));
 sky130_fd_sc_hd__and3b_1 _23056_ (.A_N(net4772),
    .B(net4742),
    .C(net4913),
    .X(_02926_));
 sky130_fd_sc_hd__a31o_1 _23057_ (.A1(_02925_),
    .A2(net4865),
    .A3(net4772),
    .B1(_02926_),
    .X(_02927_));
 sky130_fd_sc_hd__nand2_1 _23058_ (.A(net4887),
    .B(net4760),
    .Y(_02928_));
 sky130_fd_sc_hd__mux2_1 _23059_ (.A0(_02924_),
    .A1(_02927_),
    .S(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__a31o_1 _23060_ (.A1(net4913),
    .A2(net4772),
    .A3(_02922_),
    .B1(_02929_),
    .X(_02930_));
 sky130_fd_sc_hd__a21boi_1 _23061_ (.A1(_02894_),
    .A2(_02905_),
    .B1_N(_02906_),
    .Y(_02931_));
 sky130_fd_sc_hd__xnor2_2 _23062_ (.A(net2026),
    .B(net1678),
    .Y(_02932_));
 sky130_fd_sc_hd__nand2_1 _23063_ (.A(net5092),
    .B(net4588),
    .Y(_02933_));
 sky130_fd_sc_hd__nand2_1 _23064_ (.A(net5147),
    .B(net4561),
    .Y(_02934_));
 sky130_fd_sc_hd__nand2_1 _23065_ (.A(net5118),
    .B(net4574),
    .Y(_02935_));
 sky130_fd_sc_hd__xnor2_1 _23066_ (.A(_02934_),
    .B(_02935_),
    .Y(_02936_));
 sky130_fd_sc_hd__xnor2_1 _23067_ (.A(_02933_),
    .B(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__o21ai_1 _23068_ (.A1(_02876_),
    .A2(_02878_),
    .B1(_02877_),
    .Y(_02938_));
 sky130_fd_sc_hd__a21bo_1 _23069_ (.A1(_02876_),
    .A2(_02878_),
    .B1_N(_02938_),
    .X(_02939_));
 sky130_fd_sc_hd__nand2_2 _23070_ (.A(net5017),
    .B(net4655),
    .Y(_02940_));
 sky130_fd_sc_hd__nand2_1 _23071_ (.A(net5068),
    .B(net4608),
    .Y(_02941_));
 sky130_fd_sc_hd__nand2_1 _23072_ (.A(net5041),
    .B(net4634),
    .Y(_02942_));
 sky130_fd_sc_hd__xnor2_1 _23073_ (.A(_02941_),
    .B(_02942_),
    .Y(_02943_));
 sky130_fd_sc_hd__xnor2_2 _23074_ (.A(_02940_),
    .B(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__xnor2_1 _23075_ (.A(_02939_),
    .B(_02944_),
    .Y(_02945_));
 sky130_fd_sc_hd__xnor2_2 _23076_ (.A(net2432),
    .B(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__nand2_1 _23077_ (.A(_02880_),
    .B(_02885_),
    .Y(_02947_));
 sky130_fd_sc_hd__a21oi_1 _23078_ (.A1(_02947_),
    .A2(_02875_),
    .B1(_02887_),
    .Y(_02948_));
 sky130_fd_sc_hd__nand2_1 _23079_ (.A(net4949),
    .B(net4722),
    .Y(_02949_));
 sky130_fd_sc_hd__nand2_1 _23080_ (.A(net5001),
    .B(net4685),
    .Y(_02950_));
 sky130_fd_sc_hd__nand2_1 _23081_ (.A(net4969),
    .B(net4712),
    .Y(_02951_));
 sky130_fd_sc_hd__xnor2_1 _23082_ (.A(_02950_),
    .B(_02951_),
    .Y(_02952_));
 sky130_fd_sc_hd__xnor2_2 _23083_ (.A(_02949_),
    .B(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hd__nand2_1 _23084_ (.A(_02871_),
    .B(_02873_),
    .Y(_02954_));
 sky130_fd_sc_hd__nor2_1 _23085_ (.A(_02871_),
    .B(_02873_),
    .Y(_02955_));
 sky130_fd_sc_hd__a31o_1 _23086_ (.A1(net5069),
    .A2(net4629),
    .A3(_02954_),
    .B1(_02955_),
    .X(_02956_));
 sky130_fd_sc_hd__nand2_1 _23087_ (.A(_02890_),
    .B(_02891_),
    .Y(_02957_));
 sky130_fd_sc_hd__nor2_1 _23088_ (.A(_02890_),
    .B(_02891_),
    .Y(_02958_));
 sky130_fd_sc_hd__a31o_1 _23089_ (.A1(net5001),
    .A2(net4694),
    .A3(_02957_),
    .B1(_02958_),
    .X(_02959_));
 sky130_fd_sc_hd__xnor2_1 _23090_ (.A(_02956_),
    .B(_02959_),
    .Y(_02960_));
 sky130_fd_sc_hd__xnor2_2 _23091_ (.A(_02953_),
    .B(_02960_),
    .Y(_02961_));
 sky130_fd_sc_hd__xnor2_1 _23092_ (.A(_02948_),
    .B(_02961_),
    .Y(_02962_));
 sky130_fd_sc_hd__xnor2_2 _23093_ (.A(_02946_),
    .B(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__xnor2_1 _23094_ (.A(_02932_),
    .B(_02963_),
    .Y(_02964_));
 sky130_fd_sc_hd__xnor2_2 _23095_ (.A(net1032),
    .B(_02964_),
    .Y(_02965_));
 sky130_fd_sc_hd__nand2_1 _23096_ (.A(net4904),
    .B(net4771),
    .Y(_02966_));
 sky130_fd_sc_hd__nand2_1 _23097_ (.A(net4912),
    .B(net4758),
    .Y(_02967_));
 sky130_fd_sc_hd__xor2_2 _23098_ (.A(_02966_),
    .B(_02967_),
    .X(_02968_));
 sky130_fd_sc_hd__nand2_1 _23099_ (.A(net5037),
    .B(net4693),
    .Y(_02969_));
 sky130_fd_sc_hd__nand2_1 _23100_ (.A(net5015),
    .B(net4718),
    .Y(_02970_));
 sky130_fd_sc_hd__nand2_1 _23101_ (.A(_02969_),
    .B(_02970_),
    .Y(_02971_));
 sky130_fd_sc_hd__nor2_1 _23102_ (.A(_02969_),
    .B(_02970_),
    .Y(_02972_));
 sky130_fd_sc_hd__a31o_1 _23103_ (.A1(net5062),
    .A2(net4683),
    .A3(_02971_),
    .B1(_02972_),
    .X(_02973_));
 sky130_fd_sc_hd__nand2_1 _23104_ (.A(net4968),
    .B(net4755),
    .Y(_02974_));
 sky130_fd_sc_hd__nand2_1 _23105_ (.A(net4948),
    .B(net4774),
    .Y(_02975_));
 sky130_fd_sc_hd__nand2_1 _23106_ (.A(_02974_),
    .B(_02975_),
    .Y(_02976_));
 sky130_fd_sc_hd__nor2_1 _23107_ (.A(_02974_),
    .B(_02975_),
    .Y(_02977_));
 sky130_fd_sc_hd__a31o_1 _23108_ (.A1(net4981),
    .A2(net4739),
    .A3(_02976_),
    .B1(_02977_),
    .X(_02978_));
 sky130_fd_sc_hd__nand2_1 _23109_ (.A(net5000),
    .B(net4718),
    .Y(_02979_));
 sky130_fd_sc_hd__xnor2_1 _23110_ (.A(_02900_),
    .B(_02901_),
    .Y(_02980_));
 sky130_fd_sc_hd__xnor2_2 _23111_ (.A(_02979_),
    .B(_02980_),
    .Y(_02981_));
 sky130_fd_sc_hd__o21ba_1 _23112_ (.A1(_02973_),
    .A2(_02978_),
    .B1_N(_02981_),
    .X(_02982_));
 sky130_fd_sc_hd__a21o_1 _23113_ (.A1(_02973_),
    .A2(_02978_),
    .B1(_02982_),
    .X(_02983_));
 sky130_fd_sc_hd__nor2_1 _23114_ (.A(_02968_),
    .B(net1677),
    .Y(_02984_));
 sky130_fd_sc_hd__xor2_1 _23115_ (.A(_02908_),
    .B(_02919_),
    .X(_02985_));
 sky130_fd_sc_hd__xnor2_1 _23116_ (.A(_02889_),
    .B(_02985_),
    .Y(_02986_));
 sky130_fd_sc_hd__nand2_1 _23117_ (.A(_02968_),
    .B(net1677),
    .Y(_02987_));
 sky130_fd_sc_hd__a21o_1 _23118_ (.A1(net1031),
    .A2(_02987_),
    .B1(_02984_),
    .X(_02988_));
 sky130_fd_sc_hd__xnor2_1 _23119_ (.A(_02973_),
    .B(_02978_),
    .Y(_02989_));
 sky130_fd_sc_hd__xnor2_2 _23120_ (.A(_02981_),
    .B(_02989_),
    .Y(_02990_));
 sky130_fd_sc_hd__nand2_1 _23121_ (.A(net5062),
    .B(net4683),
    .Y(_02991_));
 sky130_fd_sc_hd__xnor2_1 _23122_ (.A(_02969_),
    .B(_02970_),
    .Y(_02992_));
 sky130_fd_sc_hd__xnor2_2 _23123_ (.A(_02991_),
    .B(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__xnor2_1 _23124_ (.A(_02909_),
    .B(_02910_),
    .Y(_02994_));
 sky130_fd_sc_hd__xnor2_1 _23125_ (.A(_02911_),
    .B(_02994_),
    .Y(_02995_));
 sky130_fd_sc_hd__nand2_1 _23126_ (.A(net5130),
    .B(net4657),
    .Y(_02996_));
 sky130_fd_sc_hd__nand2_1 _23127_ (.A(net5085),
    .B(net4683),
    .Y(_02997_));
 sky130_fd_sc_hd__nand2_1 _23128_ (.A(_02996_),
    .B(_02997_),
    .Y(_02998_));
 sky130_fd_sc_hd__nor2_1 _23129_ (.A(_02996_),
    .B(_02997_),
    .Y(_02999_));
 sky130_fd_sc_hd__a31o_1 _23130_ (.A1(net5143),
    .A2(net4631),
    .A3(_02998_),
    .B1(_02999_),
    .X(_03000_));
 sky130_fd_sc_hd__o21ba_1 _23131_ (.A1(_02993_),
    .A2(net2431),
    .B1_N(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__a21o_1 _23132_ (.A1(_02993_),
    .A2(net2431),
    .B1(_03001_),
    .X(_03002_));
 sky130_fd_sc_hd__xor2_1 _23133_ (.A(_02913_),
    .B(_02915_),
    .X(_03003_));
 sky130_fd_sc_hd__xnor2_1 _23134_ (.A(_02917_),
    .B(_03003_),
    .Y(_03004_));
 sky130_fd_sc_hd__o21a_1 _23135_ (.A1(_02990_),
    .A2(_03002_),
    .B1(net1676),
    .X(_03005_));
 sky130_fd_sc_hd__a21o_1 _23136_ (.A1(_02990_),
    .A2(_03002_),
    .B1(_03005_),
    .X(_03006_));
 sky130_fd_sc_hd__nor3_1 _23137_ (.A(_03006_),
    .B(net1031),
    .C(_02987_),
    .Y(_03007_));
 sky130_fd_sc_hd__a221o_1 _23138_ (.A1(_02984_),
    .A2(net1031),
    .B1(_02988_),
    .B2(_03006_),
    .C1(_03007_),
    .X(_03008_));
 sky130_fd_sc_hd__xor2_1 _23139_ (.A(_02965_),
    .B(_03008_),
    .X(_03009_));
 sky130_fd_sc_hd__nand2_1 _23140_ (.A(net5140),
    .B(net4648),
    .Y(_03010_));
 sky130_fd_sc_hd__nand2_1 _23141_ (.A(net5084),
    .B(net4697),
    .Y(_03011_));
 sky130_fd_sc_hd__nand2_1 _23142_ (.A(net5112),
    .B(net4681),
    .Y(_03012_));
 sky130_fd_sc_hd__xnor2_1 _23143_ (.A(_03011_),
    .B(_03012_),
    .Y(_03013_));
 sky130_fd_sc_hd__xnor2_2 _23144_ (.A(_03010_),
    .B(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__nand2_2 _23145_ (.A(net5084),
    .B(net4716),
    .Y(_03015_));
 sky130_fd_sc_hd__nand2_1 _23146_ (.A(net5112),
    .B(net4697),
    .Y(_03016_));
 sky130_fd_sc_hd__nand2_1 _23147_ (.A(net5140),
    .B(net4681),
    .Y(_03017_));
 sky130_fd_sc_hd__o21ai_1 _23148_ (.A1(_03015_),
    .A2(_03016_),
    .B1(_03017_),
    .Y(_03018_));
 sky130_fd_sc_hd__a21bo_1 _23149_ (.A1(_03015_),
    .A2(_03016_),
    .B1_N(_03018_),
    .X(_03019_));
 sky130_fd_sc_hd__nand2_2 _23150_ (.A(net5012),
    .B(net4754),
    .Y(_03020_));
 sky130_fd_sc_hd__nand2_1 _23151_ (.A(net5064),
    .B(net4716),
    .Y(_03021_));
 sky130_fd_sc_hd__nand2_1 _23152_ (.A(net5039),
    .B(net4738),
    .Y(_03022_));
 sky130_fd_sc_hd__xnor2_1 _23153_ (.A(_03021_),
    .B(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__xnor2_2 _23154_ (.A(_03020_),
    .B(_03023_),
    .Y(_03024_));
 sky130_fd_sc_hd__xnor2_1 _23155_ (.A(_03019_),
    .B(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__xnor2_2 _23156_ (.A(_03014_),
    .B(_03025_),
    .Y(_03026_));
 sky130_fd_sc_hd__nand2_1 _23157_ (.A(net4983),
    .B(net4776),
    .Y(_03027_));
 sky130_fd_sc_hd__nand2_1 _23158_ (.A(net5039),
    .B(net4754),
    .Y(_03028_));
 sky130_fd_sc_hd__nand2_1 _23159_ (.A(net5013),
    .B(net4776),
    .Y(_03029_));
 sky130_fd_sc_hd__nand2_1 _23160_ (.A(net5064),
    .B(net4735),
    .Y(_03030_));
 sky130_fd_sc_hd__a21o_1 _23161_ (.A1(_03028_),
    .A2(_03029_),
    .B1(_03030_),
    .X(_03031_));
 sky130_fd_sc_hd__o21ai_2 _23162_ (.A1(_03028_),
    .A2(_03029_),
    .B1(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__xor2_2 _23163_ (.A(_03027_),
    .B(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__xnor2_1 _23164_ (.A(_03016_),
    .B(_03017_),
    .Y(_03034_));
 sky130_fd_sc_hd__xnor2_2 _23165_ (.A(_03015_),
    .B(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__xnor2_1 _23166_ (.A(_03028_),
    .B(_03029_),
    .Y(_03036_));
 sky130_fd_sc_hd__xnor2_1 _23167_ (.A(_03030_),
    .B(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__or2_1 _23168_ (.A(_03035_),
    .B(_03037_),
    .X(_03038_));
 sky130_fd_sc_hd__and2_1 _23169_ (.A(net5090),
    .B(net4736),
    .X(_03039_));
 sky130_fd_sc_hd__a21o_1 _23170_ (.A1(net5116),
    .A2(net4719),
    .B1(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__a32o_1 _23171_ (.A1(net5116),
    .A2(net4719),
    .A3(_03039_),
    .B1(net4698),
    .B2(net5139),
    .X(_03041_));
 sky130_fd_sc_hd__nand2_1 _23172_ (.A(_03040_),
    .B(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__a21o_1 _23173_ (.A1(_03035_),
    .A2(_03037_),
    .B1(_03042_),
    .X(_03043_));
 sky130_fd_sc_hd__nand3_1 _23174_ (.A(_03033_),
    .B(_03038_),
    .C(_03043_),
    .Y(_03044_));
 sky130_fd_sc_hd__a21o_1 _23175_ (.A1(_03038_),
    .A2(_03043_),
    .B1(_03033_),
    .X(_03045_));
 sky130_fd_sc_hd__and3_1 _23176_ (.A(_03026_),
    .B(_03044_),
    .C(_03045_),
    .X(_03046_));
 sky130_fd_sc_hd__a21oi_1 _23177_ (.A1(_03044_),
    .A2(_03045_),
    .B1(_03026_),
    .Y(_03047_));
 sky130_fd_sc_hd__nor2_1 _23178_ (.A(_03046_),
    .B(_03047_),
    .Y(_03048_));
 sky130_fd_sc_hd__nand2_1 _23179_ (.A(net5089),
    .B(net4757),
    .Y(_03049_));
 sky130_fd_sc_hd__nand2_1 _23180_ (.A(net5115),
    .B(net4737),
    .Y(_03050_));
 sky130_fd_sc_hd__nand2_1 _23181_ (.A(_03049_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__nor2_1 _23182_ (.A(_03049_),
    .B(_03050_),
    .Y(_03052_));
 sky130_fd_sc_hd__a31o_1 _23183_ (.A1(net5145),
    .A2(net4723),
    .A3(_03051_),
    .B1(_03052_),
    .X(_03053_));
 sky130_fd_sc_hd__nand2_1 _23184_ (.A(net5040),
    .B(net4777),
    .Y(_03054_));
 sky130_fd_sc_hd__nand2_1 _23185_ (.A(net5065),
    .B(net4757),
    .Y(_03055_));
 sky130_fd_sc_hd__xor2_2 _23186_ (.A(_03054_),
    .B(_03055_),
    .X(_03056_));
 sky130_fd_sc_hd__nand2_1 _23187_ (.A(net5139),
    .B(net4698),
    .Y(_03057_));
 sky130_fd_sc_hd__nand2_1 _23188_ (.A(net5116),
    .B(net4719),
    .Y(_03058_));
 sky130_fd_sc_hd__xor2_1 _23189_ (.A(_03058_),
    .B(_03039_),
    .X(_03059_));
 sky130_fd_sc_hd__xnor2_1 _23190_ (.A(_03057_),
    .B(_03059_),
    .Y(_03060_));
 sky130_fd_sc_hd__o21ba_1 _23191_ (.A1(_03053_),
    .A2(_03056_),
    .B1_N(_03060_),
    .X(_03061_));
 sky130_fd_sc_hd__a21oi_1 _23192_ (.A1(_03053_),
    .A2(_03056_),
    .B1(_03061_),
    .Y(_03062_));
 sky130_fd_sc_hd__xor2_1 _23193_ (.A(_03037_),
    .B(_03042_),
    .X(_03063_));
 sky130_fd_sc_hd__xnor2_1 _23194_ (.A(_03035_),
    .B(_03063_),
    .Y(_03064_));
 sky130_fd_sc_hd__and2_1 _23195_ (.A(net4757),
    .B(net4777),
    .X(_03065_));
 sky130_fd_sc_hd__and3_1 _23196_ (.A(net5065),
    .B(net5040),
    .C(_03065_),
    .X(_03066_));
 sky130_fd_sc_hd__nor2_1 _23197_ (.A(_03064_),
    .B(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hd__nand2_1 _23198_ (.A(_03064_),
    .B(_03066_),
    .Y(_03068_));
 sky130_fd_sc_hd__o21a_1 _23199_ (.A1(_03062_),
    .A2(_03067_),
    .B1(_03068_),
    .X(_03069_));
 sky130_fd_sc_hd__inv_2 _23200_ (.A(_03062_),
    .Y(_03070_));
 sky130_fd_sc_hd__or3b_1 _23201_ (.A(_03046_),
    .B(_03047_),
    .C_N(_03068_),
    .X(_03071_));
 sky130_fd_sc_hd__a2bb2o_1 _23202_ (.A1_N(_03067_),
    .A2_N(_03048_),
    .B1(_03070_),
    .B2(_03071_),
    .X(_03072_));
 sky130_fd_sc_hd__a22o_1 _23203_ (.A1(net5111),
    .A2(net4756),
    .B1(net4772),
    .B2(net5089),
    .X(_03073_));
 sky130_fd_sc_hd__and2_1 _23204_ (.A(net5111),
    .B(net5083),
    .X(_03074_));
 sky130_fd_sc_hd__a32o_1 _23205_ (.A1(net5158),
    .A2(net4742),
    .A3(_03073_),
    .B1(_03074_),
    .B2(net3752),
    .X(_03075_));
 sky130_fd_sc_hd__nand2_1 _23206_ (.A(net5157),
    .B(net4723),
    .Y(_03076_));
 sky130_fd_sc_hd__xor2_1 _23207_ (.A(_03049_),
    .B(_03050_),
    .X(_03077_));
 sky130_fd_sc_hd__xnor2_1 _23208_ (.A(_03076_),
    .B(_03077_),
    .Y(_03078_));
 sky130_fd_sc_hd__nor2_1 _23209_ (.A(net5104),
    .B(net4736),
    .Y(_03079_));
 sky130_fd_sc_hd__o2111a_1 _23210_ (.A1(_03039_),
    .A2(_03079_),
    .B1(net5157),
    .C1(net5116),
    .D1(net3752),
    .X(_03080_));
 sky130_fd_sc_hd__a21o_1 _23211_ (.A1(net5070),
    .A2(net4778),
    .B1(_03080_),
    .X(_03081_));
 sky130_fd_sc_hd__o21a_1 _23212_ (.A1(_03075_),
    .A2(_03078_),
    .B1(_03081_),
    .X(_03082_));
 sky130_fd_sc_hd__and2_1 _23213_ (.A(_03075_),
    .B(_03078_),
    .X(_03083_));
 sky130_fd_sc_hd__and2_1 _23214_ (.A(net5065),
    .B(_03080_),
    .X(_03084_));
 sky130_fd_sc_hd__or3_1 _23215_ (.A(_03082_),
    .B(_03083_),
    .C(_03084_),
    .X(_03085_));
 sky130_fd_sc_hd__xnor2_1 _23216_ (.A(_03053_),
    .B(_03056_),
    .Y(_03086_));
 sky130_fd_sc_hd__or2_1 _23217_ (.A(_03060_),
    .B(_03086_),
    .X(_03087_));
 sky130_fd_sc_hd__nand2_1 _23218_ (.A(_03060_),
    .B(_03086_),
    .Y(_03088_));
 sky130_fd_sc_hd__a32o_1 _23219_ (.A1(_03085_),
    .A2(_03087_),
    .A3(_03088_),
    .B1(_03084_),
    .B2(_03083_),
    .X(_03089_));
 sky130_fd_sc_hd__a2bb2o_1 _23220_ (.A1_N(_03048_),
    .A2_N(_03069_),
    .B1(_03072_),
    .B2(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__xor2_1 _23221_ (.A(net2431),
    .B(_03000_),
    .X(_03091_));
 sky130_fd_sc_hd__xnor2_2 _23222_ (.A(_02993_),
    .B(_03091_),
    .Y(_03092_));
 sky130_fd_sc_hd__nand2_2 _23223_ (.A(net5012),
    .B(net4738),
    .Y(_03093_));
 sky130_fd_sc_hd__nand2_1 _23224_ (.A(net5063),
    .B(net4696),
    .Y(_03094_));
 sky130_fd_sc_hd__nand2_1 _23225_ (.A(net5038),
    .B(net4717),
    .Y(_03095_));
 sky130_fd_sc_hd__xnor2_1 _23226_ (.A(_03094_),
    .B(_03095_),
    .Y(_03096_));
 sky130_fd_sc_hd__xnor2_2 _23227_ (.A(_03093_),
    .B(_03096_),
    .Y(_03097_));
 sky130_fd_sc_hd__nand2_1 _23228_ (.A(net5143),
    .B(net4631),
    .Y(_03098_));
 sky130_fd_sc_hd__xnor2_1 _23229_ (.A(_02996_),
    .B(_02997_),
    .Y(_03099_));
 sky130_fd_sc_hd__xnor2_2 _23230_ (.A(_03098_),
    .B(_03099_),
    .Y(_03100_));
 sky130_fd_sc_hd__o21ai_1 _23231_ (.A1(_03011_),
    .A2(_03012_),
    .B1(_03010_),
    .Y(_03101_));
 sky130_fd_sc_hd__a21bo_1 _23232_ (.A1(_03011_),
    .A2(_03012_),
    .B1_N(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__o21a_1 _23233_ (.A1(_03097_),
    .A2(_03100_),
    .B1(net2430),
    .X(_03103_));
 sky130_fd_sc_hd__a21o_1 _23234_ (.A1(_03097_),
    .A2(_03100_),
    .B1(_03103_),
    .X(_03104_));
 sky130_fd_sc_hd__nand2_1 _23235_ (.A(net5000),
    .B(net4739),
    .Y(_03105_));
 sky130_fd_sc_hd__xnor2_1 _23236_ (.A(_02974_),
    .B(_02975_),
    .Y(_03106_));
 sky130_fd_sc_hd__xnor2_2 _23237_ (.A(_03105_),
    .B(_03106_),
    .Y(_03107_));
 sky130_fd_sc_hd__nand3_1 _23238_ (.A(net4984),
    .B(net4967),
    .C(_03065_),
    .Y(_03108_));
 sky130_fd_sc_hd__o21a_1 _23239_ (.A1(_03093_),
    .A2(_03095_),
    .B1(_03094_),
    .X(_03109_));
 sky130_fd_sc_hd__a21o_1 _23240_ (.A1(_03093_),
    .A2(_03095_),
    .B1(_03109_),
    .X(_03110_));
 sky130_fd_sc_hd__xnor2_1 _23241_ (.A(net3060),
    .B(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__xnor2_2 _23242_ (.A(_03107_),
    .B(_03111_),
    .Y(_03112_));
 sky130_fd_sc_hd__xnor2_1 _23243_ (.A(_03104_),
    .B(_03112_),
    .Y(_03113_));
 sky130_fd_sc_hd__xnor2_2 _23244_ (.A(_03092_),
    .B(_03113_),
    .Y(_03114_));
 sky130_fd_sc_hd__o21a_1 _23245_ (.A1(_03020_),
    .A2(_03022_),
    .B1(_03021_),
    .X(_03115_));
 sky130_fd_sc_hd__a21o_1 _23246_ (.A1(_03020_),
    .A2(_03022_),
    .B1(_03115_),
    .X(_03116_));
 sky130_fd_sc_hd__nand2_1 _23247_ (.A(net4966),
    .B(net4776),
    .Y(_03117_));
 sky130_fd_sc_hd__nand2_1 _23248_ (.A(net4983),
    .B(net4754),
    .Y(_03118_));
 sky130_fd_sc_hd__xnor2_2 _23249_ (.A(_03117_),
    .B(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__or2_1 _23250_ (.A(_03116_),
    .B(_03119_),
    .X(_03120_));
 sky130_fd_sc_hd__o21ai_1 _23251_ (.A1(_03014_),
    .A2(_03024_),
    .B1(_03019_),
    .Y(_03121_));
 sky130_fd_sc_hd__nand2_1 _23252_ (.A(_03014_),
    .B(_03024_),
    .Y(_03122_));
 sky130_fd_sc_hd__xor2_2 _23253_ (.A(_03116_),
    .B(_03119_),
    .X(_03123_));
 sky130_fd_sc_hd__a21o_1 _23254_ (.A1(_03121_),
    .A2(_03122_),
    .B1(_03123_),
    .X(_03124_));
 sky130_fd_sc_hd__xor2_1 _23255_ (.A(net2430),
    .B(_03100_),
    .X(_03125_));
 sky130_fd_sc_hd__xnor2_2 _23256_ (.A(_03097_),
    .B(_03125_),
    .Y(_03126_));
 sky130_fd_sc_hd__and3_1 _23257_ (.A(_03121_),
    .B(_03122_),
    .C(_03123_),
    .X(_03127_));
 sky130_fd_sc_hd__a21oi_2 _23258_ (.A1(_03124_),
    .A2(_03126_),
    .B1(_03127_),
    .Y(_03128_));
 sky130_fd_sc_hd__xnor2_1 _23259_ (.A(_03120_),
    .B(_03128_),
    .Y(_03129_));
 sky130_fd_sc_hd__xnor2_1 _23260_ (.A(_03114_),
    .B(_03129_),
    .Y(_03130_));
 sky130_fd_sc_hd__nand2_1 _23261_ (.A(_03121_),
    .B(_03122_),
    .Y(_03131_));
 sky130_fd_sc_hd__xnor2_1 _23262_ (.A(_03131_),
    .B(_03123_),
    .Y(_03132_));
 sky130_fd_sc_hd__xnor2_1 _23263_ (.A(_03126_),
    .B(_03132_),
    .Y(_03133_));
 sky130_fd_sc_hd__and3_1 _23264_ (.A(net4983),
    .B(net4776),
    .C(_03032_),
    .X(_03134_));
 sky130_fd_sc_hd__a22oi_2 _23265_ (.A1(_03026_),
    .A2(_03033_),
    .B1(_03038_),
    .B2(_03043_),
    .Y(_03135_));
 sky130_fd_sc_hd__nand2_1 _23266_ (.A(_03134_),
    .B(_03135_),
    .Y(_03136_));
 sky130_fd_sc_hd__nor2_1 _23267_ (.A(_03026_),
    .B(_03033_),
    .Y(_03137_));
 sky130_fd_sc_hd__or3_1 _23268_ (.A(_03134_),
    .B(_03137_),
    .C(_03135_),
    .X(_03138_));
 sky130_fd_sc_hd__a21bo_1 _23269_ (.A1(_03133_),
    .A2(_03136_),
    .B1_N(_03138_),
    .X(_03139_));
 sky130_fd_sc_hd__nand2_1 _23270_ (.A(_03130_),
    .B(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hd__nor2_1 _23271_ (.A(_03137_),
    .B(_03135_),
    .Y(_03141_));
 sky130_fd_sc_hd__xnor2_1 _23272_ (.A(_03134_),
    .B(_03141_),
    .Y(_03142_));
 sky130_fd_sc_hd__xnor2_1 _23273_ (.A(_03133_),
    .B(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__nor2_1 _23274_ (.A(_03130_),
    .B(_03139_),
    .Y(_03144_));
 sky130_fd_sc_hd__a31o_1 _23275_ (.A1(_03090_),
    .A2(_03140_),
    .A3(_03143_),
    .B1(_03144_),
    .X(_03145_));
 sky130_fd_sc_hd__a21o_1 _23276_ (.A1(_03114_),
    .A2(_03128_),
    .B1(_03120_),
    .X(_03146_));
 sky130_fd_sc_hd__o21a_1 _23277_ (.A1(_03114_),
    .A2(_03128_),
    .B1(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__xor2_1 _23278_ (.A(_02990_),
    .B(_03002_),
    .X(_03148_));
 sky130_fd_sc_hd__xnor2_2 _23279_ (.A(net1676),
    .B(_03148_),
    .Y(_03149_));
 sky130_fd_sc_hd__o21a_1 _23280_ (.A1(_03104_),
    .A2(_03112_),
    .B1(_03092_),
    .X(_03150_));
 sky130_fd_sc_hd__a21o_1 _23281_ (.A1(_03104_),
    .A2(_03112_),
    .B1(_03150_),
    .X(_03151_));
 sky130_fd_sc_hd__nand2_1 _23282_ (.A(net4912),
    .B(net4775),
    .Y(_03152_));
 sky130_fd_sc_hd__o21a_1 _23283_ (.A1(_03107_),
    .A2(_03110_),
    .B1(net3060),
    .X(_03153_));
 sky130_fd_sc_hd__a21o_1 _23284_ (.A1(_03107_),
    .A2(_03110_),
    .B1(_03153_),
    .X(_03154_));
 sky130_fd_sc_hd__xor2_1 _23285_ (.A(_03152_),
    .B(_03154_),
    .X(_03155_));
 sky130_fd_sc_hd__xnor2_1 _23286_ (.A(_03151_),
    .B(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__xnor2_1 _23287_ (.A(_03149_),
    .B(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__nand2_1 _23288_ (.A(_03147_),
    .B(_03157_),
    .Y(_03158_));
 sky130_fd_sc_hd__nor2_1 _23289_ (.A(_03147_),
    .B(_03157_),
    .Y(_03159_));
 sky130_fd_sc_hd__a21o_1 _23290_ (.A1(_03145_),
    .A2(_03158_),
    .B1(_03159_),
    .X(_03160_));
 sky130_fd_sc_hd__or2b_1 _23291_ (.A(_02984_),
    .B_N(_02987_),
    .X(_03161_));
 sky130_fd_sc_hd__xnor2_1 _23292_ (.A(_03006_),
    .B(_03161_),
    .Y(_03162_));
 sky130_fd_sc_hd__nand2_1 _23293_ (.A(net1031),
    .B(_03162_),
    .Y(_03163_));
 sky130_fd_sc_hd__or2_1 _23294_ (.A(net1031),
    .B(_03162_),
    .X(_03164_));
 sky130_fd_sc_hd__and2_1 _23295_ (.A(_03163_),
    .B(_03164_),
    .X(_03165_));
 sky130_fd_sc_hd__a211o_1 _23296_ (.A1(_03145_),
    .A2(_03158_),
    .B1(_03159_),
    .C1(_03165_),
    .X(_03166_));
 sky130_fd_sc_hd__nor2_1 _23297_ (.A(_03154_),
    .B(_03151_),
    .Y(_03167_));
 sky130_fd_sc_hd__nand2_1 _23298_ (.A(_03154_),
    .B(_03151_),
    .Y(_03168_));
 sky130_fd_sc_hd__o21ai_1 _23299_ (.A1(_03149_),
    .A2(_03167_),
    .B1(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__o2bb2a_1 _23300_ (.A1_N(_03152_),
    .A2_N(_03169_),
    .B1(_03168_),
    .B2(_03149_),
    .X(_03170_));
 sky130_fd_sc_hd__a32o_1 _23301_ (.A1(_03160_),
    .A2(_03163_),
    .A3(_03164_),
    .B1(_03166_),
    .B2(_03170_),
    .X(_03171_));
 sky130_fd_sc_hd__a21o_1 _23302_ (.A1(_03160_),
    .A2(_03165_),
    .B1(_03009_),
    .X(_03172_));
 sky130_fd_sc_hd__and3b_1 _23303_ (.A_N(_03152_),
    .B(_03149_),
    .C(_03167_),
    .X(_03173_));
 sky130_fd_sc_hd__a22o_1 _23304_ (.A1(_03009_),
    .A2(_03171_),
    .B1(_03172_),
    .B2(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__inv_2 _23305_ (.A(net1031),
    .Y(_03175_));
 sky130_fd_sc_hd__nor2_1 _23306_ (.A(_02968_),
    .B(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__a21bo_1 _23307_ (.A1(_02968_),
    .A2(_03175_),
    .B1_N(_02965_),
    .X(_03177_));
 sky130_fd_sc_hd__a2bb2o_1 _23308_ (.A1_N(_02965_),
    .A2_N(_03176_),
    .B1(_03177_),
    .B2(net1677),
    .X(_03178_));
 sky130_fd_sc_hd__inv_2 _23309_ (.A(_03006_),
    .Y(_03179_));
 sky130_fd_sc_hd__a2bb2o_1 _23310_ (.A1_N(_02965_),
    .A2_N(_02988_),
    .B1(_03178_),
    .B2(_03179_),
    .X(_03180_));
 sky130_fd_sc_hd__or2_1 _23311_ (.A(net697),
    .B(net755),
    .X(_03181_));
 sky130_fd_sc_hd__a21o_1 _23312_ (.A1(_02946_),
    .A2(_02961_),
    .B1(_02948_),
    .X(_03182_));
 sky130_fd_sc_hd__o21ai_1 _23313_ (.A1(_02946_),
    .A2(_02961_),
    .B1(_03182_),
    .Y(_03183_));
 sky130_fd_sc_hd__o21ba_1 _23314_ (.A1(_02956_),
    .A2(_02959_),
    .B1_N(_02953_),
    .X(_03184_));
 sky130_fd_sc_hd__a21oi_1 _23315_ (.A1(_02956_),
    .A2(_02959_),
    .B1(_03184_),
    .Y(_03185_));
 sky130_fd_sc_hd__nand2_1 _23316_ (.A(net4864),
    .B(net4760),
    .Y(_03186_));
 sky130_fd_sc_hd__nand2_1 _23317_ (.A(net4887),
    .B(net4743),
    .Y(_03187_));
 sky130_fd_sc_hd__nand2_1 _23318_ (.A(net4723),
    .B(net4913),
    .Y(_03188_));
 sky130_fd_sc_hd__xnor2_1 _23319_ (.A(_03187_),
    .B(_03188_),
    .Y(_03189_));
 sky130_fd_sc_hd__xnor2_1 _23320_ (.A(_03186_),
    .B(_03189_),
    .Y(_03190_));
 sky130_fd_sc_hd__a22o_1 _23321_ (.A1(net4887),
    .A2(net4760),
    .B1(net4771),
    .B2(net4864),
    .X(_03191_));
 sky130_fd_sc_hd__and4_1 _23322_ (.A(net4887),
    .B(net4880),
    .C(net4760),
    .D(net4771),
    .X(_03192_));
 sky130_fd_sc_hd__a31oi_2 _23323_ (.A1(net4926),
    .A2(net4743),
    .A3(_03191_),
    .B1(_03192_),
    .Y(_03193_));
 sky130_fd_sc_hd__nand2_1 _23324_ (.A(net4850),
    .B(net4771),
    .Y(_03194_));
 sky130_fd_sc_hd__xnor2_1 _23325_ (.A(_03193_),
    .B(_03194_),
    .Y(_03195_));
 sky130_fd_sc_hd__xnor2_1 _23326_ (.A(_03190_),
    .B(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__inv_2 _23327_ (.A(net4888),
    .Y(_03197_));
 sky130_fd_sc_hd__or4b_1 _23328_ (.A(_02925_),
    .B(_03197_),
    .C(_02922_),
    .D_N(net3751),
    .X(_03198_));
 sky130_fd_sc_hd__xnor2_1 _23329_ (.A(_03196_),
    .B(net3059),
    .Y(_03199_));
 sky130_fd_sc_hd__xnor2_2 _23330_ (.A(net1675),
    .B(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__nand2_1 _23331_ (.A(net5108),
    .B(net4576),
    .Y(_03201_));
 sky130_fd_sc_hd__nand2_1 _23332_ (.A(net5124),
    .B(net4568),
    .Y(_03202_));
 sky130_fd_sc_hd__nand2_1 _23333_ (.A(net5162),
    .B(net4540),
    .Y(_03203_));
 sky130_fd_sc_hd__xnor2_1 _23334_ (.A(_03202_),
    .B(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__xnor2_1 _23335_ (.A(_03201_),
    .B(_03204_),
    .Y(_03205_));
 sky130_fd_sc_hd__o21ai_1 _23336_ (.A1(_02933_),
    .A2(_02935_),
    .B1(_02934_),
    .Y(_03206_));
 sky130_fd_sc_hd__a21bo_1 _23337_ (.A1(_02933_),
    .A2(_02935_),
    .B1_N(_03206_),
    .X(_03207_));
 sky130_fd_sc_hd__nand2_2 _23338_ (.A(net5022),
    .B(net4638),
    .Y(_03208_));
 sky130_fd_sc_hd__nand2_1 _23339_ (.A(net5057),
    .B(net4618),
    .Y(_03209_));
 sky130_fd_sc_hd__nand2_1 _23340_ (.A(net5077),
    .B(net4599),
    .Y(_03210_));
 sky130_fd_sc_hd__xnor2_1 _23341_ (.A(_03209_),
    .B(_03210_),
    .Y(_03211_));
 sky130_fd_sc_hd__xnor2_2 _23342_ (.A(_03208_),
    .B(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__xnor2_1 _23343_ (.A(_03207_),
    .B(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hd__xnor2_1 _23344_ (.A(net2429),
    .B(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__o21a_1 _23345_ (.A1(_02939_),
    .A2(_02944_),
    .B1(net2432),
    .X(_03215_));
 sky130_fd_sc_hd__a21o_1 _23346_ (.A1(_02939_),
    .A2(_02944_),
    .B1(_03215_),
    .X(_03216_));
 sky130_fd_sc_hd__nand2_2 _23347_ (.A(net4941),
    .B(net4707),
    .Y(_03217_));
 sky130_fd_sc_hd__nand2_1 _23348_ (.A(net4957),
    .B(net4673),
    .Y(_03218_));
 sky130_fd_sc_hd__nand2_1 _23349_ (.A(net4990),
    .B(net4667),
    .Y(_03219_));
 sky130_fd_sc_hd__xnor2_1 _23350_ (.A(_03218_),
    .B(_03219_),
    .Y(_03220_));
 sky130_fd_sc_hd__xnor2_2 _23351_ (.A(_03217_),
    .B(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__o21a_1 _23352_ (.A1(_02940_),
    .A2(_02942_),
    .B1(_02941_),
    .X(_03222_));
 sky130_fd_sc_hd__a21oi_2 _23353_ (.A1(_02940_),
    .A2(_02942_),
    .B1(_03222_),
    .Y(_03223_));
 sky130_fd_sc_hd__o21a_1 _23354_ (.A1(_02949_),
    .A2(_02951_),
    .B1(_02950_),
    .X(_03224_));
 sky130_fd_sc_hd__a21oi_1 _23355_ (.A1(_02949_),
    .A2(_02951_),
    .B1(_03224_),
    .Y(_03225_));
 sky130_fd_sc_hd__xnor2_1 _23356_ (.A(_03223_),
    .B(net2428),
    .Y(_03226_));
 sky130_fd_sc_hd__xnor2_2 _23357_ (.A(_03221_),
    .B(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__xnor2_1 _23358_ (.A(_03216_),
    .B(_03227_),
    .Y(_03228_));
 sky130_fd_sc_hd__xnor2_2 _23359_ (.A(net1674),
    .B(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__xnor2_1 _23360_ (.A(_03200_),
    .B(_03229_),
    .Y(_03230_));
 sky130_fd_sc_hd__xnor2_1 _23361_ (.A(_03183_),
    .B(_03230_),
    .Y(_03231_));
 sky130_fd_sc_hd__nand2_1 _23362_ (.A(net2026),
    .B(net1678),
    .Y(_03232_));
 sky130_fd_sc_hd__o21a_1 _23363_ (.A1(_02932_),
    .A2(_02963_),
    .B1(net1032),
    .X(_03233_));
 sky130_fd_sc_hd__a21o_1 _23364_ (.A1(_02932_),
    .A2(_02963_),
    .B1(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__xnor2_1 _23365_ (.A(_03232_),
    .B(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__and2_1 _23366_ (.A(_03231_),
    .B(_03235_),
    .X(_03236_));
 sky130_fd_sc_hd__nor2_1 _23367_ (.A(_03231_),
    .B(_03235_),
    .Y(_03237_));
 sky130_fd_sc_hd__a211o_1 _23368_ (.A1(net697),
    .A2(net755),
    .B1(_03236_),
    .C1(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__o21ba_1 _23369_ (.A1(_03232_),
    .A2(_03234_),
    .B1_N(_03231_),
    .X(_03239_));
 sky130_fd_sc_hd__a21o_1 _23370_ (.A1(_03232_),
    .A2(_03234_),
    .B1(_03239_),
    .X(_03240_));
 sky130_fd_sc_hd__nand2_1 _23371_ (.A(net4863),
    .B(net4741),
    .Y(_03241_));
 sky130_fd_sc_hd__nand2_1 _23372_ (.A(net4721),
    .B(net4886),
    .Y(_03242_));
 sky130_fd_sc_hd__nand2_1 _23373_ (.A(net4700),
    .B(net4914),
    .Y(_03243_));
 sky130_fd_sc_hd__xnor2_1 _23374_ (.A(_03242_),
    .B(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__xnor2_1 _23375_ (.A(_03241_),
    .B(_03244_),
    .Y(_03245_));
 sky130_fd_sc_hd__o21a_1 _23376_ (.A1(_03186_),
    .A2(_03187_),
    .B1(_03188_),
    .X(_03246_));
 sky130_fd_sc_hd__a21oi_1 _23377_ (.A1(_03186_),
    .A2(_03187_),
    .B1(_03246_),
    .Y(_03247_));
 sky130_fd_sc_hd__nand2_1 _23378_ (.A(net4833),
    .B(net4773),
    .Y(_03248_));
 sky130_fd_sc_hd__nand2_1 _23379_ (.A(net4759),
    .B(net4850),
    .Y(_03249_));
 sky130_fd_sc_hd__xor2_1 _23380_ (.A(_03248_),
    .B(_03249_),
    .X(_03250_));
 sky130_fd_sc_hd__nor2_1 _23381_ (.A(_03247_),
    .B(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__nand2_1 _23382_ (.A(_03247_),
    .B(_03250_),
    .Y(_03252_));
 sky130_fd_sc_hd__and2b_1 _23383_ (.A_N(_03251_),
    .B(_03252_),
    .X(_03253_));
 sky130_fd_sc_hd__xnor2_1 _23384_ (.A(_03245_),
    .B(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__a21o_1 _23385_ (.A1(_03193_),
    .A2(_03190_),
    .B1(_03194_),
    .X(_03255_));
 sky130_fd_sc_hd__o21a_1 _23386_ (.A1(_03193_),
    .A2(_03190_),
    .B1(_03255_),
    .X(_03256_));
 sky130_fd_sc_hd__a21bo_1 _23387_ (.A1(_03223_),
    .A2(net2428),
    .B1_N(_03221_),
    .X(_03257_));
 sky130_fd_sc_hd__o21ai_1 _23388_ (.A1(_03223_),
    .A2(net2428),
    .B1(_03257_),
    .Y(_03258_));
 sky130_fd_sc_hd__nor2_1 _23389_ (.A(_03256_),
    .B(_03258_),
    .Y(_03259_));
 sky130_fd_sc_hd__nand2_1 _23390_ (.A(_03256_),
    .B(_03258_),
    .Y(_03260_));
 sky130_fd_sc_hd__or2b_1 _23391_ (.A(_03259_),
    .B_N(_03260_),
    .X(_03261_));
 sky130_fd_sc_hd__xnor2_1 _23392_ (.A(_03254_),
    .B(_03261_),
    .Y(_03262_));
 sky130_fd_sc_hd__o21a_1 _23393_ (.A1(_03216_),
    .A2(_03227_),
    .B1(net1674),
    .X(_03263_));
 sky130_fd_sc_hd__a21o_1 _23394_ (.A1(_03216_),
    .A2(_03227_),
    .B1(_03263_),
    .X(_03264_));
 sky130_fd_sc_hd__nand2_2 _23395_ (.A(net5099),
    .B(net4563),
    .Y(_03265_));
 sky130_fd_sc_hd__nand2_1 _23396_ (.A(net5124),
    .B(net4550),
    .Y(_03266_));
 sky130_fd_sc_hd__nand2_1 _23397_ (.A(net5150),
    .B(net4525),
    .Y(_03267_));
 sky130_fd_sc_hd__xor2_1 _23398_ (.A(_03266_),
    .B(_03267_),
    .X(_03268_));
 sky130_fd_sc_hd__xnor2_2 _23399_ (.A(_03265_),
    .B(_03268_),
    .Y(_03269_));
 sky130_fd_sc_hd__o21ai_1 _23400_ (.A1(_03201_),
    .A2(_03202_),
    .B1(_03203_),
    .Y(_03270_));
 sky130_fd_sc_hd__a21bo_1 _23401_ (.A1(_03201_),
    .A2(_03202_),
    .B1_N(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__nand2_1 _23402_ (.A(net5033),
    .B(net4614),
    .Y(_03272_));
 sky130_fd_sc_hd__nand2_1 _23403_ (.A(net5054),
    .B(net4597),
    .Y(_03273_));
 sky130_fd_sc_hd__nand2_1 _23404_ (.A(net4575),
    .B(net5080),
    .Y(_03274_));
 sky130_fd_sc_hd__xnor2_1 _23405_ (.A(_03273_),
    .B(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__xnor2_1 _23406_ (.A(_03272_),
    .B(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__nor2_1 _23407_ (.A(net2427),
    .B(_03276_),
    .Y(_03277_));
 sky130_fd_sc_hd__nand2_1 _23408_ (.A(net2427),
    .B(_03276_),
    .Y(_03278_));
 sky130_fd_sc_hd__or2b_1 _23409_ (.A(_03277_),
    .B_N(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__xor2_1 _23410_ (.A(_03269_),
    .B(_03279_),
    .X(_03280_));
 sky130_fd_sc_hd__o21a_1 _23411_ (.A1(_03207_),
    .A2(_03212_),
    .B1(net2429),
    .X(_03281_));
 sky130_fd_sc_hd__a21o_1 _23412_ (.A1(_03207_),
    .A2(_03212_),
    .B1(_03281_),
    .X(_03282_));
 sky130_fd_sc_hd__nand2_2 _23413_ (.A(net4934),
    .B(net4679),
    .Y(_03283_));
 sky130_fd_sc_hd__nand2_1 _23414_ (.A(net4963),
    .B(net4666),
    .Y(_03284_));
 sky130_fd_sc_hd__nand2_1 _23415_ (.A(net4637),
    .B(net4989),
    .Y(_03285_));
 sky130_fd_sc_hd__xnor2_1 _23416_ (.A(_03284_),
    .B(_03285_),
    .Y(_03286_));
 sky130_fd_sc_hd__xnor2_2 _23417_ (.A(_03283_),
    .B(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__o21a_1 _23418_ (.A1(_03217_),
    .A2(_03218_),
    .B1(_03219_),
    .X(_03288_));
 sky130_fd_sc_hd__a21oi_2 _23419_ (.A1(_03217_),
    .A2(_03218_),
    .B1(_03288_),
    .Y(_03289_));
 sky130_fd_sc_hd__o21a_1 _23420_ (.A1(_03208_),
    .A2(_03209_),
    .B1(_03210_),
    .X(_03290_));
 sky130_fd_sc_hd__a21oi_2 _23421_ (.A1(_03208_),
    .A2(_03209_),
    .B1(_03290_),
    .Y(_03291_));
 sky130_fd_sc_hd__xnor2_1 _23422_ (.A(_03289_),
    .B(_03291_),
    .Y(_03292_));
 sky130_fd_sc_hd__xnor2_2 _23423_ (.A(_03287_),
    .B(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__xnor2_1 _23424_ (.A(_03282_),
    .B(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__xnor2_1 _23425_ (.A(net1385),
    .B(_03294_),
    .Y(_03295_));
 sky130_fd_sc_hd__and2_1 _23426_ (.A(_03264_),
    .B(net1167),
    .X(_03296_));
 sky130_fd_sc_hd__nor2_1 _23427_ (.A(_03264_),
    .B(net1167),
    .Y(_03297_));
 sky130_fd_sc_hd__nor2_1 _23428_ (.A(_03296_),
    .B(_03297_),
    .Y(_03298_));
 sky130_fd_sc_hd__xnor2_1 _23429_ (.A(_03262_),
    .B(_03298_),
    .Y(_03299_));
 sky130_fd_sc_hd__o21a_1 _23430_ (.A1(net1675),
    .A2(net3059),
    .B1(_03196_),
    .X(_03300_));
 sky130_fd_sc_hd__a21o_1 _23431_ (.A1(net1675),
    .A2(net3059),
    .B1(_03300_),
    .X(_03301_));
 sky130_fd_sc_hd__a21bo_1 _23432_ (.A1(_03200_),
    .A2(_03229_),
    .B1_N(_03183_),
    .X(_03302_));
 sky130_fd_sc_hd__o21a_1 _23433_ (.A1(_03200_),
    .A2(_03229_),
    .B1(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__xnor2_1 _23434_ (.A(net1166),
    .B(net938),
    .Y(_03304_));
 sky130_fd_sc_hd__xnor2_1 _23435_ (.A(_03299_),
    .B(_03304_),
    .Y(_03305_));
 sky130_fd_sc_hd__xnor2_1 _23436_ (.A(net749),
    .B(net796),
    .Y(_03306_));
 sky130_fd_sc_hd__inv_2 _23437_ (.A(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__a21oi_1 _23438_ (.A1(net646),
    .A2(net640),
    .B1(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hd__and3_1 _23439_ (.A(_03307_),
    .B(net646),
    .C(net640),
    .X(_03309_));
 sky130_fd_sc_hd__nor2_1 _23440_ (.A(_03308_),
    .B(_03309_),
    .Y(_03310_));
 sky130_fd_sc_hd__xor2_1 _23441_ (.A(\pid_q.curr_int[0] ),
    .B(\pid_q.prev_int[0] ),
    .X(_03311_));
 sky130_fd_sc_hd__xnor2_1 _23442_ (.A(\pid_q.prev_error[0] ),
    .B(\pid_q.curr_error[0] ),
    .Y(_03312_));
 sky130_fd_sc_hd__nor2_1 _23443_ (.A(net3999),
    .B(_03312_),
    .Y(_03313_));
 sky130_fd_sc_hd__a221o_1 _23444_ (.A1(net7466),
    .A2(net545),
    .B1(_03311_),
    .B2(net7526),
    .C1(net3056),
    .X(_03314_));
 sky130_fd_sc_hd__a22o_1 _23445_ (.A1(\pid_q.curr_int[0] ),
    .A2(net3061),
    .B1(net2028),
    .B2(_03314_),
    .X(_00665_));
 sky130_fd_sc_hd__nand2_1 _23446_ (.A(\pid_q.curr_int[0] ),
    .B(\pid_q.prev_int[0] ),
    .Y(_03315_));
 sky130_fd_sc_hd__xor2_1 _23447_ (.A(\pid_q.curr_int[1] ),
    .B(\pid_q.prev_int[1] ),
    .X(_03316_));
 sky130_fd_sc_hd__xnor2_1 _23448_ (.A(_03315_),
    .B(_03316_),
    .Y(_03317_));
 sky130_fd_sc_hd__or2_1 _23449_ (.A(net749),
    .B(net796),
    .X(_03318_));
 sky130_fd_sc_hd__o21bai_1 _23450_ (.A1(_03262_),
    .A2(_03297_),
    .B1_N(_03296_),
    .Y(_03319_));
 sky130_fd_sc_hd__o21a_1 _23451_ (.A1(_03282_),
    .A2(_03293_),
    .B1(net1385),
    .X(_03320_));
 sky130_fd_sc_hd__a21o_1 _23452_ (.A1(_03282_),
    .A2(_03293_),
    .B1(_03320_),
    .X(_03321_));
 sky130_fd_sc_hd__nand2_2 _23453_ (.A(net4597),
    .B(net5024),
    .Y(_03322_));
 sky130_fd_sc_hd__nand2_1 _23454_ (.A(net4575),
    .B(net5054),
    .Y(_03323_));
 sky130_fd_sc_hd__nand2_1 _23455_ (.A(net4563),
    .B(net5080),
    .Y(_03324_));
 sky130_fd_sc_hd__xnor2_1 _23456_ (.A(_03323_),
    .B(_03324_),
    .Y(_03325_));
 sky130_fd_sc_hd__xnor2_2 _23457_ (.A(_03322_),
    .B(_03325_),
    .Y(_03326_));
 sky130_fd_sc_hd__o21ai_1 _23458_ (.A1(_03265_),
    .A2(_03266_),
    .B1(_03267_),
    .Y(_03327_));
 sky130_fd_sc_hd__a21bo_1 _23459_ (.A1(_03265_),
    .A2(_03266_),
    .B1_N(_03327_),
    .X(_03328_));
 sky130_fd_sc_hd__nand2_1 _23460_ (.A(net5162),
    .B(net4513),
    .Y(_03329_));
 sky130_fd_sc_hd__nand2_1 _23461_ (.A(net4550),
    .B(net5099),
    .Y(_03330_));
 sky130_fd_sc_hd__nand2_1 _23462_ (.A(net4532),
    .B(net5128),
    .Y(_03331_));
 sky130_fd_sc_hd__xnor2_1 _23463_ (.A(_03330_),
    .B(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__xnor2_1 _23464_ (.A(_03329_),
    .B(_03332_),
    .Y(_03333_));
 sky130_fd_sc_hd__xnor2_1 _23465_ (.A(_03328_),
    .B(net2426),
    .Y(_03334_));
 sky130_fd_sc_hd__xnor2_2 _23466_ (.A(_03326_),
    .B(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__a21oi_2 _23467_ (.A1(_03269_),
    .A2(_03278_),
    .B1(_03277_),
    .Y(_03336_));
 sky130_fd_sc_hd__nand2_2 _23468_ (.A(net4662),
    .B(net4944),
    .Y(_03337_));
 sky130_fd_sc_hd__nand2_1 _23469_ (.A(net4641),
    .B(net4962),
    .Y(_03338_));
 sky130_fd_sc_hd__nand2_1 _23470_ (.A(net4619),
    .B(net4996),
    .Y(_03339_));
 sky130_fd_sc_hd__xnor2_1 _23471_ (.A(_03338_),
    .B(_03339_),
    .Y(_03340_));
 sky130_fd_sc_hd__xnor2_2 _23472_ (.A(_03337_),
    .B(_03340_),
    .Y(_03341_));
 sky130_fd_sc_hd__o21a_1 _23473_ (.A1(_03283_),
    .A2(_03284_),
    .B1(_03285_),
    .X(_03342_));
 sky130_fd_sc_hd__a21oi_1 _23474_ (.A1(_03283_),
    .A2(_03284_),
    .B1(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__o21a_1 _23475_ (.A1(_03272_),
    .A2(_03273_),
    .B1(_03274_),
    .X(_03344_));
 sky130_fd_sc_hd__a21oi_2 _23476_ (.A1(_03272_),
    .A2(_03273_),
    .B1(_03344_),
    .Y(_03345_));
 sky130_fd_sc_hd__xnor2_1 _23477_ (.A(net2424),
    .B(_03345_),
    .Y(_03346_));
 sky130_fd_sc_hd__xnor2_2 _23478_ (.A(_03341_),
    .B(_03346_),
    .Y(_03347_));
 sky130_fd_sc_hd__xnor2_1 _23479_ (.A(_03336_),
    .B(_03347_),
    .Y(_03348_));
 sky130_fd_sc_hd__xnor2_2 _23480_ (.A(_03335_),
    .B(_03348_),
    .Y(_03349_));
 sky130_fd_sc_hd__nand2_2 _23481_ (.A(net4727),
    .B(net4876),
    .Y(_03350_));
 sky130_fd_sc_hd__nand2_1 _23482_ (.A(net4677),
    .B(net4920),
    .Y(_03351_));
 sky130_fd_sc_hd__nand2_1 _23483_ (.A(net4702),
    .B(net4900),
    .Y(_03352_));
 sky130_fd_sc_hd__xnor2_1 _23484_ (.A(_03351_),
    .B(_03352_),
    .Y(_03353_));
 sky130_fd_sc_hd__xnor2_2 _23485_ (.A(_03350_),
    .B(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__o21ai_1 _23486_ (.A1(_03241_),
    .A2(_03242_),
    .B1(_03243_),
    .Y(_03355_));
 sky130_fd_sc_hd__a21bo_1 _23487_ (.A1(_03241_),
    .A2(_03242_),
    .B1_N(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__nand2_2 _23488_ (.A(net4784),
    .B(net4813),
    .Y(_03357_));
 sky130_fd_sc_hd__nand2_1 _23489_ (.A(net4768),
    .B(net4826),
    .Y(_03358_));
 sky130_fd_sc_hd__nand2_1 _23490_ (.A(net4749),
    .B(net4845),
    .Y(_03359_));
 sky130_fd_sc_hd__xnor2_1 _23491_ (.A(_03358_),
    .B(_03359_),
    .Y(_03360_));
 sky130_fd_sc_hd__xnor2_2 _23492_ (.A(_03357_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__xnor2_1 _23493_ (.A(net2420),
    .B(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__xnor2_2 _23494_ (.A(_03354_),
    .B(_03362_),
    .Y(_03363_));
 sky130_fd_sc_hd__a21oi_1 _23495_ (.A1(_03245_),
    .A2(_03252_),
    .B1(_03251_),
    .Y(_03364_));
 sky130_fd_sc_hd__a21bo_1 _23496_ (.A1(_03289_),
    .A2(_03291_),
    .B1_N(_03287_),
    .X(_03365_));
 sky130_fd_sc_hd__o21a_1 _23497_ (.A1(_03289_),
    .A2(_03291_),
    .B1(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__xnor2_1 _23498_ (.A(net1670),
    .B(net1667),
    .Y(_03367_));
 sky130_fd_sc_hd__xnor2_2 _23499_ (.A(_03363_),
    .B(_03367_),
    .Y(_03368_));
 sky130_fd_sc_hd__xor2_1 _23500_ (.A(_03349_),
    .B(_03368_),
    .X(_03369_));
 sky130_fd_sc_hd__xnor2_1 _23501_ (.A(net1028),
    .B(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__o21ai_1 _23502_ (.A1(_03254_),
    .A2(_03259_),
    .B1(_03260_),
    .Y(_03371_));
 sky130_fd_sc_hd__and2_1 _23503_ (.A(net4842),
    .B(net4827),
    .X(_03372_));
 sky130_fd_sc_hd__buf_1 _23504_ (.A(_03372_),
    .X(_03373_));
 sky130_fd_sc_hd__nand2_1 _23505_ (.A(net3750),
    .B(net3050),
    .Y(_03374_));
 sky130_fd_sc_hd__xor2_1 _23506_ (.A(_03371_),
    .B(_03374_),
    .X(_03375_));
 sky130_fd_sc_hd__nand2_1 _23507_ (.A(_03370_),
    .B(net1024),
    .Y(_03376_));
 sky130_fd_sc_hd__or2_1 _23508_ (.A(_03370_),
    .B(net1024),
    .X(_03377_));
 sky130_fd_sc_hd__nand2_1 _23509_ (.A(_03376_),
    .B(_03377_),
    .Y(_03378_));
 sky130_fd_sc_hd__xnor2_2 _23510_ (.A(net934),
    .B(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__o21a_1 _23511_ (.A1(net1166),
    .A2(net938),
    .B1(_03299_),
    .X(_03380_));
 sky130_fd_sc_hd__a21o_1 _23512_ (.A1(net1166),
    .A2(net938),
    .B1(_03380_),
    .X(_03381_));
 sky130_fd_sc_hd__xnor2_1 _23513_ (.A(_03379_),
    .B(net745),
    .Y(_03382_));
 sky130_fd_sc_hd__xnor2_1 _23514_ (.A(_03318_),
    .B(_03382_),
    .Y(_03383_));
 sky130_fd_sc_hd__xnor2_1 _23515_ (.A(_03309_),
    .B(_03383_),
    .Y(_03384_));
 sky130_fd_sc_hd__xnor2_1 _23516_ (.A(\pid_q.prev_error[1] ),
    .B(net5168),
    .Y(_03385_));
 sky130_fd_sc_hd__and3_1 _23517_ (.A(\pid_q.prev_error[0] ),
    .B(\pid_q.curr_error[0] ),
    .C(_03385_),
    .X(_03386_));
 sky130_fd_sc_hd__a21oi_1 _23518_ (.A1(\pid_q.prev_error[0] ),
    .A2(\pid_q.curr_error[0] ),
    .B1(_03385_),
    .Y(_03387_));
 sky130_fd_sc_hd__o21a_1 _23519_ (.A1(_03386_),
    .A2(_03387_),
    .B1(net7511),
    .X(_03388_));
 sky130_fd_sc_hd__a221o_1 _23520_ (.A1(net7526),
    .A2(_03317_),
    .B1(net540),
    .B2(net7466),
    .C1(net2417),
    .X(_03389_));
 sky130_fd_sc_hd__a22o_1 _23521_ (.A1(\pid_q.curr_int[1] ),
    .A2(net3061),
    .B1(net2028),
    .B2(_03389_),
    .X(_00666_));
 sky130_fd_sc_hd__a22o_1 _23522_ (.A1(\pid_q.curr_int[0] ),
    .A2(\pid_q.prev_int[0] ),
    .B1(\pid_q.prev_int[1] ),
    .B2(\pid_q.curr_int[1] ),
    .X(_03390_));
 sky130_fd_sc_hd__o21a_1 _23523_ (.A1(\pid_q.curr_int[1] ),
    .A2(\pid_q.prev_int[1] ),
    .B1(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__xnor2_1 _23524_ (.A(net5180),
    .B(\pid_q.prev_int[2] ),
    .Y(_03392_));
 sky130_fd_sc_hd__xnor2_1 _23525_ (.A(_03391_),
    .B(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__nand2_1 _23526_ (.A(net5163),
    .B(net4496),
    .Y(_03394_));
 sky130_fd_sc_hd__nand2_1 _23527_ (.A(net5129),
    .B(net4512),
    .Y(_03395_));
 sky130_fd_sc_hd__xnor2_1 _23528_ (.A(_03394_),
    .B(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__xnor2_1 _23529_ (.A(net4795),
    .B(_03396_),
    .Y(_03397_));
 sky130_fd_sc_hd__o21ai_1 _23530_ (.A1(_03330_),
    .A2(_03331_),
    .B1(_03329_),
    .Y(_03398_));
 sky130_fd_sc_hd__a21bo_1 _23531_ (.A1(_03330_),
    .A2(_03331_),
    .B1_N(_03398_),
    .X(_03399_));
 sky130_fd_sc_hd__nand2_1 _23532_ (.A(net4557),
    .B(net5053),
    .Y(_03400_));
 sky130_fd_sc_hd__nand2_1 _23533_ (.A(net4540),
    .B(net5079),
    .Y(_03401_));
 sky130_fd_sc_hd__nand2_1 _23534_ (.A(net4532),
    .B(net5108),
    .Y(_03402_));
 sky130_fd_sc_hd__xnor2_1 _23535_ (.A(_03401_),
    .B(_03402_),
    .Y(_03403_));
 sky130_fd_sc_hd__xnor2_1 _23536_ (.A(_03400_),
    .B(_03403_),
    .Y(_03404_));
 sky130_fd_sc_hd__nor2_1 _23537_ (.A(_03399_),
    .B(_03404_),
    .Y(_03405_));
 sky130_fd_sc_hd__nand2_1 _23538_ (.A(_03399_),
    .B(_03404_),
    .Y(_03406_));
 sky130_fd_sc_hd__or2b_1 _23539_ (.A(_03405_),
    .B_N(_03406_),
    .X(_03407_));
 sky130_fd_sc_hd__xnor2_1 _23540_ (.A(_03397_),
    .B(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__o21a_1 _23541_ (.A1(_03328_),
    .A2(net2426),
    .B1(_03326_),
    .X(_03409_));
 sky130_fd_sc_hd__a21o_1 _23542_ (.A1(_03328_),
    .A2(net2426),
    .B1(_03409_),
    .X(_03410_));
 sky130_fd_sc_hd__nand2_2 _23543_ (.A(net4619),
    .B(net4962),
    .Y(_03411_));
 sky130_fd_sc_hd__nand2_1 _23544_ (.A(net4597),
    .B(net4996),
    .Y(_03412_));
 sky130_fd_sc_hd__nand2_1 _23545_ (.A(net4575),
    .B(net5024),
    .Y(_03413_));
 sky130_fd_sc_hd__xnor2_1 _23546_ (.A(_03412_),
    .B(_03413_),
    .Y(_03414_));
 sky130_fd_sc_hd__xnor2_2 _23547_ (.A(_03411_),
    .B(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__o21a_1 _23548_ (.A1(_03337_),
    .A2(_03338_),
    .B1(_03339_),
    .X(_03416_));
 sky130_fd_sc_hd__a21oi_2 _23549_ (.A1(_03337_),
    .A2(_03338_),
    .B1(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__o21a_1 _23550_ (.A1(_03322_),
    .A2(_03323_),
    .B1(_03324_),
    .X(_03418_));
 sky130_fd_sc_hd__a21oi_2 _23551_ (.A1(_03322_),
    .A2(_03323_),
    .B1(_03418_),
    .Y(_03419_));
 sky130_fd_sc_hd__xnor2_1 _23552_ (.A(_03417_),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__xnor2_2 _23553_ (.A(_03415_),
    .B(_03420_),
    .Y(_03421_));
 sky130_fd_sc_hd__xnor2_1 _23554_ (.A(_03410_),
    .B(_03421_),
    .Y(_03422_));
 sky130_fd_sc_hd__xnor2_2 _23555_ (.A(net1384),
    .B(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__a21o_1 _23556_ (.A1(_03336_),
    .A2(_03347_),
    .B1(_03335_),
    .X(_03424_));
 sky130_fd_sc_hd__o21a_1 _23557_ (.A1(_03336_),
    .A2(_03347_),
    .B1(_03424_),
    .X(_03425_));
 sky130_fd_sc_hd__nand2_1 _23558_ (.A(net4677),
    .B(net4900),
    .Y(_03426_));
 sky130_fd_sc_hd__nand2_1 _23559_ (.A(net4664),
    .B(net4920),
    .Y(_03427_));
 sky130_fd_sc_hd__nand2_1 _23560_ (.A(net4641),
    .B(net4944),
    .Y(_03428_));
 sky130_fd_sc_hd__xnor2_1 _23561_ (.A(_03427_),
    .B(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__xnor2_1 _23562_ (.A(_03426_),
    .B(_03429_),
    .Y(_03430_));
 sky130_fd_sc_hd__o21ai_1 _23563_ (.A1(_03350_),
    .A2(_03352_),
    .B1(_03351_),
    .Y(_03431_));
 sky130_fd_sc_hd__a21bo_1 _23564_ (.A1(_03350_),
    .A2(_03352_),
    .B1_N(_03431_),
    .X(_03432_));
 sky130_fd_sc_hd__nand2_2 _23565_ (.A(net4749),
    .B(net4826),
    .Y(_03433_));
 sky130_fd_sc_hd__nand2_1 _23566_ (.A(net4727),
    .B(net4845),
    .Y(_03434_));
 sky130_fd_sc_hd__nand2_1 _23567_ (.A(net4702),
    .B(net4876),
    .Y(_03435_));
 sky130_fd_sc_hd__xnor2_1 _23568_ (.A(_03434_),
    .B(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__xnor2_2 _23569_ (.A(_03433_),
    .B(_03436_),
    .Y(_03437_));
 sky130_fd_sc_hd__xnor2_1 _23570_ (.A(_03432_),
    .B(_03437_),
    .Y(_03438_));
 sky130_fd_sc_hd__xnor2_1 _23571_ (.A(_03430_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__o21a_1 _23572_ (.A1(net2420),
    .A2(_03361_),
    .B1(_03354_),
    .X(_03440_));
 sky130_fd_sc_hd__a21o_1 _23573_ (.A1(net2420),
    .A2(_03361_),
    .B1(_03440_),
    .X(_03441_));
 sky130_fd_sc_hd__a21bo_1 _23574_ (.A1(net2424),
    .A2(_03345_),
    .B1_N(_03341_),
    .X(_03442_));
 sky130_fd_sc_hd__o21ai_2 _23575_ (.A1(net2424),
    .A2(_03345_),
    .B1(_03442_),
    .Y(_03443_));
 sky130_fd_sc_hd__xnor2_1 _23576_ (.A(_03441_),
    .B(_03443_),
    .Y(_03444_));
 sky130_fd_sc_hd__xnor2_1 _23577_ (.A(_03439_),
    .B(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__nor2_1 _23578_ (.A(_03425_),
    .B(_03445_),
    .Y(_03446_));
 sky130_fd_sc_hd__nand2_1 _23579_ (.A(_03425_),
    .B(_03445_),
    .Y(_03447_));
 sky130_fd_sc_hd__and2b_1 _23580_ (.A_N(_03446_),
    .B(_03447_),
    .X(_03448_));
 sky130_fd_sc_hd__xnor2_2 _23581_ (.A(_03423_),
    .B(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__o21a_1 _23582_ (.A1(_03349_),
    .A2(_03368_),
    .B1(net1028),
    .X(_03450_));
 sky130_fd_sc_hd__a21o_1 _23583_ (.A1(_03349_),
    .A2(_03368_),
    .B1(_03450_),
    .X(_03451_));
 sky130_fd_sc_hd__a21bo_1 _23584_ (.A1(net1670),
    .A2(net1667),
    .B1_N(_03363_),
    .X(_03452_));
 sky130_fd_sc_hd__o21ai_2 _23585_ (.A1(net1670),
    .A2(net1667),
    .B1(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__o21a_1 _23586_ (.A1(_03357_),
    .A2(_03358_),
    .B1(_03359_),
    .X(_03454_));
 sky130_fd_sc_hd__a21o_1 _23587_ (.A1(_03357_),
    .A2(_03358_),
    .B1(_03454_),
    .X(_03455_));
 sky130_fd_sc_hd__inv_2 _23588_ (.A(net4795),
    .Y(_03456_));
 sky130_fd_sc_hd__or2_1 _23589_ (.A(net4784),
    .B(net3746),
    .X(_03457_));
 sky130_fd_sc_hd__nand2_1 _23590_ (.A(net4768),
    .B(net4813),
    .Y(_03458_));
 sky130_fd_sc_hd__xnor2_1 _23591_ (.A(_03457_),
    .B(_03458_),
    .Y(_03459_));
 sky130_fd_sc_hd__xnor2_2 _23592_ (.A(_03455_),
    .B(_03459_),
    .Y(_03460_));
 sky130_fd_sc_hd__xnor2_2 _23593_ (.A(_03453_),
    .B(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__xor2_1 _23594_ (.A(_03451_),
    .B(_03461_),
    .X(_03462_));
 sky130_fd_sc_hd__xnor2_2 _23595_ (.A(_03449_),
    .B(_03462_),
    .Y(_03463_));
 sky130_fd_sc_hd__nor2_1 _23596_ (.A(_03370_),
    .B(net1024),
    .Y(_03464_));
 sky130_fd_sc_hd__o21ai_2 _23597_ (.A1(net934),
    .A2(_03464_),
    .B1(_03376_),
    .Y(_03465_));
 sky130_fd_sc_hd__nor2_1 _23598_ (.A(_03371_),
    .B(_03374_),
    .Y(_03466_));
 sky130_fd_sc_hd__xnor2_1 _23599_ (.A(_03465_),
    .B(net1020),
    .Y(_03467_));
 sky130_fd_sc_hd__xnor2_1 _23600_ (.A(_03463_),
    .B(_03467_),
    .Y(_03468_));
 sky130_fd_sc_hd__nand2_1 _23601_ (.A(_03379_),
    .B(net745),
    .Y(_03469_));
 sky130_fd_sc_hd__or2b_1 _23602_ (.A(_03469_),
    .B_N(_03318_),
    .X(_03470_));
 sky130_fd_sc_hd__o21ai_1 _23603_ (.A1(_03379_),
    .A2(net745),
    .B1(_03318_),
    .Y(_03471_));
 sky130_fd_sc_hd__a32o_1 _23604_ (.A1(_03307_),
    .A2(net646),
    .A3(net640),
    .B1(_03469_),
    .B2(_03471_),
    .X(_03472_));
 sky130_fd_sc_hd__and2_1 _23605_ (.A(_03470_),
    .B(_03472_),
    .X(_03473_));
 sky130_fd_sc_hd__xor2_1 _23606_ (.A(net696),
    .B(_03473_),
    .X(_03474_));
 sky130_fd_sc_hd__nand2_1 _23607_ (.A(\pid_q.prev_error[1] ),
    .B(net5168),
    .Y(_03475_));
 sky130_fd_sc_hd__o211ai_4 _23608_ (.A1(\pid_q.prev_error[1] ),
    .A2(net5168),
    .B1(\pid_q.prev_error[0] ),
    .C1(\pid_q.curr_error[0] ),
    .Y(_03476_));
 sky130_fd_sc_hd__xor2_1 _23609_ (.A(\pid_q.prev_error[2] ),
    .B(\pid_q.curr_error[2] ),
    .X(_03477_));
 sky130_fd_sc_hd__and3_1 _23610_ (.A(_03475_),
    .B(_03476_),
    .C(_03477_),
    .X(_03478_));
 sky130_fd_sc_hd__a21oi_1 _23611_ (.A1(_03475_),
    .A2(_03476_),
    .B1(_03477_),
    .Y(_03479_));
 sky130_fd_sc_hd__o21a_1 _23612_ (.A1(_03478_),
    .A2(_03479_),
    .B1(net7510),
    .X(_03480_));
 sky130_fd_sc_hd__a221o_1 _23613_ (.A1(net7527),
    .A2(_03393_),
    .B1(net514),
    .B2(net7468),
    .C1(net2414),
    .X(_03481_));
 sky130_fd_sc_hd__a22o_1 _23614_ (.A1(net8996),
    .A2(net3062),
    .B1(net2028),
    .B2(_03481_),
    .X(_00667_));
 sky130_fd_sc_hd__a21o_1 _23615_ (.A1(\pid_q.prev_int[2] ),
    .A2(_03391_),
    .B1(net5180),
    .X(_03482_));
 sky130_fd_sc_hd__o21ai_2 _23616_ (.A1(\pid_q.prev_int[2] ),
    .A2(_03391_),
    .B1(_03482_),
    .Y(_03483_));
 sky130_fd_sc_hd__xor2_1 _23617_ (.A(\pid_q.curr_int[3] ),
    .B(\pid_q.prev_int[3] ),
    .X(_03484_));
 sky130_fd_sc_hd__xnor2_1 _23618_ (.A(_03483_),
    .B(_03484_),
    .Y(_03485_));
 sky130_fd_sc_hd__nand2_1 _23619_ (.A(net696),
    .B(_03473_),
    .Y(_03486_));
 sky130_fd_sc_hd__o21a_1 _23620_ (.A1(_03465_),
    .A2(_03463_),
    .B1(net1020),
    .X(_03487_));
 sky130_fd_sc_hd__a21oi_1 _23621_ (.A1(_03465_),
    .A2(_03463_),
    .B1(_03487_),
    .Y(_03488_));
 sky130_fd_sc_hd__nand2_2 _23622_ (.A(net4677),
    .B(net4875),
    .Y(_03489_));
 sky130_fd_sc_hd__nand2_1 _23623_ (.A(net4636),
    .B(net4922),
    .Y(_03490_));
 sky130_fd_sc_hd__nand2_1 _23624_ (.A(net4664),
    .B(net4899),
    .Y(_03491_));
 sky130_fd_sc_hd__xnor2_1 _23625_ (.A(_03490_),
    .B(_03491_),
    .Y(_03492_));
 sky130_fd_sc_hd__xnor2_2 _23626_ (.A(_03489_),
    .B(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__nand2_1 _23627_ (.A(_03426_),
    .B(_03427_),
    .Y(_03494_));
 sky130_fd_sc_hd__nor2_1 _23628_ (.A(_03426_),
    .B(_03427_),
    .Y(_03495_));
 sky130_fd_sc_hd__a31o_1 _23629_ (.A1(net4641),
    .A2(net4940),
    .A3(_03494_),
    .B1(_03495_),
    .X(_03496_));
 sky130_fd_sc_hd__nand2_1 _23630_ (.A(net4703),
    .B(net4846),
    .Y(_03497_));
 sky130_fd_sc_hd__nand2_1 _23631_ (.A(net4728),
    .B(net4822),
    .Y(_03498_));
 sky130_fd_sc_hd__xor2_1 _23632_ (.A(_03497_),
    .B(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__nand2_1 _23633_ (.A(net4748),
    .B(net4812),
    .Y(_03500_));
 sky130_fd_sc_hd__xor2_1 _23634_ (.A(_03499_),
    .B(_03500_),
    .X(_03501_));
 sky130_fd_sc_hd__xor2_1 _23635_ (.A(_03496_),
    .B(net2413),
    .X(_03502_));
 sky130_fd_sc_hd__xnor2_2 _23636_ (.A(_03493_),
    .B(_03502_),
    .Y(_03503_));
 sky130_fd_sc_hd__a21bo_1 _23637_ (.A1(_03417_),
    .A2(_03419_),
    .B1_N(_03415_),
    .X(_03504_));
 sky130_fd_sc_hd__o21ai_1 _23638_ (.A1(_03417_),
    .A2(_03419_),
    .B1(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__o21a_1 _23639_ (.A1(_03432_),
    .A2(_03437_),
    .B1(_03430_),
    .X(_03506_));
 sky130_fd_sc_hd__a21o_1 _23640_ (.A1(_03432_),
    .A2(_03437_),
    .B1(_03506_),
    .X(_03507_));
 sky130_fd_sc_hd__xnor2_1 _23641_ (.A(net1666),
    .B(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__xnor2_2 _23642_ (.A(_03503_),
    .B(_03508_),
    .Y(_03509_));
 sky130_fd_sc_hd__a21bo_1 _23643_ (.A1(_03410_),
    .A2(_03421_),
    .B1_N(net1384),
    .X(_03510_));
 sky130_fd_sc_hd__o21ai_1 _23644_ (.A1(_03410_),
    .A2(_03421_),
    .B1(_03510_),
    .Y(_03511_));
 sky130_fd_sc_hd__nand2_1 _23645_ (.A(net4558),
    .B(net5023),
    .Y(_03512_));
 sky130_fd_sc_hd__nand2_1 _23646_ (.A(net4530),
    .B(net5078),
    .Y(_03513_));
 sky130_fd_sc_hd__nand2_1 _23647_ (.A(net4548),
    .B(net5052),
    .Y(_03514_));
 sky130_fd_sc_hd__xor2_1 _23648_ (.A(_03513_),
    .B(_03514_),
    .X(_03515_));
 sky130_fd_sc_hd__xnor2_1 _23649_ (.A(_03512_),
    .B(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__o21ai_1 _23650_ (.A1(net3748),
    .A2(_03395_),
    .B1(_03394_),
    .Y(_03517_));
 sky130_fd_sc_hd__a21bo_1 _23651_ (.A1(net3748),
    .A2(_03395_),
    .B1_N(_03517_),
    .X(_03518_));
 sky130_fd_sc_hd__xor2_1 _23652_ (.A(net5154),
    .B(net5120),
    .X(_03519_));
 sky130_fd_sc_hd__nand2_1 _23653_ (.A(net4495),
    .B(_03519_),
    .Y(_03520_));
 sky130_fd_sc_hd__nand2_1 _23654_ (.A(net5094),
    .B(net4511),
    .Y(_03521_));
 sky130_fd_sc_hd__xnor2_2 _23655_ (.A(_03520_),
    .B(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__xnor2_1 _23656_ (.A(_03518_),
    .B(_03522_),
    .Y(_03523_));
 sky130_fd_sc_hd__xnor2_1 _23657_ (.A(_03516_),
    .B(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__a21oi_1 _23658_ (.A1(_03397_),
    .A2(_03406_),
    .B1(_03405_),
    .Y(_03525_));
 sky130_fd_sc_hd__nand2_1 _23659_ (.A(net4615),
    .B(net4934),
    .Y(_03526_));
 sky130_fd_sc_hd__nand2_1 _23660_ (.A(net4576),
    .B(net4998),
    .Y(_03527_));
 sky130_fd_sc_hd__nand2_1 _23661_ (.A(net4598),
    .B(net4964),
    .Y(_03528_));
 sky130_fd_sc_hd__xnor2_1 _23662_ (.A(_03527_),
    .B(_03528_),
    .Y(_03529_));
 sky130_fd_sc_hd__xnor2_1 _23663_ (.A(_03526_),
    .B(_03529_),
    .Y(_03530_));
 sky130_fd_sc_hd__o21a_1 _23664_ (.A1(_03411_),
    .A2(_03412_),
    .B1(_03413_),
    .X(_03531_));
 sky130_fd_sc_hd__a21oi_2 _23665_ (.A1(_03411_),
    .A2(_03412_),
    .B1(_03531_),
    .Y(_03532_));
 sky130_fd_sc_hd__o21a_1 _23666_ (.A1(_03400_),
    .A2(_03401_),
    .B1(_03402_),
    .X(_03533_));
 sky130_fd_sc_hd__a21oi_2 _23667_ (.A1(_03400_),
    .A2(_03401_),
    .B1(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__xnor2_1 _23668_ (.A(_03532_),
    .B(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__xnor2_1 _23669_ (.A(_03530_),
    .B(_03535_),
    .Y(_03536_));
 sky130_fd_sc_hd__nor2_1 _23670_ (.A(_03525_),
    .B(_03536_),
    .Y(_03537_));
 sky130_fd_sc_hd__nand2_1 _23671_ (.A(_03525_),
    .B(_03536_),
    .Y(_03538_));
 sky130_fd_sc_hd__or2b_1 _23672_ (.A(_03537_),
    .B_N(_03538_),
    .X(_03539_));
 sky130_fd_sc_hd__xnor2_1 _23673_ (.A(_03524_),
    .B(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hd__xnor2_1 _23674_ (.A(net1019),
    .B(net1018),
    .Y(_03541_));
 sky130_fd_sc_hd__xnor2_2 _23675_ (.A(_03509_),
    .B(_03541_),
    .Y(_03542_));
 sky130_fd_sc_hd__a21o_1 _23676_ (.A1(_03423_),
    .A2(_03447_),
    .B1(_03446_),
    .X(_03543_));
 sky130_fd_sc_hd__o21a_1 _23677_ (.A1(_03441_),
    .A2(_03443_),
    .B1(_03439_),
    .X(_03544_));
 sky130_fd_sc_hd__a21o_1 _23678_ (.A1(_03441_),
    .A2(_03443_),
    .B1(_03544_),
    .X(_03545_));
 sky130_fd_sc_hd__a21o_1 _23679_ (.A1(_03455_),
    .A2(_03457_),
    .B1(_03458_),
    .X(_03546_));
 sky130_fd_sc_hd__o21ai_1 _23680_ (.A1(_03455_),
    .A2(_03457_),
    .B1(_03546_),
    .Y(_03547_));
 sky130_fd_sc_hd__or2_1 _23681_ (.A(net4768),
    .B(net3746),
    .X(_03548_));
 sky130_fd_sc_hd__o21a_1 _23682_ (.A1(_03433_),
    .A2(_03434_),
    .B1(_03435_),
    .X(_03549_));
 sky130_fd_sc_hd__a21oi_1 _23683_ (.A1(_03433_),
    .A2(_03434_),
    .B1(_03549_),
    .Y(_03550_));
 sky130_fd_sc_hd__xnor2_1 _23684_ (.A(_03548_),
    .B(_03550_),
    .Y(_03551_));
 sky130_fd_sc_hd__nor2_1 _23685_ (.A(_03547_),
    .B(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__nand2_1 _23686_ (.A(_03547_),
    .B(_03551_),
    .Y(_03553_));
 sky130_fd_sc_hd__and2b_1 _23687_ (.A_N(_03552_),
    .B(_03553_),
    .X(_03554_));
 sky130_fd_sc_hd__xnor2_1 _23688_ (.A(net1165),
    .B(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__nor2_1 _23689_ (.A(net933),
    .B(_03555_),
    .Y(_03556_));
 sky130_fd_sc_hd__nand2_1 _23690_ (.A(net933),
    .B(_03555_),
    .Y(_03557_));
 sky130_fd_sc_hd__or2b_1 _23691_ (.A(_03556_),
    .B_N(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__xnor2_2 _23692_ (.A(_03542_),
    .B(_03558_),
    .Y(_03559_));
 sky130_fd_sc_hd__o21a_1 _23693_ (.A1(_03451_),
    .A2(_03461_),
    .B1(_03449_),
    .X(_03560_));
 sky130_fd_sc_hd__a21o_1 _23694_ (.A1(_03451_),
    .A2(_03461_),
    .B1(_03560_),
    .X(_03561_));
 sky130_fd_sc_hd__or2_1 _23695_ (.A(_03453_),
    .B(_03460_),
    .X(_03562_));
 sky130_fd_sc_hd__xor2_1 _23696_ (.A(net744),
    .B(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__xnor2_1 _23697_ (.A(_03559_),
    .B(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__xnor2_1 _23698_ (.A(net639),
    .B(_03564_),
    .Y(_03565_));
 sky130_fd_sc_hd__xnor2_1 _23699_ (.A(_03486_),
    .B(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__inv_2 _23700_ (.A(\pid_q.curr_error[2] ),
    .Y(_03567_));
 sky130_fd_sc_hd__a21o_1 _23701_ (.A1(_03475_),
    .A2(_03476_),
    .B1(_03567_),
    .X(_03568_));
 sky130_fd_sc_hd__inv_2 _23702_ (.A(\pid_q.prev_error[2] ),
    .Y(_03569_));
 sky130_fd_sc_hd__a31o_1 _23703_ (.A1(_03567_),
    .A2(_03475_),
    .A3(_03476_),
    .B1(_03569_),
    .X(_03570_));
 sky130_fd_sc_hd__and2_1 _23704_ (.A(_03568_),
    .B(_03570_),
    .X(_03571_));
 sky130_fd_sc_hd__xnor2_1 _23705_ (.A(\pid_q.prev_error[3] ),
    .B(\pid_q.curr_error[3] ),
    .Y(_03572_));
 sky130_fd_sc_hd__nand2_1 _23706_ (.A(_03571_),
    .B(_03572_),
    .Y(_03573_));
 sky130_fd_sc_hd__or2_1 _23707_ (.A(_03571_),
    .B(_03572_),
    .X(_03574_));
 sky130_fd_sc_hd__and3_1 _23708_ (.A(net7503),
    .B(_03573_),
    .C(_03574_),
    .X(_03575_));
 sky130_fd_sc_hd__a221o_1 _23709_ (.A1(net7527),
    .A2(_03485_),
    .B1(net467),
    .B2(net7468),
    .C1(net1663),
    .X(_03576_));
 sky130_fd_sc_hd__a22o_1 _23710_ (.A1(\pid_q.curr_int[3] ),
    .A2(net3062),
    .B1(net2029),
    .B2(_03576_),
    .X(_00668_));
 sky130_fd_sc_hd__inv_2 _23711_ (.A(\pid_q.prev_int[3] ),
    .Y(_03577_));
 sky130_fd_sc_hd__inv_2 _23712_ (.A(\pid_q.curr_int[3] ),
    .Y(_03578_));
 sky130_fd_sc_hd__o21a_1 _23713_ (.A1(_03577_),
    .A2(_03483_),
    .B1(_03578_),
    .X(_03579_));
 sky130_fd_sc_hd__a21o_1 _23714_ (.A1(_03577_),
    .A2(_03483_),
    .B1(_03579_),
    .X(_03580_));
 sky130_fd_sc_hd__xor2_1 _23715_ (.A(\pid_q.curr_int[4] ),
    .B(\pid_q.prev_int[4] ),
    .X(_03581_));
 sky130_fd_sc_hd__xnor2_1 _23716_ (.A(_03580_),
    .B(_03581_),
    .Y(_03582_));
 sky130_fd_sc_hd__and2b_1 _23717_ (.A_N(net639),
    .B(_03564_),
    .X(_03583_));
 sky130_fd_sc_hd__a31o_1 _23718_ (.A1(net696),
    .A2(_03470_),
    .A3(_03472_),
    .B1(_03583_),
    .X(_03584_));
 sky130_fd_sc_hd__or2b_1 _23719_ (.A(_03564_),
    .B_N(net639),
    .X(_03585_));
 sky130_fd_sc_hd__nand2_1 _23720_ (.A(_03584_),
    .B(_03585_),
    .Y(_03586_));
 sky130_fd_sc_hd__o21ba_1 _23721_ (.A1(_03518_),
    .A2(_03522_),
    .B1_N(_03516_),
    .X(_03587_));
 sky130_fd_sc_hd__a21oi_2 _23722_ (.A1(_03518_),
    .A2(_03522_),
    .B1(_03587_),
    .Y(_03588_));
 sky130_fd_sc_hd__nand2_1 _23723_ (.A(net4600),
    .B(net4942),
    .Y(_03589_));
 sky130_fd_sc_hd__nand2_1 _23724_ (.A(net4562),
    .B(net4997),
    .Y(_03590_));
 sky130_fd_sc_hd__nand2_1 _23725_ (.A(net4587),
    .B(net4963),
    .Y(_03591_));
 sky130_fd_sc_hd__xnor2_1 _23726_ (.A(_03590_),
    .B(_03591_),
    .Y(_03592_));
 sky130_fd_sc_hd__xnor2_1 _23727_ (.A(_03589_),
    .B(_03592_),
    .Y(_03593_));
 sky130_fd_sc_hd__o21a_1 _23728_ (.A1(_03512_),
    .A2(_03514_),
    .B1(_03513_),
    .X(_03594_));
 sky130_fd_sc_hd__a21oi_2 _23729_ (.A1(_03512_),
    .A2(_03514_),
    .B1(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__o21a_1 _23730_ (.A1(_03526_),
    .A2(_03528_),
    .B1(_03527_),
    .X(_03596_));
 sky130_fd_sc_hd__a21oi_2 _23731_ (.A1(_03526_),
    .A2(_03528_),
    .B1(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__xnor2_1 _23732_ (.A(_03595_),
    .B(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hd__xnor2_1 _23733_ (.A(_03593_),
    .B(_03598_),
    .Y(_03599_));
 sky130_fd_sc_hd__nand2_1 _23734_ (.A(net5077),
    .B(net4508),
    .Y(_03600_));
 sky130_fd_sc_hd__nand2_1 _23735_ (.A(net4527),
    .B(net5051),
    .Y(_03601_));
 sky130_fd_sc_hd__nand2_1 _23736_ (.A(net4543),
    .B(net5031),
    .Y(_03602_));
 sky130_fd_sc_hd__xnor2_1 _23737_ (.A(_03601_),
    .B(_03602_),
    .Y(_03603_));
 sky130_fd_sc_hd__xnor2_1 _23738_ (.A(_03600_),
    .B(_03603_),
    .Y(_03604_));
 sky130_fd_sc_hd__inv_2 _23739_ (.A(net4504),
    .Y(_03605_));
 sky130_fd_sc_hd__o21a_1 _23740_ (.A1(net5120),
    .A2(net3744),
    .B1(net5155),
    .X(_03606_));
 sky130_fd_sc_hd__a21o_1 _23741_ (.A1(net5120),
    .A2(net3744),
    .B1(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__o31ai_1 _23742_ (.A1(net5146),
    .A2(net5122),
    .A3(net5097),
    .B1(net4482),
    .Y(_03608_));
 sky130_fd_sc_hd__a21o_1 _23743_ (.A1(net5096),
    .A2(_03607_),
    .B1(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__xnor2_1 _23744_ (.A(net2412),
    .B(_03609_),
    .Y(_03610_));
 sky130_fd_sc_hd__nor2_1 _23745_ (.A(net1662),
    .B(_03610_),
    .Y(_03611_));
 sky130_fd_sc_hd__nand2_1 _23746_ (.A(net1662),
    .B(_03610_),
    .Y(_03612_));
 sky130_fd_sc_hd__and2b_1 _23747_ (.A_N(_03611_),
    .B(_03612_),
    .X(_03613_));
 sky130_fd_sc_hd__xnor2_1 _23748_ (.A(_03588_),
    .B(_03613_),
    .Y(_03614_));
 sky130_fd_sc_hd__o21ai_1 _23749_ (.A1(_03524_),
    .A2(_03537_),
    .B1(_03538_),
    .Y(_03615_));
 sky130_fd_sc_hd__nand2_1 _23750_ (.A(net4729),
    .B(net4812),
    .Y(_03616_));
 sky130_fd_sc_hd__nand2_1 _23751_ (.A(net4674),
    .B(net4859),
    .Y(_03617_));
 sky130_fd_sc_hd__nand2_1 _23752_ (.A(net4703),
    .B(net4828),
    .Y(_03618_));
 sky130_fd_sc_hd__xnor2_1 _23753_ (.A(_03617_),
    .B(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__xnor2_2 _23754_ (.A(_03616_),
    .B(_03619_),
    .Y(_03620_));
 sky130_fd_sc_hd__o21ai_1 _23755_ (.A1(_03489_),
    .A2(_03491_),
    .B1(_03490_),
    .Y(_03621_));
 sky130_fd_sc_hd__a21bo_1 _23756_ (.A1(_03489_),
    .A2(_03491_),
    .B1_N(_03621_),
    .X(_03622_));
 sky130_fd_sc_hd__nand2_1 _23757_ (.A(net4665),
    .B(net4875),
    .Y(_03623_));
 sky130_fd_sc_hd__nand2_1 _23758_ (.A(net4616),
    .B(net4922),
    .Y(_03624_));
 sky130_fd_sc_hd__nand2_1 _23759_ (.A(net4636),
    .B(net4899),
    .Y(_03625_));
 sky130_fd_sc_hd__xnor2_1 _23760_ (.A(_03624_),
    .B(_03625_),
    .Y(_03626_));
 sky130_fd_sc_hd__xnor2_2 _23761_ (.A(_03623_),
    .B(_03626_),
    .Y(_03627_));
 sky130_fd_sc_hd__xnor2_1 _23762_ (.A(_03622_),
    .B(_03627_),
    .Y(_03628_));
 sky130_fd_sc_hd__xnor2_2 _23763_ (.A(_03620_),
    .B(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__a21bo_1 _23764_ (.A1(_03532_),
    .A2(_03534_),
    .B1_N(_03530_),
    .X(_03630_));
 sky130_fd_sc_hd__o21ai_1 _23765_ (.A1(_03532_),
    .A2(_03534_),
    .B1(_03630_),
    .Y(_03631_));
 sky130_fd_sc_hd__o21ba_1 _23766_ (.A1(_03493_),
    .A2(net2413),
    .B1_N(_03496_),
    .X(_03632_));
 sky130_fd_sc_hd__a21o_1 _23767_ (.A1(_03493_),
    .A2(net2413),
    .B1(_03632_),
    .X(_03633_));
 sky130_fd_sc_hd__and2_1 _23768_ (.A(net1661),
    .B(_03633_),
    .X(_03634_));
 sky130_fd_sc_hd__or2_1 _23769_ (.A(net1661),
    .B(_03633_),
    .X(_03635_));
 sky130_fd_sc_hd__or2b_1 _23770_ (.A(_03634_),
    .B_N(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__xnor2_2 _23771_ (.A(_03629_),
    .B(_03636_),
    .Y(_03637_));
 sky130_fd_sc_hd__xor2_1 _23772_ (.A(net1164),
    .B(_03637_),
    .X(_03638_));
 sky130_fd_sc_hd__xnor2_1 _23773_ (.A(_03614_),
    .B(_03638_),
    .Y(_03639_));
 sky130_fd_sc_hd__a21bo_1 _23774_ (.A1(net1019),
    .A2(net1018),
    .B1_N(_03509_),
    .X(_03640_));
 sky130_fd_sc_hd__o21a_1 _23775_ (.A1(net1019),
    .A2(net1018),
    .B1(_03640_),
    .X(_03641_));
 sky130_fd_sc_hd__o21a_1 _23776_ (.A1(net1666),
    .A2(_03507_),
    .B1(_03503_),
    .X(_03642_));
 sky130_fd_sc_hd__a21o_1 _23777_ (.A1(net1666),
    .A2(_03507_),
    .B1(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__and3_1 _23778_ (.A(net4708),
    .B(net4729),
    .C(_03372_),
    .X(_03644_));
 sky130_fd_sc_hd__xnor2_1 _23779_ (.A(net4796),
    .B(net3049),
    .Y(_03645_));
 sky130_fd_sc_hd__a21oi_1 _23780_ (.A1(net4810),
    .A2(_03499_),
    .B1(net3049),
    .Y(_03646_));
 sky130_fd_sc_hd__mux2_1 _23781_ (.A0(_03645_),
    .A1(_03646_),
    .S(net4748),
    .X(_03647_));
 sky130_fd_sc_hd__and2b_1 _23782_ (.A_N(_03548_),
    .B(_03550_),
    .X(_03648_));
 sky130_fd_sc_hd__xnor2_1 _23783_ (.A(_03647_),
    .B(_03648_),
    .Y(_03649_));
 sky130_fd_sc_hd__xnor2_2 _23784_ (.A(net1163),
    .B(_03649_),
    .Y(_03650_));
 sky130_fd_sc_hd__xnor2_1 _23785_ (.A(_03641_),
    .B(_03650_),
    .Y(_03651_));
 sky130_fd_sc_hd__xnor2_2 _23786_ (.A(net855),
    .B(_03651_),
    .Y(_03652_));
 sky130_fd_sc_hd__a21oi_1 _23787_ (.A1(_03542_),
    .A2(_03557_),
    .B1(_03556_),
    .Y(_03653_));
 sky130_fd_sc_hd__a21oi_1 _23788_ (.A1(net1165),
    .A2(_03553_),
    .B1(_03552_),
    .Y(_03654_));
 sky130_fd_sc_hd__xnor2_1 _23789_ (.A(_03653_),
    .B(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__xnor2_2 _23790_ (.A(_03652_),
    .B(_03655_),
    .Y(_03656_));
 sky130_fd_sc_hd__o21a_1 _23791_ (.A1(net744),
    .A2(_03559_),
    .B1(_03562_),
    .X(_03657_));
 sky130_fd_sc_hd__a21oi_1 _23792_ (.A1(net744),
    .A2(_03559_),
    .B1(_03657_),
    .Y(_03658_));
 sky130_fd_sc_hd__xor2_1 _23793_ (.A(_03656_),
    .B(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__xnor2_1 _23794_ (.A(_03586_),
    .B(_03659_),
    .Y(_03660_));
 sky130_fd_sc_hd__inv_2 _23795_ (.A(\pid_q.curr_error[3] ),
    .Y(_03661_));
 sky130_fd_sc_hd__inv_2 _23796_ (.A(\pid_q.prev_error[3] ),
    .Y(_03662_));
 sky130_fd_sc_hd__a31o_1 _23797_ (.A1(_03661_),
    .A2(_03568_),
    .A3(_03570_),
    .B1(_03662_),
    .X(_03663_));
 sky130_fd_sc_hd__o21a_1 _23798_ (.A1(_03661_),
    .A2(_03571_),
    .B1(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__xnor2_1 _23799_ (.A(\pid_q.prev_error[4] ),
    .B(\pid_q.curr_error[4] ),
    .Y(_03665_));
 sky130_fd_sc_hd__nand2_1 _23800_ (.A(_03664_),
    .B(_03665_),
    .Y(_03666_));
 sky130_fd_sc_hd__or2_1 _23801_ (.A(_03664_),
    .B(_03665_),
    .X(_03667_));
 sky130_fd_sc_hd__and3_1 _23802_ (.A(net7503),
    .B(_03666_),
    .C(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__a221o_1 _23803_ (.A1(net7527),
    .A2(_03582_),
    .B1(net463),
    .B2(net7468),
    .C1(net1381),
    .X(_03669_));
 sky130_fd_sc_hd__a22o_1 _23804_ (.A1(\pid_q.curr_int[4] ),
    .A2(net3062),
    .B1(net2028),
    .B2(_03669_),
    .X(_00669_));
 sky130_fd_sc_hd__inv_2 _23805_ (.A(\pid_q.prev_int[4] ),
    .Y(_03670_));
 sky130_fd_sc_hd__inv_2 _23806_ (.A(\pid_q.curr_int[4] ),
    .Y(_03671_));
 sky130_fd_sc_hd__o21a_1 _23807_ (.A1(_03670_),
    .A2(_03580_),
    .B1(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__a21o_1 _23808_ (.A1(_03670_),
    .A2(_03580_),
    .B1(_03672_),
    .X(_03673_));
 sky130_fd_sc_hd__xor2_1 _23809_ (.A(\pid_q.curr_int[5] ),
    .B(\pid_q.prev_int[5] ),
    .X(_03674_));
 sky130_fd_sc_hd__xnor2_1 _23810_ (.A(_03673_),
    .B(_03674_),
    .Y(_03675_));
 sky130_fd_sc_hd__a21o_1 _23811_ (.A1(_03584_),
    .A2(_03585_),
    .B1(_03658_),
    .X(_03676_));
 sky130_fd_sc_hd__and3_1 _23812_ (.A(_03584_),
    .B(_03585_),
    .C(_03658_),
    .X(_03677_));
 sky130_fd_sc_hd__a21o_1 _23813_ (.A1(_03656_),
    .A2(_03676_),
    .B1(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__a21o_1 _23814_ (.A1(_03652_),
    .A2(_03654_),
    .B1(_03653_),
    .X(_03679_));
 sky130_fd_sc_hd__or2_1 _23815_ (.A(_03652_),
    .B(_03654_),
    .X(_03680_));
 sky130_fd_sc_hd__nand2_1 _23816_ (.A(net4573),
    .B(net4941),
    .Y(_03681_));
 sky130_fd_sc_hd__nand2_1 _23817_ (.A(net4542),
    .B(net4991),
    .Y(_03682_));
 sky130_fd_sc_hd__nand2_1 _23818_ (.A(net4560),
    .B(net4957),
    .Y(_03683_));
 sky130_fd_sc_hd__xnor2_1 _23819_ (.A(_03682_),
    .B(_03683_),
    .Y(_03684_));
 sky130_fd_sc_hd__xnor2_1 _23820_ (.A(_03681_),
    .B(_03684_),
    .Y(_03685_));
 sky130_fd_sc_hd__nand2_1 _23821_ (.A(_03600_),
    .B(_03602_),
    .Y(_03686_));
 sky130_fd_sc_hd__nor2_1 _23822_ (.A(_03600_),
    .B(_03602_),
    .Y(_03687_));
 sky130_fd_sc_hd__a31o_1 _23823_ (.A1(net4527),
    .A2(net5057),
    .A3(_03686_),
    .B1(_03687_),
    .X(_03688_));
 sky130_fd_sc_hd__nand2_1 _23824_ (.A(_03589_),
    .B(_03591_),
    .Y(_03689_));
 sky130_fd_sc_hd__nor2_1 _23825_ (.A(_03589_),
    .B(_03591_),
    .Y(_03690_));
 sky130_fd_sc_hd__a31o_1 _23826_ (.A1(net4562),
    .A2(net4997),
    .A3(_03689_),
    .B1(_03690_),
    .X(_03691_));
 sky130_fd_sc_hd__xnor2_1 _23827_ (.A(_03688_),
    .B(_03691_),
    .Y(_03692_));
 sky130_fd_sc_hd__xnor2_1 _23828_ (.A(_03685_),
    .B(_03692_),
    .Y(_03693_));
 sky130_fd_sc_hd__nand2_2 _23829_ (.A(net5066),
    .B(net4483),
    .Y(_03694_));
 sky130_fd_sc_hd__nand2_1 _23830_ (.A(net4526),
    .B(net5020),
    .Y(_03695_));
 sky130_fd_sc_hd__nand2_1 _23831_ (.A(net5036),
    .B(net4499),
    .Y(_03696_));
 sky130_fd_sc_hd__xnor2_1 _23832_ (.A(_03695_),
    .B(_03696_),
    .Y(_03697_));
 sky130_fd_sc_hd__xnor2_2 _23833_ (.A(_03694_),
    .B(_03697_),
    .Y(_03698_));
 sky130_fd_sc_hd__a21oi_4 _23834_ (.A1(net5149),
    .A2(net3749),
    .B1(net3743),
    .Y(_03699_));
 sky130_fd_sc_hd__xnor2_2 _23835_ (.A(_03698_),
    .B(_03699_),
    .Y(_03700_));
 sky130_fd_sc_hd__nand2_1 _23836_ (.A(net5121),
    .B(net5095),
    .Y(_03701_));
 sky130_fd_sc_hd__and3_1 _23837_ (.A(net5096),
    .B(net3744),
    .C(_03519_),
    .X(_03702_));
 sky130_fd_sc_hd__nor2_1 _23838_ (.A(net5121),
    .B(net5095),
    .Y(_03703_));
 sky130_fd_sc_hd__o21ba_1 _23839_ (.A1(net2412),
    .A2(_03703_),
    .B1_N(net5155),
    .X(_03704_));
 sky130_fd_sc_hd__inv_2 _23840_ (.A(net4490),
    .Y(_03705_));
 sky130_fd_sc_hd__a2111oi_2 _23841_ (.A1(_03701_),
    .A2(net2412),
    .B1(_03702_),
    .C1(_03704_),
    .D1(net3741),
    .Y(_03706_));
 sky130_fd_sc_hd__xor2_1 _23842_ (.A(_03700_),
    .B(_03706_),
    .X(_03707_));
 sky130_fd_sc_hd__xnor2_1 _23843_ (.A(net1660),
    .B(_03707_),
    .Y(_03708_));
 sky130_fd_sc_hd__nand2_1 _23844_ (.A(net4688),
    .B(net4827),
    .Y(_03709_));
 sky130_fd_sc_hd__nand2_1 _23845_ (.A(net4669),
    .B(net4854),
    .Y(_03710_));
 sky130_fd_sc_hd__xor2_2 _23846_ (.A(_03709_),
    .B(_03710_),
    .X(_03711_));
 sky130_fd_sc_hd__nand2_1 _23847_ (.A(net4704),
    .B(net4811),
    .Y(_03712_));
 sky130_fd_sc_hd__xor2_2 _23848_ (.A(_03711_),
    .B(_03712_),
    .X(_03713_));
 sky130_fd_sc_hd__o21ai_1 _23849_ (.A1(_03623_),
    .A2(_03625_),
    .B1(_03624_),
    .Y(_03714_));
 sky130_fd_sc_hd__a21bo_1 _23850_ (.A1(_03623_),
    .A2(_03625_),
    .B1_N(_03714_),
    .X(_03715_));
 sky130_fd_sc_hd__nand2_1 _23851_ (.A(net4639),
    .B(net4868),
    .Y(_03716_));
 sky130_fd_sc_hd__nand2_1 _23852_ (.A(net4596),
    .B(net4921),
    .Y(_03717_));
 sky130_fd_sc_hd__nand2_1 _23853_ (.A(net4617),
    .B(net4891),
    .Y(_03718_));
 sky130_fd_sc_hd__xnor2_1 _23854_ (.A(_03717_),
    .B(_03718_),
    .Y(_03719_));
 sky130_fd_sc_hd__xnor2_1 _23855_ (.A(_03716_),
    .B(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__xnor2_1 _23856_ (.A(_03715_),
    .B(_03720_),
    .Y(_03721_));
 sky130_fd_sc_hd__xnor2_2 _23857_ (.A(_03713_),
    .B(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__o21a_1 _23858_ (.A1(_03622_),
    .A2(_03627_),
    .B1(_03620_),
    .X(_03723_));
 sky130_fd_sc_hd__a21o_1 _23859_ (.A1(_03622_),
    .A2(_03627_),
    .B1(_03723_),
    .X(_03724_));
 sky130_fd_sc_hd__a21bo_1 _23860_ (.A1(_03595_),
    .A2(_03597_),
    .B1_N(_03593_),
    .X(_03725_));
 sky130_fd_sc_hd__o21ai_1 _23861_ (.A1(_03595_),
    .A2(_03597_),
    .B1(_03725_),
    .Y(_03726_));
 sky130_fd_sc_hd__or2_1 _23862_ (.A(_03724_),
    .B(_03726_),
    .X(_03727_));
 sky130_fd_sc_hd__and2_1 _23863_ (.A(_03724_),
    .B(_03726_),
    .X(_03728_));
 sky130_fd_sc_hd__inv_2 _23864_ (.A(_03728_),
    .Y(_03729_));
 sky130_fd_sc_hd__nand2_1 _23865_ (.A(_03727_),
    .B(_03729_),
    .Y(_03730_));
 sky130_fd_sc_hd__xnor2_2 _23866_ (.A(_03722_),
    .B(_03730_),
    .Y(_03731_));
 sky130_fd_sc_hd__a21oi_2 _23867_ (.A1(_03588_),
    .A2(_03612_),
    .B1(_03611_),
    .Y(_03732_));
 sky130_fd_sc_hd__xnor2_1 _23868_ (.A(_03731_),
    .B(_03732_),
    .Y(_03733_));
 sky130_fd_sc_hd__xnor2_2 _23869_ (.A(net1162),
    .B(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__o21a_1 _23870_ (.A1(net1164),
    .A2(_03637_),
    .B1(_03614_),
    .X(_03735_));
 sky130_fd_sc_hd__a21o_1 _23871_ (.A1(net1164),
    .A2(_03637_),
    .B1(_03735_),
    .X(_03736_));
 sky130_fd_sc_hd__a21o_1 _23872_ (.A1(_03629_),
    .A2(_03635_),
    .B1(_03634_),
    .X(_03737_));
 sky130_fd_sc_hd__nand3_1 _23873_ (.A(net4674),
    .B(net4704),
    .C(_03373_),
    .Y(_03738_));
 sky130_fd_sc_hd__clkbuf_1 _23874_ (.A(net3747),
    .X(_03739_));
 sky130_fd_sc_hd__a21o_1 _23875_ (.A1(_03617_),
    .A2(_03618_),
    .B1(_03616_),
    .X(_03740_));
 sky130_fd_sc_hd__o21a_1 _23876_ (.A1(net4729),
    .A2(net3048),
    .B1(_03740_),
    .X(_03741_));
 sky130_fd_sc_hd__or3_1 _23877_ (.A(net4729),
    .B(net3747),
    .C(_03738_),
    .X(_03742_));
 sky130_fd_sc_hd__a21bo_1 _23878_ (.A1(_03738_),
    .A2(_03741_),
    .B1_N(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__or3b_1 _23879_ (.A(net4748),
    .B(_03739_),
    .C_N(net3049),
    .X(_03744_));
 sky130_fd_sc_hd__xor2_1 _23880_ (.A(_03743_),
    .B(_03744_),
    .X(_03745_));
 sky130_fd_sc_hd__xnor2_2 _23881_ (.A(_03737_),
    .B(_03745_),
    .Y(_03746_));
 sky130_fd_sc_hd__xnor2_1 _23882_ (.A(_03736_),
    .B(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__xnor2_1 _23883_ (.A(_03734_),
    .B(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__o21a_1 _23884_ (.A1(_03641_),
    .A2(_03650_),
    .B1(net855),
    .X(_03749_));
 sky130_fd_sc_hd__a21o_1 _23885_ (.A1(_03641_),
    .A2(_03650_),
    .B1(_03749_),
    .X(_03750_));
 sky130_fd_sc_hd__o21ba_1 _23886_ (.A1(net1163),
    .A2(_03647_),
    .B1_N(_03648_),
    .X(_03751_));
 sky130_fd_sc_hd__a21oi_1 _23887_ (.A1(net1163),
    .A2(_03647_),
    .B1(_03751_),
    .Y(_03752_));
 sky130_fd_sc_hd__nand2_1 _23888_ (.A(_03750_),
    .B(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__inv_2 _23889_ (.A(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__nor2_1 _23890_ (.A(_03750_),
    .B(_03752_),
    .Y(_03755_));
 sky130_fd_sc_hd__nor2_1 _23891_ (.A(_03754_),
    .B(_03755_),
    .Y(_03756_));
 sky130_fd_sc_hd__xnor2_1 _23892_ (.A(_03748_),
    .B(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__a21oi_1 _23893_ (.A1(_03679_),
    .A2(_03680_),
    .B1(_03757_),
    .Y(_03758_));
 sky130_fd_sc_hd__and3_1 _23894_ (.A(_03757_),
    .B(_03679_),
    .C(_03680_),
    .X(_03759_));
 sky130_fd_sc_hd__nor2_1 _23895_ (.A(_03758_),
    .B(_03759_),
    .Y(_03760_));
 sky130_fd_sc_hd__xor2_1 _23896_ (.A(_03678_),
    .B(_03760_),
    .X(_03761_));
 sky130_fd_sc_hd__inv_2 _23897_ (.A(\pid_q.curr_error[4] ),
    .Y(_03762_));
 sky130_fd_sc_hd__o21ba_1 _23898_ (.A1(_03762_),
    .A2(_03664_),
    .B1_N(\pid_q.prev_error[4] ),
    .X(_03763_));
 sky130_fd_sc_hd__a21o_1 _23899_ (.A1(_03762_),
    .A2(_03664_),
    .B1(_03763_),
    .X(_03764_));
 sky130_fd_sc_hd__xnor2_1 _23900_ (.A(\pid_q.prev_error[5] ),
    .B(\pid_q.curr_error[5] ),
    .Y(_03765_));
 sky130_fd_sc_hd__nand2_1 _23901_ (.A(_03764_),
    .B(_03765_),
    .Y(_03766_));
 sky130_fd_sc_hd__or2_1 _23902_ (.A(_03764_),
    .B(_03765_),
    .X(_03767_));
 sky130_fd_sc_hd__and3_1 _23903_ (.A(net7504),
    .B(_03766_),
    .C(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__a221o_1 _23904_ (.A1(net7526),
    .A2(_03675_),
    .B1(net408),
    .B2(net7466),
    .C1(net1016),
    .X(_03769_));
 sky130_fd_sc_hd__a22o_1 _23905_ (.A1(\pid_q.curr_int[5] ),
    .A2(net3061),
    .B1(net2027),
    .B2(_03769_),
    .X(_00670_));
 sky130_fd_sc_hd__inv_2 _23906_ (.A(\pid_q.prev_int[5] ),
    .Y(_03770_));
 sky130_fd_sc_hd__inv_2 _23907_ (.A(\pid_q.curr_int[5] ),
    .Y(_03771_));
 sky130_fd_sc_hd__o21a_1 _23908_ (.A1(_03770_),
    .A2(_03673_),
    .B1(_03771_),
    .X(_03772_));
 sky130_fd_sc_hd__a21o_1 _23909_ (.A1(_03770_),
    .A2(_03673_),
    .B1(_03772_),
    .X(_03773_));
 sky130_fd_sc_hd__xor2_1 _23910_ (.A(\pid_q.curr_int[6] ),
    .B(\pid_q.prev_int[6] ),
    .X(_03774_));
 sky130_fd_sc_hd__xnor2_1 _23911_ (.A(_03773_),
    .B(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__inv_2 _23912_ (.A(_03759_),
    .Y(_03776_));
 sky130_fd_sc_hd__o21ai_1 _23913_ (.A1(_03656_),
    .A2(_03677_),
    .B1(_03676_),
    .Y(_03777_));
 sky130_fd_sc_hd__a21o_1 _23914_ (.A1(_03776_),
    .A2(_03777_),
    .B1(_03758_),
    .X(_03778_));
 sky130_fd_sc_hd__or2_1 _23915_ (.A(_03748_),
    .B(_03755_),
    .X(_03779_));
 sky130_fd_sc_hd__a21bo_1 _23916_ (.A1(_03731_),
    .A2(_03732_),
    .B1_N(net1162),
    .X(_03780_));
 sky130_fd_sc_hd__o21a_1 _23917_ (.A1(_03731_),
    .A2(_03732_),
    .B1(_03780_),
    .X(_03781_));
 sky130_fd_sc_hd__nand2_1 _23918_ (.A(net4611),
    .B(net4880),
    .Y(_03782_));
 sky130_fd_sc_hd__nand2_1 _23919_ (.A(net4572),
    .B(net4915),
    .Y(_03783_));
 sky130_fd_sc_hd__nand2_1 _23920_ (.A(net4592),
    .B(net4905),
    .Y(_03784_));
 sky130_fd_sc_hd__xnor2_1 _23921_ (.A(_03783_),
    .B(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__xnor2_1 _23922_ (.A(_03782_),
    .B(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__o21ai_1 _23923_ (.A1(_03716_),
    .A2(_03718_),
    .B1(_03717_),
    .Y(_03787_));
 sky130_fd_sc_hd__a21bo_1 _23924_ (.A1(_03716_),
    .A2(_03718_),
    .B1_N(_03787_),
    .X(_03788_));
 sky130_fd_sc_hd__nand2_1 _23925_ (.A(net4661),
    .B(net4830),
    .Y(_03789_));
 sky130_fd_sc_hd__nand2_1 _23926_ (.A(net4635),
    .B(net4855),
    .Y(_03790_));
 sky130_fd_sc_hd__xor2_2 _23927_ (.A(_03789_),
    .B(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__nand2_1 _23928_ (.A(net4676),
    .B(net4799),
    .Y(_03792_));
 sky130_fd_sc_hd__xor2_2 _23929_ (.A(_03791_),
    .B(_03792_),
    .X(_03793_));
 sky130_fd_sc_hd__xnor2_1 _23930_ (.A(_03788_),
    .B(_03793_),
    .Y(_03794_));
 sky130_fd_sc_hd__xnor2_1 _23931_ (.A(net2411),
    .B(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__o21ba_1 _23932_ (.A1(_03688_),
    .A2(_03691_),
    .B1_N(_03685_),
    .X(_03796_));
 sky130_fd_sc_hd__a21oi_1 _23933_ (.A1(_03688_),
    .A2(_03691_),
    .B1(_03796_),
    .Y(_03797_));
 sky130_fd_sc_hd__o21a_1 _23934_ (.A1(_03715_),
    .A2(_03720_),
    .B1(_03713_),
    .X(_03798_));
 sky130_fd_sc_hd__a21o_1 _23935_ (.A1(_03715_),
    .A2(_03720_),
    .B1(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__and2_1 _23936_ (.A(_03797_),
    .B(_03799_),
    .X(_03800_));
 sky130_fd_sc_hd__or2_1 _23937_ (.A(_03797_),
    .B(_03799_),
    .X(_03801_));
 sky130_fd_sc_hd__and2b_1 _23938_ (.A_N(_03800_),
    .B(_03801_),
    .X(_03802_));
 sky130_fd_sc_hd__xnor2_1 _23939_ (.A(_03795_),
    .B(_03802_),
    .Y(_03803_));
 sky130_fd_sc_hd__nand2_1 _23940_ (.A(_03701_),
    .B(_03698_),
    .Y(_03804_));
 sky130_fd_sc_hd__o2bb2a_1 _23941_ (.A1_N(net5155),
    .A2_N(_03804_),
    .B1(_03698_),
    .B2(_03703_),
    .X(_03805_));
 sky130_fd_sc_hd__nor2_1 _23942_ (.A(net3741),
    .B(_03805_),
    .Y(_03806_));
 sky130_fd_sc_hd__nand2_2 _23943_ (.A(net4559),
    .B(net4951),
    .Y(_03807_));
 sky130_fd_sc_hd__nand2_1 _23944_ (.A(net4518),
    .B(net4986),
    .Y(_03808_));
 sky130_fd_sc_hd__nand2_1 _23945_ (.A(net4541),
    .B(net4972),
    .Y(_03809_));
 sky130_fd_sc_hd__xnor2_1 _23946_ (.A(_03808_),
    .B(_03809_),
    .Y(_03810_));
 sky130_fd_sc_hd__xnor2_2 _23947_ (.A(_03807_),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__o21a_1 _23948_ (.A1(_03694_),
    .A2(_03696_),
    .B1(_03695_),
    .X(_03812_));
 sky130_fd_sc_hd__a21oi_2 _23949_ (.A1(_03694_),
    .A2(_03696_),
    .B1(_03812_),
    .Y(_03813_));
 sky130_fd_sc_hd__o21a_1 _23950_ (.A1(_03681_),
    .A2(_03683_),
    .B1(_03682_),
    .X(_03814_));
 sky130_fd_sc_hd__a21oi_2 _23951_ (.A1(_03681_),
    .A2(_03683_),
    .B1(_03814_),
    .Y(_03815_));
 sky130_fd_sc_hd__xor2_1 _23952_ (.A(_03813_),
    .B(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__xnor2_2 _23953_ (.A(_03811_),
    .B(_03816_),
    .Y(_03817_));
 sky130_fd_sc_hd__nand2_1 _23954_ (.A(net5020),
    .B(net4499),
    .Y(_03818_));
 sky130_fd_sc_hd__xor2_1 _23955_ (.A(net5071),
    .B(net5036),
    .X(_03819_));
 sky130_fd_sc_hd__nand2_1 _23956_ (.A(net4488),
    .B(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hd__xor2_2 _23957_ (.A(_03818_),
    .B(_03820_),
    .X(_03821_));
 sky130_fd_sc_hd__xor2_2 _23958_ (.A(_03699_),
    .B(_03821_),
    .X(_03822_));
 sky130_fd_sc_hd__xor2_1 _23959_ (.A(_03817_),
    .B(_03822_),
    .X(_03823_));
 sky130_fd_sc_hd__xnor2_2 _23960_ (.A(_03806_),
    .B(_03823_),
    .Y(_03824_));
 sky130_fd_sc_hd__a21bo_1 _23961_ (.A1(_03700_),
    .A2(net1659),
    .B1_N(net1660),
    .X(_03825_));
 sky130_fd_sc_hd__o21ai_2 _23962_ (.A1(_03700_),
    .A2(net1659),
    .B1(_03825_),
    .Y(_03826_));
 sky130_fd_sc_hd__xnor2_1 _23963_ (.A(_03824_),
    .B(_03826_),
    .Y(_03827_));
 sky130_fd_sc_hd__xnor2_1 _23964_ (.A(_03803_),
    .B(_03827_),
    .Y(_03828_));
 sky130_fd_sc_hd__a21oi_1 _23965_ (.A1(_03722_),
    .A2(_03727_),
    .B1(_03728_),
    .Y(_03829_));
 sky130_fd_sc_hd__and3_1 _23966_ (.A(net4663),
    .B(net4688),
    .C(_03373_),
    .X(_03830_));
 sky130_fd_sc_hd__xnor2_1 _23967_ (.A(net3048),
    .B(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__a21o_1 _23968_ (.A1(net4811),
    .A2(_03711_),
    .B1(_03830_),
    .X(_03832_));
 sky130_fd_sc_hd__mux2_1 _23969_ (.A0(_03831_),
    .A1(_03832_),
    .S(net4704),
    .X(_03833_));
 sky130_fd_sc_hd__xnor2_1 _23970_ (.A(_03742_),
    .B(_03833_),
    .Y(_03834_));
 sky130_fd_sc_hd__xnor2_2 _23971_ (.A(net1161),
    .B(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__xnor2_1 _23972_ (.A(net932),
    .B(_03835_),
    .Y(_03836_));
 sky130_fd_sc_hd__xnor2_1 _23973_ (.A(net795),
    .B(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__a21bo_1 _23974_ (.A1(_03734_),
    .A2(_03746_),
    .B1_N(_03736_),
    .X(_03838_));
 sky130_fd_sc_hd__o21ai_1 _23975_ (.A1(_03734_),
    .A2(_03746_),
    .B1(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__o21a_1 _23976_ (.A1(_03737_),
    .A2(_03743_),
    .B1(_03744_),
    .X(_03840_));
 sky130_fd_sc_hd__a21o_1 _23977_ (.A1(_03737_),
    .A2(_03743_),
    .B1(_03840_),
    .X(_03841_));
 sky130_fd_sc_hd__nand2_1 _23978_ (.A(_03839_),
    .B(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__inv_2 _23979_ (.A(_03842_),
    .Y(_03843_));
 sky130_fd_sc_hd__nor2_1 _23980_ (.A(_03839_),
    .B(_03841_),
    .Y(_03844_));
 sky130_fd_sc_hd__nor2_1 _23981_ (.A(_03843_),
    .B(_03844_),
    .Y(_03845_));
 sky130_fd_sc_hd__xnor2_1 _23982_ (.A(_03837_),
    .B(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__a21o_1 _23983_ (.A1(_03753_),
    .A2(_03779_),
    .B1(net511),
    .X(_03847_));
 sky130_fd_sc_hd__inv_2 _23984_ (.A(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__and3_1 _23985_ (.A(_03753_),
    .B(net511),
    .C(_03779_),
    .X(_03849_));
 sky130_fd_sc_hd__nor2_1 _23986_ (.A(_03848_),
    .B(_03849_),
    .Y(_03850_));
 sky130_fd_sc_hd__xnor2_1 _23987_ (.A(_03778_),
    .B(_03850_),
    .Y(_03851_));
 sky130_fd_sc_hd__inv_2 _23988_ (.A(\pid_q.curr_error[5] ),
    .Y(_03852_));
 sky130_fd_sc_hd__o21ba_1 _23989_ (.A1(_03852_),
    .A2(_03764_),
    .B1_N(\pid_q.prev_error[5] ),
    .X(_03853_));
 sky130_fd_sc_hd__a21o_1 _23990_ (.A1(_03852_),
    .A2(_03764_),
    .B1(_03853_),
    .X(_03854_));
 sky130_fd_sc_hd__xnor2_1 _23991_ (.A(\pid_q.prev_error[6] ),
    .B(\pid_q.curr_error[6] ),
    .Y(_03855_));
 sky130_fd_sc_hd__nand2_1 _23992_ (.A(_03854_),
    .B(_03855_),
    .Y(_03856_));
 sky130_fd_sc_hd__or2_1 _23993_ (.A(_03854_),
    .B(_03855_),
    .X(_03857_));
 sky130_fd_sc_hd__and3_1 _23994_ (.A(net7504),
    .B(_03856_),
    .C(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__a221o_1 _23995_ (.A1(net7526),
    .A2(_03775_),
    .B1(net333),
    .B2(net7466),
    .C1(net854),
    .X(_03859_));
 sky130_fd_sc_hd__a22o_1 _23996_ (.A1(\pid_q.curr_int[6] ),
    .A2(net3061),
    .B1(net2027),
    .B2(_03859_),
    .X(_00671_));
 sky130_fd_sc_hd__inv_2 _23997_ (.A(\pid_q.prev_int[6] ),
    .Y(_03860_));
 sky130_fd_sc_hd__inv_2 _23998_ (.A(\pid_q.curr_int[6] ),
    .Y(_03861_));
 sky130_fd_sc_hd__o21a_1 _23999_ (.A1(_03860_),
    .A2(_03773_),
    .B1(_03861_),
    .X(_03862_));
 sky130_fd_sc_hd__a21o_1 _24000_ (.A1(_03860_),
    .A2(_03773_),
    .B1(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__xor2_1 _24001_ (.A(net5178),
    .B(\pid_q.prev_int[7] ),
    .X(_03864_));
 sky130_fd_sc_hd__xnor2_1 _24002_ (.A(net743),
    .B(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__a21oi_1 _24003_ (.A1(_03778_),
    .A2(_03847_),
    .B1(_03849_),
    .Y(_03866_));
 sky130_fd_sc_hd__nor2_1 _24004_ (.A(net795),
    .B(_03835_),
    .Y(_03867_));
 sky130_fd_sc_hd__nand2_1 _24005_ (.A(net795),
    .B(_03835_),
    .Y(_03868_));
 sky130_fd_sc_hd__o21ai_2 _24006_ (.A1(net932),
    .A2(_03867_),
    .B1(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__o21ai_1 _24007_ (.A1(net3749),
    .A2(_03821_),
    .B1(net5149),
    .Y(_03870_));
 sky130_fd_sc_hd__or2b_1 _24008_ (.A(_03703_),
    .B_N(_03821_),
    .X(_03871_));
 sky130_fd_sc_hd__a21oi_1 _24009_ (.A1(_03870_),
    .A2(_03871_),
    .B1(net3741),
    .Y(_03872_));
 sky130_fd_sc_hd__a21o_1 _24010_ (.A1(net5027),
    .A2(net4500),
    .B1(net5048),
    .X(_03873_));
 sky130_fd_sc_hd__and3_1 _24011_ (.A(net5048),
    .B(net5027),
    .C(net4500),
    .X(_03874_));
 sky130_fd_sc_hd__a21o_1 _24012_ (.A1(net5067),
    .A2(_03873_),
    .B1(_03874_),
    .X(_03875_));
 sky130_fd_sc_hd__nand2_1 _24013_ (.A(net4488),
    .B(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hd__o21ai_1 _24014_ (.A1(_03807_),
    .A2(_03809_),
    .B1(_03808_),
    .Y(_03877_));
 sky130_fd_sc_hd__a21bo_1 _24015_ (.A1(_03807_),
    .A2(_03809_),
    .B1_N(_03877_),
    .X(_03878_));
 sky130_fd_sc_hd__nand2_1 _24016_ (.A(net4987),
    .B(net4500),
    .Y(_03879_));
 sky130_fd_sc_hd__nand2_1 _24017_ (.A(net4519),
    .B(net4971),
    .Y(_03880_));
 sky130_fd_sc_hd__nand2_1 _24018_ (.A(net4534),
    .B(net4952),
    .Y(_03881_));
 sky130_fd_sc_hd__xnor2_1 _24019_ (.A(_03880_),
    .B(_03881_),
    .Y(_03882_));
 sky130_fd_sc_hd__xnor2_1 _24020_ (.A(_03879_),
    .B(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__xnor2_1 _24021_ (.A(_03878_),
    .B(_03883_),
    .Y(_03884_));
 sky130_fd_sc_hd__xnor2_2 _24022_ (.A(_03876_),
    .B(_03884_),
    .Y(_03885_));
 sky130_fd_sc_hd__xor2_1 _24023_ (.A(net5011),
    .B(_03819_),
    .X(_03886_));
 sky130_fd_sc_hd__nand2_2 _24024_ (.A(net4486),
    .B(_03886_),
    .Y(_03887_));
 sky130_fd_sc_hd__xor2_2 _24025_ (.A(_03699_),
    .B(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__xor2_1 _24026_ (.A(_03885_),
    .B(_03888_),
    .X(_03889_));
 sky130_fd_sc_hd__xnor2_1 _24027_ (.A(_03872_),
    .B(_03889_),
    .Y(_03890_));
 sky130_fd_sc_hd__a21o_1 _24028_ (.A1(_03817_),
    .A2(_03822_),
    .B1(_03806_),
    .X(_03891_));
 sky130_fd_sc_hd__o21ai_2 _24029_ (.A1(_03817_),
    .A2(_03822_),
    .B1(_03891_),
    .Y(_03892_));
 sky130_fd_sc_hd__nand2_2 _24030_ (.A(net4591),
    .B(net4881),
    .Y(_03893_));
 sky130_fd_sc_hd__nand2_1 _24031_ (.A(net4552),
    .B(net4911),
    .Y(_03894_));
 sky130_fd_sc_hd__nand2_1 _24032_ (.A(net4578),
    .B(net4906),
    .Y(_03895_));
 sky130_fd_sc_hd__xnor2_1 _24033_ (.A(_03894_),
    .B(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__xnor2_2 _24034_ (.A(_03893_),
    .B(_03896_),
    .Y(_03897_));
 sky130_fd_sc_hd__o21ai_1 _24035_ (.A1(_03782_),
    .A2(_03784_),
    .B1(_03783_),
    .Y(_03898_));
 sky130_fd_sc_hd__a21bo_1 _24036_ (.A1(_03782_),
    .A2(_03784_),
    .B1_N(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__nand2_1 _24037_ (.A(net4626),
    .B(net4834),
    .Y(_03900_));
 sky130_fd_sc_hd__nand2_1 _24038_ (.A(net4606),
    .B(net4851),
    .Y(_03901_));
 sky130_fd_sc_hd__xor2_1 _24039_ (.A(_03900_),
    .B(_03901_),
    .X(_03902_));
 sky130_fd_sc_hd__and3_1 _24040_ (.A(net4652),
    .B(net4815),
    .C(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__a21oi_1 _24041_ (.A1(net4652),
    .A2(net4801),
    .B1(_03902_),
    .Y(_03904_));
 sky130_fd_sc_hd__or2_1 _24042_ (.A(_03903_),
    .B(_03904_),
    .X(_03905_));
 sky130_fd_sc_hd__or2_1 _24043_ (.A(_03899_),
    .B(_03905_),
    .X(_03906_));
 sky130_fd_sc_hd__nand2_1 _24044_ (.A(_03899_),
    .B(_03905_),
    .Y(_03907_));
 sky130_fd_sc_hd__and2_1 _24045_ (.A(_03906_),
    .B(_03907_),
    .X(_03908_));
 sky130_fd_sc_hd__xnor2_2 _24046_ (.A(_03897_),
    .B(_03908_),
    .Y(_03909_));
 sky130_fd_sc_hd__a21bo_1 _24047_ (.A1(_03813_),
    .A2(_03815_),
    .B1_N(_03811_),
    .X(_03910_));
 sky130_fd_sc_hd__o21ai_1 _24048_ (.A1(_03813_),
    .A2(_03815_),
    .B1(_03910_),
    .Y(_03911_));
 sky130_fd_sc_hd__o21a_1 _24049_ (.A1(_03788_),
    .A2(_03793_),
    .B1(net2411),
    .X(_03912_));
 sky130_fd_sc_hd__a21o_1 _24050_ (.A1(_03788_),
    .A2(_03793_),
    .B1(_03912_),
    .X(_03913_));
 sky130_fd_sc_hd__nand2_1 _24051_ (.A(_03911_),
    .B(_03913_),
    .Y(_03914_));
 sky130_fd_sc_hd__inv_2 _24052_ (.A(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__nor2_1 _24053_ (.A(_03911_),
    .B(_03913_),
    .Y(_03916_));
 sky130_fd_sc_hd__nor2_1 _24054_ (.A(_03915_),
    .B(_03916_),
    .Y(_03917_));
 sky130_fd_sc_hd__xnor2_2 _24055_ (.A(_03909_),
    .B(_03917_),
    .Y(_03918_));
 sky130_fd_sc_hd__xor2_1 _24056_ (.A(_03892_),
    .B(_03918_),
    .X(_03919_));
 sky130_fd_sc_hd__xnor2_1 _24057_ (.A(_03890_),
    .B(_03919_),
    .Y(_03920_));
 sky130_fd_sc_hd__o21ba_1 _24058_ (.A1(_03824_),
    .A2(_03826_),
    .B1_N(_03803_),
    .X(_03921_));
 sky130_fd_sc_hd__a21o_1 _24059_ (.A1(_03824_),
    .A2(_03826_),
    .B1(_03921_),
    .X(_03922_));
 sky130_fd_sc_hd__o21a_1 _24060_ (.A1(_03795_),
    .A2(_03800_),
    .B1(_03801_),
    .X(_03923_));
 sky130_fd_sc_hd__and3_1 _24061_ (.A(net4640),
    .B(net4669),
    .C(_03372_),
    .X(_03924_));
 sky130_fd_sc_hd__xnor2_1 _24062_ (.A(net4790),
    .B(_03924_),
    .Y(_03925_));
 sky130_fd_sc_hd__a21oi_1 _24063_ (.A1(net4816),
    .A2(net3042),
    .B1(_03924_),
    .Y(_03926_));
 sky130_fd_sc_hd__mux2_1 _24064_ (.A0(_03925_),
    .A1(_03926_),
    .S(net4675),
    .X(_03927_));
 sky130_fd_sc_hd__or3b_1 _24065_ (.A(net4704),
    .B(net3747),
    .C_N(_03830_),
    .X(_03928_));
 sky130_fd_sc_hd__xor2_1 _24066_ (.A(_03927_),
    .B(_03928_),
    .X(_03929_));
 sky130_fd_sc_hd__xnor2_1 _24067_ (.A(net1160),
    .B(_03929_),
    .Y(_03930_));
 sky130_fd_sc_hd__inv_2 _24068_ (.A(_03930_),
    .Y(_03931_));
 sky130_fd_sc_hd__nand2_1 _24069_ (.A(_03922_),
    .B(_03931_),
    .Y(_03932_));
 sky130_fd_sc_hd__or2_1 _24070_ (.A(_03922_),
    .B(_03931_),
    .X(_03933_));
 sky130_fd_sc_hd__nand2_1 _24071_ (.A(_03932_),
    .B(_03933_),
    .Y(_03934_));
 sky130_fd_sc_hd__xnor2_1 _24072_ (.A(_03920_),
    .B(_03934_),
    .Y(_03935_));
 sky130_fd_sc_hd__a21bo_1 _24073_ (.A1(net1161),
    .A2(_03833_),
    .B1_N(_03742_),
    .X(_03936_));
 sky130_fd_sc_hd__o21ai_2 _24074_ (.A1(net1161),
    .A2(_03833_),
    .B1(_03936_),
    .Y(_03937_));
 sky130_fd_sc_hd__xor2_1 _24075_ (.A(_03935_),
    .B(_03937_),
    .X(_03938_));
 sky130_fd_sc_hd__xnor2_1 _24076_ (.A(_03869_),
    .B(_03938_),
    .Y(_03939_));
 sky130_fd_sc_hd__o21ai_1 _24077_ (.A1(_03837_),
    .A2(_03844_),
    .B1(_03842_),
    .Y(_03940_));
 sky130_fd_sc_hd__nand2_1 _24078_ (.A(net595),
    .B(net592),
    .Y(_03941_));
 sky130_fd_sc_hd__nor2_1 _24079_ (.A(net595),
    .B(net592),
    .Y(_03942_));
 sky130_fd_sc_hd__inv_2 _24080_ (.A(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__nand2_1 _24081_ (.A(_03941_),
    .B(_03943_),
    .Y(_03944_));
 sky130_fd_sc_hd__xnor2_1 _24082_ (.A(net376),
    .B(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__inv_2 _24083_ (.A(\pid_q.curr_error[6] ),
    .Y(_03946_));
 sky130_fd_sc_hd__o21ba_1 _24084_ (.A1(_03946_),
    .A2(_03854_),
    .B1_N(\pid_q.prev_error[6] ),
    .X(_03947_));
 sky130_fd_sc_hd__a21o_1 _24085_ (.A1(_03946_),
    .A2(_03854_),
    .B1(_03947_),
    .X(_03948_));
 sky130_fd_sc_hd__xnor2_1 _24086_ (.A(\pid_q.prev_error[7] ),
    .B(\pid_q.curr_error[7] ),
    .Y(_03949_));
 sky130_fd_sc_hd__nand2_1 _24087_ (.A(_03948_),
    .B(_03949_),
    .Y(_03950_));
 sky130_fd_sc_hd__or2_1 _24088_ (.A(_03948_),
    .B(_03949_),
    .X(_03951_));
 sky130_fd_sc_hd__and3_1 _24089_ (.A(net7505),
    .B(_03950_),
    .C(_03951_),
    .X(_03952_));
 sky130_fd_sc_hd__a221o_1 _24090_ (.A1(net7523),
    .A2(_03865_),
    .B1(net329),
    .B2(net7462),
    .C1(net741),
    .X(_03953_));
 sky130_fd_sc_hd__a22o_1 _24091_ (.A1(net5178),
    .A2(net3063),
    .B1(net2029),
    .B2(_03953_),
    .X(_00672_));
 sky130_fd_sc_hd__inv_2 _24092_ (.A(\pid_q.prev_int[7] ),
    .Y(_03954_));
 sky130_fd_sc_hd__inv_2 _24093_ (.A(net5178),
    .Y(_03955_));
 sky130_fd_sc_hd__o21a_1 _24094_ (.A1(_03954_),
    .A2(net743),
    .B1(_03955_),
    .X(_03956_));
 sky130_fd_sc_hd__a21o_1 _24095_ (.A1(_03954_),
    .A2(net743),
    .B1(_03956_),
    .X(_03957_));
 sky130_fd_sc_hd__xor2_1 _24096_ (.A(\pid_q.curr_int[8] ),
    .B(\pid_q.prev_int[8] ),
    .X(_03958_));
 sky130_fd_sc_hd__xnor2_1 _24097_ (.A(_03957_),
    .B(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__or2_1 _24098_ (.A(net376),
    .B(_03942_),
    .X(_03960_));
 sky130_fd_sc_hd__nand2_1 _24099_ (.A(_03941_),
    .B(_03960_),
    .Y(_03961_));
 sky130_fd_sc_hd__and4_1 _24100_ (.A(net5149),
    .B(net4483),
    .C(net3749),
    .D(_03886_),
    .X(_03962_));
 sky130_fd_sc_hd__a21oi_1 _24101_ (.A1(net3743),
    .A2(_03887_),
    .B1(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__nand2_2 _24102_ (.A(net4980),
    .B(net4484),
    .Y(_03964_));
 sky130_fd_sc_hd__nand2_1 _24103_ (.A(net4521),
    .B(net4953),
    .Y(_03965_));
 sky130_fd_sc_hd__nand2_1 _24104_ (.A(net4970),
    .B(net4501),
    .Y(_03966_));
 sky130_fd_sc_hd__xnor2_1 _24105_ (.A(_03965_),
    .B(_03966_),
    .Y(_03967_));
 sky130_fd_sc_hd__xnor2_2 _24106_ (.A(_03964_),
    .B(_03967_),
    .Y(_03968_));
 sky130_fd_sc_hd__o21ai_1 _24107_ (.A1(net5059),
    .A2(net5028),
    .B1(net5075),
    .Y(_03969_));
 sky130_fd_sc_hd__nand2_1 _24108_ (.A(net5059),
    .B(net5028),
    .Y(_03970_));
 sky130_fd_sc_hd__a21oi_1 _24109_ (.A1(_03969_),
    .A2(_03970_),
    .B1(net3742),
    .Y(_03971_));
 sky130_fd_sc_hd__o21a_1 _24110_ (.A1(_03879_),
    .A2(_03881_),
    .B1(_03880_),
    .X(_03972_));
 sky130_fd_sc_hd__a21oi_2 _24111_ (.A1(_03879_),
    .A2(_03881_),
    .B1(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__xnor2_1 _24112_ (.A(net3040),
    .B(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__xnor2_2 _24113_ (.A(_03968_),
    .B(_03974_),
    .Y(_03975_));
 sky130_fd_sc_hd__xnor2_2 _24114_ (.A(net2025),
    .B(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__o21ba_1 _24115_ (.A1(_03885_),
    .A2(_03888_),
    .B1_N(_03872_),
    .X(_03977_));
 sky130_fd_sc_hd__a21o_1 _24116_ (.A1(_03885_),
    .A2(_03888_),
    .B1(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__nand2_1 _24117_ (.A(net4590),
    .B(net4852),
    .Y(_03979_));
 sky130_fd_sc_hd__nand2_1 _24118_ (.A(net4604),
    .B(net4835),
    .Y(_03980_));
 sky130_fd_sc_hd__xor2_2 _24119_ (.A(_03979_),
    .B(_03980_),
    .X(_03981_));
 sky130_fd_sc_hd__nand2_1 _24120_ (.A(net4624),
    .B(net4802),
    .Y(_03982_));
 sky130_fd_sc_hd__xnor2_2 _24121_ (.A(_03981_),
    .B(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hd__o21ai_1 _24122_ (.A1(_03893_),
    .A2(_03895_),
    .B1(_03894_),
    .Y(_03984_));
 sky130_fd_sc_hd__a21bo_1 _24123_ (.A1(_03893_),
    .A2(_03895_),
    .B1_N(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__nand2_1 _24124_ (.A(net4579),
    .B(net4866),
    .Y(_03986_));
 sky130_fd_sc_hd__nand2_1 _24125_ (.A(net4534),
    .B(net4928),
    .Y(_03987_));
 sky130_fd_sc_hd__nand2_1 _24126_ (.A(net4553),
    .B(net4889),
    .Y(_03988_));
 sky130_fd_sc_hd__xnor2_1 _24127_ (.A(_03987_),
    .B(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__xnor2_1 _24128_ (.A(_03986_),
    .B(_03989_),
    .Y(_03990_));
 sky130_fd_sc_hd__nor2_1 _24129_ (.A(net2408),
    .B(_03990_),
    .Y(_03991_));
 sky130_fd_sc_hd__nand2_1 _24130_ (.A(net2408),
    .B(_03990_),
    .Y(_03992_));
 sky130_fd_sc_hd__or2b_1 _24131_ (.A(_03991_),
    .B_N(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__xnor2_2 _24132_ (.A(_03983_),
    .B(_03993_),
    .Y(_03994_));
 sky130_fd_sc_hd__o21a_1 _24133_ (.A1(_03878_),
    .A2(_03883_),
    .B1(_03876_),
    .X(_03995_));
 sky130_fd_sc_hd__a21o_1 _24134_ (.A1(_03878_),
    .A2(_03883_),
    .B1(_03995_),
    .X(_03996_));
 sky130_fd_sc_hd__a21bo_1 _24135_ (.A1(_03897_),
    .A2(_03906_),
    .B1_N(_03907_),
    .X(_03997_));
 sky130_fd_sc_hd__nor2_1 _24136_ (.A(_03996_),
    .B(_03997_),
    .Y(_03998_));
 sky130_fd_sc_hd__nand2_1 _24137_ (.A(_03996_),
    .B(_03997_),
    .Y(_03999_));
 sky130_fd_sc_hd__and2b_1 _24138_ (.A_N(_03998_),
    .B(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__xnor2_2 _24139_ (.A(_03994_),
    .B(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__xnor2_1 _24140_ (.A(_03978_),
    .B(_04001_),
    .Y(_04002_));
 sky130_fd_sc_hd__xnor2_2 _24141_ (.A(_03976_),
    .B(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__o21a_1 _24142_ (.A1(_03892_),
    .A2(_03918_),
    .B1(_03890_),
    .X(_04004_));
 sky130_fd_sc_hd__a21oi_1 _24143_ (.A1(_03892_),
    .A2(_03918_),
    .B1(_04004_),
    .Y(_04005_));
 sky130_fd_sc_hd__o21a_1 _24144_ (.A1(_03909_),
    .A2(_03916_),
    .B1(_03914_),
    .X(_04006_));
 sky130_fd_sc_hd__inv_2 _24145_ (.A(net4651),
    .Y(_04007_));
 sky130_fd_sc_hd__a32o_1 _24146_ (.A1(net4605),
    .A2(net4625),
    .A3(net3052),
    .B1(net4788),
    .B2(_04007_),
    .X(_04008_));
 sky130_fd_sc_hd__nand2_1 _24147_ (.A(net4788),
    .B(net3052),
    .Y(_04009_));
 sky130_fd_sc_hd__or4bb_1 _24148_ (.A(net4651),
    .B(_04009_),
    .C_N(net4605),
    .D_N(net4625),
    .X(_04010_));
 sky130_fd_sc_hd__o21a_1 _24149_ (.A1(_03903_),
    .A2(_04008_),
    .B1(net2023),
    .X(_04011_));
 sky130_fd_sc_hd__or3b_1 _24150_ (.A(net4675),
    .B(net3043),
    .C_N(_03924_),
    .X(_04012_));
 sky130_fd_sc_hd__xor2_1 _24151_ (.A(net1658),
    .B(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__xnor2_2 _24152_ (.A(net1015),
    .B(_04013_),
    .Y(_04014_));
 sky130_fd_sc_hd__xnor2_1 _24153_ (.A(_04005_),
    .B(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__xnor2_1 _24154_ (.A(_04003_),
    .B(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__nor2_1 _24155_ (.A(_03922_),
    .B(_03931_),
    .Y(_04017_));
 sky130_fd_sc_hd__o21ai_1 _24156_ (.A1(_03920_),
    .A2(_04017_),
    .B1(_03932_),
    .Y(_04018_));
 sky130_fd_sc_hd__o21a_1 _24157_ (.A1(net1160),
    .A2(_03927_),
    .B1(_03928_),
    .X(_04019_));
 sky130_fd_sc_hd__a21oi_1 _24158_ (.A1(net1160),
    .A2(_03927_),
    .B1(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__xnor2_1 _24159_ (.A(net739),
    .B(net930),
    .Y(_04021_));
 sky130_fd_sc_hd__xnor2_2 _24160_ (.A(net694),
    .B(_04021_),
    .Y(_04022_));
 sky130_fd_sc_hd__nor2_1 _24161_ (.A(_03869_),
    .B(_03937_),
    .Y(_04023_));
 sky130_fd_sc_hd__nand2_1 _24162_ (.A(_03869_),
    .B(_03937_),
    .Y(_04024_));
 sky130_fd_sc_hd__o21ai_1 _24163_ (.A1(_03935_),
    .A2(_04023_),
    .B1(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__xnor2_1 _24164_ (.A(_04022_),
    .B(net590),
    .Y(_04026_));
 sky130_fd_sc_hd__xnor2_1 _24165_ (.A(_03961_),
    .B(_04026_),
    .Y(_04027_));
 sky130_fd_sc_hd__inv_2 _24166_ (.A(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__inv_2 _24167_ (.A(\pid_q.curr_error[7] ),
    .Y(_04029_));
 sky130_fd_sc_hd__o21ba_1 _24168_ (.A1(_04029_),
    .A2(_03948_),
    .B1_N(\pid_q.prev_error[7] ),
    .X(_04030_));
 sky130_fd_sc_hd__a21o_1 _24169_ (.A1(_04029_),
    .A2(_03948_),
    .B1(_04030_),
    .X(_04031_));
 sky130_fd_sc_hd__xnor2_1 _24170_ (.A(\pid_q.prev_error[8] ),
    .B(\pid_q.curr_error[8] ),
    .Y(_04032_));
 sky130_fd_sc_hd__nand2_1 _24171_ (.A(_04031_),
    .B(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__or2_1 _24172_ (.A(_04031_),
    .B(_04032_),
    .X(_04034_));
 sky130_fd_sc_hd__and3_1 _24173_ (.A(net7511),
    .B(_04033_),
    .C(_04034_),
    .X(_04035_));
 sky130_fd_sc_hd__a221o_1 _24174_ (.A1(net7525),
    .A2(_03959_),
    .B1(net241),
    .B2(net7467),
    .C1(net636),
    .X(_04036_));
 sky130_fd_sc_hd__a22o_1 _24175_ (.A1(\pid_q.curr_int[8] ),
    .A2(net3757),
    .B1(_02870_),
    .B2(_04036_),
    .X(_00673_));
 sky130_fd_sc_hd__inv_2 _24176_ (.A(\pid_q.prev_int[8] ),
    .Y(_04037_));
 sky130_fd_sc_hd__inv_2 _24177_ (.A(\pid_q.curr_int[8] ),
    .Y(_04038_));
 sky130_fd_sc_hd__o21a_1 _24178_ (.A1(_04037_),
    .A2(_03957_),
    .B1(_04038_),
    .X(_04039_));
 sky130_fd_sc_hd__a21o_1 _24179_ (.A1(_04037_),
    .A2(_03957_),
    .B1(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__xor2_1 _24180_ (.A(\pid_q.curr_int[9] ),
    .B(\pid_q.prev_int[9] ),
    .X(_04041_));
 sky130_fd_sc_hd__xnor2_1 _24181_ (.A(_04040_),
    .B(_04041_),
    .Y(_04042_));
 sky130_fd_sc_hd__nand2_1 _24182_ (.A(_04022_),
    .B(net590),
    .Y(_04043_));
 sky130_fd_sc_hd__nor2_1 _24183_ (.A(_04022_),
    .B(net590),
    .Y(_04044_));
 sky130_fd_sc_hd__a31o_1 _24184_ (.A1(_03941_),
    .A2(_03960_),
    .A3(_04043_),
    .B1(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__inv_2 _24185_ (.A(net930),
    .Y(_04046_));
 sky130_fd_sc_hd__a21bo_1 _24186_ (.A1(net739),
    .A2(_04046_),
    .B1_N(net694),
    .X(_04047_));
 sky130_fd_sc_hd__o21ai_1 _24187_ (.A1(net739),
    .A2(_04046_),
    .B1(_04047_),
    .Y(_04048_));
 sky130_fd_sc_hd__a21o_1 _24188_ (.A1(_04003_),
    .A2(_04014_),
    .B1(_04005_),
    .X(_04049_));
 sky130_fd_sc_hd__o21ai_1 _24189_ (.A1(_04003_),
    .A2(_04014_),
    .B1(_04049_),
    .Y(_04050_));
 sky130_fd_sc_hd__inv_2 _24190_ (.A(_03976_),
    .Y(_04051_));
 sky130_fd_sc_hd__o21a_1 _24191_ (.A1(_04051_),
    .A2(_04001_),
    .B1(_03978_),
    .X(_04052_));
 sky130_fd_sc_hd__a21o_1 _24192_ (.A1(_04051_),
    .A2(_04001_),
    .B1(_04052_),
    .X(_04053_));
 sky130_fd_sc_hd__nand2_1 _24193_ (.A(net4590),
    .B(net4836),
    .Y(_04054_));
 sky130_fd_sc_hd__nand2_1 _24194_ (.A(net4580),
    .B(net4853),
    .Y(_04055_));
 sky130_fd_sc_hd__xor2_2 _24195_ (.A(_04054_),
    .B(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__nand2_1 _24196_ (.A(net4603),
    .B(net4803),
    .Y(_04057_));
 sky130_fd_sc_hd__xor2_2 _24197_ (.A(_04056_),
    .B(_04057_),
    .X(_04058_));
 sky130_fd_sc_hd__o21ai_1 _24198_ (.A1(_03986_),
    .A2(_03988_),
    .B1(_03987_),
    .Y(_04059_));
 sky130_fd_sc_hd__a21bo_1 _24199_ (.A1(_03986_),
    .A2(_03988_),
    .B1_N(_04059_),
    .X(_04060_));
 sky130_fd_sc_hd__nand2_1 _24200_ (.A(net4553),
    .B(net4867),
    .Y(_04061_));
 sky130_fd_sc_hd__nand2_1 _24201_ (.A(net4520),
    .B(net4928),
    .Y(_04062_));
 sky130_fd_sc_hd__nand2_1 _24202_ (.A(net4535),
    .B(net4890),
    .Y(_04063_));
 sky130_fd_sc_hd__xnor2_1 _24203_ (.A(_04062_),
    .B(_04063_),
    .Y(_04064_));
 sky130_fd_sc_hd__xnor2_1 _24204_ (.A(_04061_),
    .B(_04064_),
    .Y(_04065_));
 sky130_fd_sc_hd__xnor2_1 _24205_ (.A(_04060_),
    .B(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__xnor2_2 _24206_ (.A(_04058_),
    .B(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__a21bo_1 _24207_ (.A1(net3040),
    .A2(_03973_),
    .B1_N(_03968_),
    .X(_04068_));
 sky130_fd_sc_hd__o21ai_1 _24208_ (.A1(net3040),
    .A2(_03973_),
    .B1(_04068_),
    .Y(_04069_));
 sky130_fd_sc_hd__a21oi_1 _24209_ (.A1(_03983_),
    .A2(_03992_),
    .B1(_03991_),
    .Y(_04070_));
 sky130_fd_sc_hd__and2_1 _24210_ (.A(_04069_),
    .B(_04070_),
    .X(_04071_));
 sky130_fd_sc_hd__or2_1 _24211_ (.A(_04069_),
    .B(_04070_),
    .X(_04072_));
 sky130_fd_sc_hd__or2b_1 _24212_ (.A(net1380),
    .B_N(net1379),
    .X(_04073_));
 sky130_fd_sc_hd__xnor2_2 _24213_ (.A(_04067_),
    .B(_04073_),
    .Y(_04074_));
 sky130_fd_sc_hd__inv_2 _24214_ (.A(_03975_),
    .Y(_04075_));
 sky130_fd_sc_hd__nand2_1 _24215_ (.A(net3743),
    .B(_03887_),
    .Y(_04076_));
 sky130_fd_sc_hd__o21ai_1 _24216_ (.A1(net2410),
    .A2(_04075_),
    .B1(net2021),
    .Y(_04077_));
 sky130_fd_sc_hd__xor2_1 _24217_ (.A(net4993),
    .B(net4959),
    .X(_04078_));
 sky130_fd_sc_hd__nand2_1 _24218_ (.A(net4484),
    .B(_04078_),
    .Y(_04079_));
 sky130_fd_sc_hd__nand2_1 _24219_ (.A(net4937),
    .B(net4501),
    .Y(_04080_));
 sky130_fd_sc_hd__xor2_2 _24220_ (.A(_04079_),
    .B(_04080_),
    .X(_04081_));
 sky130_fd_sc_hd__o21a_1 _24221_ (.A1(_03964_),
    .A2(_03966_),
    .B1(_03965_),
    .X(_04082_));
 sky130_fd_sc_hd__a21oi_2 _24222_ (.A1(_03964_),
    .A2(_03966_),
    .B1(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__xnor2_1 _24223_ (.A(net3040),
    .B(_04083_),
    .Y(_04084_));
 sky130_fd_sc_hd__xnor2_1 _24224_ (.A(_04081_),
    .B(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__xnor2_2 _24225_ (.A(net2024),
    .B(net1657),
    .Y(_04086_));
 sky130_fd_sc_hd__xnor2_1 _24226_ (.A(net1159),
    .B(_04086_),
    .Y(_04087_));
 sky130_fd_sc_hd__xnor2_1 _24227_ (.A(_04074_),
    .B(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__o21ai_1 _24228_ (.A1(_03994_),
    .A2(_03998_),
    .B1(_03999_),
    .Y(_04089_));
 sky130_fd_sc_hd__and3_1 _24229_ (.A(net4590),
    .B(net4604),
    .C(net3053),
    .X(_04090_));
 sky130_fd_sc_hd__xnor2_1 _24230_ (.A(net4789),
    .B(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__a21oi_1 _24231_ (.A1(net4802),
    .A2(_03981_),
    .B1(_04090_),
    .Y(_04092_));
 sky130_fd_sc_hd__mux2_1 _24232_ (.A0(_04091_),
    .A1(_04092_),
    .S(net4624),
    .X(_04093_));
 sky130_fd_sc_hd__xnor2_1 _24233_ (.A(net2022),
    .B(net1656),
    .Y(_04094_));
 sky130_fd_sc_hd__xnor2_2 _24234_ (.A(net1013),
    .B(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__xnor2_1 _24235_ (.A(_04088_),
    .B(_04095_),
    .Y(_04096_));
 sky130_fd_sc_hd__xnor2_1 _24236_ (.A(net793),
    .B(_04096_),
    .Y(_04097_));
 sky130_fd_sc_hd__nor2_1 _24237_ (.A(net1015),
    .B(net1658),
    .Y(_04098_));
 sky130_fd_sc_hd__nand2_1 _24238_ (.A(net1015),
    .B(net1658),
    .Y(_04099_));
 sky130_fd_sc_hd__o21a_1 _24239_ (.A1(_04012_),
    .A2(_04098_),
    .B1(_04099_),
    .X(_04100_));
 sky130_fd_sc_hd__and2_1 _24240_ (.A(_04097_),
    .B(net852),
    .X(_04101_));
 sky130_fd_sc_hd__or2_1 _24241_ (.A(_04097_),
    .B(net852),
    .X(_04102_));
 sky130_fd_sc_hd__and2b_1 _24242_ (.A_N(_04101_),
    .B(_04102_),
    .X(_04103_));
 sky130_fd_sc_hd__xnor2_1 _24243_ (.A(net692),
    .B(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hd__nor2_1 _24244_ (.A(_04048_),
    .B(net589),
    .Y(_04105_));
 sky130_fd_sc_hd__and2_1 _24245_ (.A(_04048_),
    .B(net589),
    .X(_04106_));
 sky130_fd_sc_hd__or2_1 _24246_ (.A(_04105_),
    .B(_04106_),
    .X(_04107_));
 sky130_fd_sc_hd__xnor2_1 _24247_ (.A(_04045_),
    .B(_04107_),
    .Y(_04108_));
 sky130_fd_sc_hd__inv_2 _24248_ (.A(\pid_q.curr_error[8] ),
    .Y(_04109_));
 sky130_fd_sc_hd__a21bo_1 _24249_ (.A1(_04109_),
    .A2(_04031_),
    .B1_N(\pid_q.prev_error[8] ),
    .X(_04110_));
 sky130_fd_sc_hd__o21a_1 _24250_ (.A1(_04109_),
    .A2(_04031_),
    .B1(_04110_),
    .X(_04111_));
 sky130_fd_sc_hd__xnor2_1 _24251_ (.A(\pid_q.prev_error[9] ),
    .B(\pid_q.curr_error[9] ),
    .Y(_04112_));
 sky130_fd_sc_hd__nand2_1 _24252_ (.A(_04111_),
    .B(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__or2_1 _24253_ (.A(_04111_),
    .B(_04112_),
    .X(_04114_));
 sky130_fd_sc_hd__and3_1 _24254_ (.A(net7505),
    .B(_04113_),
    .C(_04114_),
    .X(_04115_));
 sky130_fd_sc_hd__a221o_1 _24255_ (.A1(net7523),
    .A2(_04042_),
    .B1(net269),
    .B2(net7467),
    .C1(net536),
    .X(_04116_));
 sky130_fd_sc_hd__a22o_1 _24256_ (.A1(\pid_q.curr_int[9] ),
    .A2(net3758),
    .B1(_02870_),
    .B2(_04116_),
    .X(_00674_));
 sky130_fd_sc_hd__inv_2 _24257_ (.A(\pid_q.curr_int[10] ),
    .Y(_04117_));
 sky130_fd_sc_hd__nor2_1 _24258_ (.A(_04117_),
    .B(_02868_),
    .Y(_04118_));
 sky130_fd_sc_hd__or2_1 _24259_ (.A(_04048_),
    .B(net589),
    .X(_04119_));
 sky130_fd_sc_hd__o21a_1 _24260_ (.A1(net793),
    .A2(_04095_),
    .B1(_04088_),
    .X(_04120_));
 sky130_fd_sc_hd__a21o_1 _24261_ (.A1(net793),
    .A2(_04095_),
    .B1(_04120_),
    .X(_04121_));
 sky130_fd_sc_hd__o21a_1 _24262_ (.A1(net1159),
    .A2(_04086_),
    .B1(_04074_),
    .X(_04122_));
 sky130_fd_sc_hd__a21o_1 _24263_ (.A1(net1159),
    .A2(_04086_),
    .B1(_04122_),
    .X(_04123_));
 sky130_fd_sc_hd__nand2_1 _24264_ (.A(net4580),
    .B(net4836),
    .Y(_04124_));
 sky130_fd_sc_hd__nand2_1 _24265_ (.A(net4554),
    .B(net4853),
    .Y(_04125_));
 sky130_fd_sc_hd__xor2_2 _24266_ (.A(_04124_),
    .B(_04125_),
    .X(_04126_));
 sky130_fd_sc_hd__nand2_1 _24267_ (.A(net4589),
    .B(net4803),
    .Y(_04127_));
 sky130_fd_sc_hd__xor2_2 _24268_ (.A(_04126_),
    .B(_04127_),
    .X(_04128_));
 sky130_fd_sc_hd__o21ai_1 _24269_ (.A1(_04061_),
    .A2(_04063_),
    .B1(_04062_),
    .Y(_04129_));
 sky130_fd_sc_hd__a21bo_1 _24270_ (.A1(_04061_),
    .A2(_04063_),
    .B1_N(_04129_),
    .X(_04130_));
 sky130_fd_sc_hd__nand2_2 _24271_ (.A(net4917),
    .B(net4502),
    .Y(_04131_));
 sky130_fd_sc_hd__nand2_1 _24272_ (.A(net4522),
    .B(net4885),
    .Y(_04132_));
 sky130_fd_sc_hd__nand2_1 _24273_ (.A(net4536),
    .B(net4862),
    .Y(_04133_));
 sky130_fd_sc_hd__xnor2_1 _24274_ (.A(_04132_),
    .B(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hd__xnor2_2 _24275_ (.A(_04131_),
    .B(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__xnor2_1 _24276_ (.A(net2405),
    .B(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__xnor2_2 _24277_ (.A(_04128_),
    .B(_04136_),
    .Y(_04137_));
 sky130_fd_sc_hd__a21o_1 _24278_ (.A1(_04081_),
    .A2(_04083_),
    .B1(net3040),
    .X(_04138_));
 sky130_fd_sc_hd__o21ai_1 _24279_ (.A1(_04081_),
    .A2(_04083_),
    .B1(_04138_),
    .Y(_04139_));
 sky130_fd_sc_hd__o21a_1 _24280_ (.A1(_04060_),
    .A2(_04065_),
    .B1(_04058_),
    .X(_04140_));
 sky130_fd_sc_hd__a21o_1 _24281_ (.A1(_04060_),
    .A2(_04065_),
    .B1(_04140_),
    .X(_04141_));
 sky130_fd_sc_hd__xnor2_1 _24282_ (.A(net1655),
    .B(net1654),
    .Y(_04142_));
 sky130_fd_sc_hd__xnor2_2 _24283_ (.A(_04137_),
    .B(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__a21o_1 _24284_ (.A1(net2020),
    .A2(net1657),
    .B1(net2409),
    .X(_04144_));
 sky130_fd_sc_hd__o21a_1 _24285_ (.A1(net4960),
    .A2(_03605_),
    .B1(net4994),
    .X(_04145_));
 sky130_fd_sc_hd__a21o_1 _24286_ (.A1(net4959),
    .A2(_03605_),
    .B1(_04145_),
    .X(_04146_));
 sky130_fd_sc_hd__o31ai_1 _24287_ (.A1(net4993),
    .A2(net4959),
    .A3(net4937),
    .B1(net4484),
    .Y(_04147_));
 sky130_fd_sc_hd__a21o_1 _24288_ (.A1(net4937),
    .A2(_04146_),
    .B1(_04147_),
    .X(_04148_));
 sky130_fd_sc_hd__xnor2_1 _24289_ (.A(net3041),
    .B(_04148_),
    .Y(_04149_));
 sky130_fd_sc_hd__xor2_2 _24290_ (.A(net2024),
    .B(net1653),
    .X(_04150_));
 sky130_fd_sc_hd__xnor2_1 _24291_ (.A(_04144_),
    .B(_04150_),
    .Y(_04151_));
 sky130_fd_sc_hd__xnor2_2 _24292_ (.A(_04143_),
    .B(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__a21oi_2 _24293_ (.A1(_04067_),
    .A2(net1379),
    .B1(net1380),
    .Y(_04153_));
 sky130_fd_sc_hd__and3_1 _24294_ (.A(net4580),
    .B(net4590),
    .C(net3053),
    .X(_04154_));
 sky130_fd_sc_hd__xnor2_1 _24295_ (.A(net3044),
    .B(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__a21o_1 _24296_ (.A1(net4803),
    .A2(_04056_),
    .B1(_04154_),
    .X(_04156_));
 sky130_fd_sc_hd__mux2_1 _24297_ (.A0(_04155_),
    .A1(_04156_),
    .S(net4603),
    .X(_04157_));
 sky130_fd_sc_hd__or3b_1 _24298_ (.A(net4624),
    .B(net3044),
    .C_N(_04090_),
    .X(_04158_));
 sky130_fd_sc_hd__xnor2_1 _24299_ (.A(_04157_),
    .B(_04158_),
    .Y(_04159_));
 sky130_fd_sc_hd__xnor2_2 _24300_ (.A(_04153_),
    .B(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__xnor2_1 _24301_ (.A(_04152_),
    .B(_04160_),
    .Y(_04161_));
 sky130_fd_sc_hd__xnor2_2 _24302_ (.A(_04123_),
    .B(_04161_),
    .Y(_04162_));
 sky130_fd_sc_hd__o21a_1 _24303_ (.A1(net1013),
    .A2(net1656),
    .B1(net2022),
    .X(_04163_));
 sky130_fd_sc_hd__a21o_1 _24304_ (.A1(net1013),
    .A2(net1656),
    .B1(_04163_),
    .X(_04164_));
 sky130_fd_sc_hd__xnor2_1 _24305_ (.A(_04162_),
    .B(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__xnor2_1 _24306_ (.A(_04121_),
    .B(_04165_),
    .Y(_04166_));
 sky130_fd_sc_hd__a21o_1 _24307_ (.A1(net692),
    .A2(_04102_),
    .B1(_04101_),
    .X(_04167_));
 sky130_fd_sc_hd__xnor2_2 _24308_ (.A(net634),
    .B(net633),
    .Y(_04168_));
 sky130_fd_sc_hd__nor3_1 _24309_ (.A(_04045_),
    .B(_04106_),
    .C(_04168_),
    .Y(_04169_));
 sky130_fd_sc_hd__a31o_1 _24310_ (.A1(_04045_),
    .A2(_04119_),
    .A3(_04168_),
    .B1(_04169_),
    .X(_04170_));
 sky130_fd_sc_hd__inv_2 _24311_ (.A(\pid_q.prev_int[9] ),
    .Y(_04171_));
 sky130_fd_sc_hd__inv_2 _24312_ (.A(\pid_q.curr_int[9] ),
    .Y(_04172_));
 sky130_fd_sc_hd__o21a_1 _24313_ (.A1(_04171_),
    .A2(_04040_),
    .B1(_04172_),
    .X(_04173_));
 sky130_fd_sc_hd__a21o_1 _24314_ (.A1(_04171_),
    .A2(_04040_),
    .B1(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__xor2_1 _24315_ (.A(\pid_q.curr_int[10] ),
    .B(\pid_q.prev_int[10] ),
    .X(_04175_));
 sky130_fd_sc_hd__xnor2_1 _24316_ (.A(_04174_),
    .B(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hd__mux2_1 _24317_ (.A0(_04105_),
    .A1(_04106_),
    .S(_04168_),
    .X(_04177_));
 sky130_fd_sc_hd__inv_2 _24318_ (.A(\pid_q.curr_error[9] ),
    .Y(_04178_));
 sky130_fd_sc_hd__o21ba_1 _24319_ (.A1(_04178_),
    .A2(_04111_),
    .B1_N(\pid_q.prev_error[9] ),
    .X(_04179_));
 sky130_fd_sc_hd__a21o_1 _24320_ (.A1(_04178_),
    .A2(_04111_),
    .B1(_04179_),
    .X(_04180_));
 sky130_fd_sc_hd__xnor2_1 _24321_ (.A(\pid_q.prev_error[10] ),
    .B(\pid_q.curr_error[10] ),
    .Y(_04181_));
 sky130_fd_sc_hd__nand2_1 _24322_ (.A(_04180_),
    .B(_04181_),
    .Y(_04182_));
 sky130_fd_sc_hd__or2_1 _24323_ (.A(_04180_),
    .B(_04181_),
    .X(_04183_));
 sky130_fd_sc_hd__and3_1 _24324_ (.A(net7506),
    .B(_04182_),
    .C(_04183_),
    .X(_04184_));
 sky130_fd_sc_hd__a221o_1 _24325_ (.A1(net7524),
    .A2(_04176_),
    .B1(net510),
    .B2(net7464),
    .C1(net460),
    .X(_04185_));
 sky130_fd_sc_hd__a211o_1 _24326_ (.A1(net7464),
    .A2(net238),
    .B1(_04185_),
    .C1(_04118_),
    .X(_04186_));
 sky130_fd_sc_hd__o21a_1 _24327_ (.A1(_02869_),
    .A2(_04118_),
    .B1(_04186_),
    .X(_00675_));
 sky130_fd_sc_hd__inv_2 _24328_ (.A(\pid_q.prev_int[10] ),
    .Y(_04187_));
 sky130_fd_sc_hd__o21a_1 _24329_ (.A1(_04187_),
    .A2(_04174_),
    .B1(net3736),
    .X(_04188_));
 sky130_fd_sc_hd__a21oi_2 _24330_ (.A1(_04187_),
    .A2(_04174_),
    .B1(_04188_),
    .Y(_04189_));
 sky130_fd_sc_hd__xnor2_1 _24331_ (.A(net5177),
    .B(\pid_q.prev_int[11] ),
    .Y(_04190_));
 sky130_fd_sc_hd__xnor2_1 _24332_ (.A(_04189_),
    .B(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__nor2_1 _24333_ (.A(_04026_),
    .B(_04107_),
    .Y(_04192_));
 sky130_fd_sc_hd__nor2_1 _24334_ (.A(_03944_),
    .B(_04168_),
    .Y(_04193_));
 sky130_fd_sc_hd__a211oi_1 _24335_ (.A1(_03942_),
    .A2(_04043_),
    .B1(_04106_),
    .C1(_04044_),
    .Y(_04194_));
 sky130_fd_sc_hd__a211o_1 _24336_ (.A1(net634),
    .A2(net633),
    .B1(_04194_),
    .C1(_04105_),
    .X(_04195_));
 sky130_fd_sc_hd__o21ai_1 _24337_ (.A1(net634),
    .A2(net633),
    .B1(_04195_),
    .Y(_04196_));
 sky130_fd_sc_hd__a31o_1 _24338_ (.A1(net376),
    .A2(_04192_),
    .A3(_04193_),
    .B1(_04196_),
    .X(_04197_));
 sky130_fd_sc_hd__o21ba_1 _24339_ (.A1(_04144_),
    .A2(_04150_),
    .B1_N(_04143_),
    .X(_04198_));
 sky130_fd_sc_hd__a21oi_1 _24340_ (.A1(_04144_),
    .A2(_04150_),
    .B1(_04198_),
    .Y(_04199_));
 sky130_fd_sc_hd__nand2_1 _24341_ (.A(net4917),
    .B(net4485),
    .Y(_04200_));
 sky130_fd_sc_hd__nand2_1 _24342_ (.A(net4522),
    .B(net4873),
    .Y(_04201_));
 sky130_fd_sc_hd__nand2_1 _24343_ (.A(net4895),
    .B(net4504),
    .Y(_04202_));
 sky130_fd_sc_hd__xnor2_1 _24344_ (.A(_04201_),
    .B(_04202_),
    .Y(_04203_));
 sky130_fd_sc_hd__xnor2_2 _24345_ (.A(_04200_),
    .B(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__o21ai_1 _24346_ (.A1(_04131_),
    .A2(_04133_),
    .B1(_04132_),
    .Y(_04205_));
 sky130_fd_sc_hd__a21bo_1 _24347_ (.A1(_04131_),
    .A2(_04133_),
    .B1_N(_04205_),
    .X(_04206_));
 sky130_fd_sc_hd__nand2_1 _24348_ (.A(net4536),
    .B(net4857),
    .Y(_04207_));
 sky130_fd_sc_hd__nand2_1 _24349_ (.A(net4555),
    .B(net4837),
    .Y(_04208_));
 sky130_fd_sc_hd__xor2_2 _24350_ (.A(_04207_),
    .B(_04208_),
    .X(_04209_));
 sky130_fd_sc_hd__nand2_1 _24351_ (.A(net4581),
    .B(net4805),
    .Y(_04210_));
 sky130_fd_sc_hd__xor2_2 _24352_ (.A(_04209_),
    .B(_04210_),
    .X(_04211_));
 sky130_fd_sc_hd__xor2_1 _24353_ (.A(_04206_),
    .B(_04211_),
    .X(_04212_));
 sky130_fd_sc_hd__xnor2_2 _24354_ (.A(_04204_),
    .B(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__o21a_1 _24355_ (.A1(net4960),
    .A2(net4937),
    .B1(net3041),
    .X(_04214_));
 sky130_fd_sc_hd__a31oi_1 _24356_ (.A1(net4937),
    .A2(_03605_),
    .A3(_04078_),
    .B1(net3742),
    .Y(_04215_));
 sky130_fd_sc_hd__a21o_1 _24357_ (.A1(net4960),
    .A2(net4937),
    .B1(net3041),
    .X(_04216_));
 sky130_fd_sc_hd__o211a_1 _24358_ (.A1(net4994),
    .A2(_04214_),
    .B1(_04215_),
    .C1(_04216_),
    .X(_04217_));
 sky130_fd_sc_hd__o21a_1 _24359_ (.A1(net2405),
    .A2(_04135_),
    .B1(_04128_),
    .X(_04218_));
 sky130_fd_sc_hd__a21oi_1 _24360_ (.A1(net2405),
    .A2(_04135_),
    .B1(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hd__xnor2_1 _24361_ (.A(net2019),
    .B(net1652),
    .Y(_04220_));
 sky130_fd_sc_hd__xnor2_2 _24362_ (.A(_04213_),
    .B(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__a21o_1 _24363_ (.A1(net2020),
    .A2(net1653),
    .B1(net2409),
    .X(_04222_));
 sky130_fd_sc_hd__a31o_1 _24364_ (.A1(net4993),
    .A2(net4959),
    .A3(net4937),
    .B1(_04147_),
    .X(_04223_));
 sky130_fd_sc_hd__xnor2_1 _24365_ (.A(net3041),
    .B(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__xor2_2 _24366_ (.A(net2024),
    .B(net2404),
    .X(_04225_));
 sky130_fd_sc_hd__xnor2_1 _24367_ (.A(_04222_),
    .B(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__xnor2_2 _24368_ (.A(_04221_),
    .B(_04226_),
    .Y(_04227_));
 sky130_fd_sc_hd__a21o_1 _24369_ (.A1(net1655),
    .A2(net1654),
    .B1(_04137_),
    .X(_04228_));
 sky130_fd_sc_hd__o21a_1 _24370_ (.A1(net1655),
    .A2(net1654),
    .B1(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__and3_1 _24371_ (.A(net4554),
    .B(net4581),
    .C(net3053),
    .X(_04230_));
 sky130_fd_sc_hd__xnor2_1 _24372_ (.A(net4789),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__a21oi_1 _24373_ (.A1(net4804),
    .A2(_04126_),
    .B1(_04230_),
    .Y(_04232_));
 sky130_fd_sc_hd__mux2_1 _24374_ (.A0(_04231_),
    .A1(_04232_),
    .S(net4589),
    .X(_04233_));
 sky130_fd_sc_hd__or3b_1 _24375_ (.A(net4603),
    .B(net3044),
    .C_N(_04154_),
    .X(_04234_));
 sky130_fd_sc_hd__xor2_1 _24376_ (.A(_04233_),
    .B(_04234_),
    .X(_04235_));
 sky130_fd_sc_hd__xnor2_1 _24377_ (.A(_04229_),
    .B(_04235_),
    .Y(_04236_));
 sky130_fd_sc_hd__xnor2_1 _24378_ (.A(_04227_),
    .B(net1012),
    .Y(_04237_));
 sky130_fd_sc_hd__xnor2_1 _24379_ (.A(_04199_),
    .B(_04237_),
    .Y(_04238_));
 sky130_fd_sc_hd__a21o_1 _24380_ (.A1(_04152_),
    .A2(_04160_),
    .B1(_04123_),
    .X(_04239_));
 sky130_fd_sc_hd__o21ai_1 _24381_ (.A1(_04152_),
    .A2(_04160_),
    .B1(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__a21bo_1 _24382_ (.A1(_04153_),
    .A2(_04157_),
    .B1_N(_04158_),
    .X(_04241_));
 sky130_fd_sc_hd__o21a_1 _24383_ (.A1(_04153_),
    .A2(_04157_),
    .B1(_04241_),
    .X(_04242_));
 sky130_fd_sc_hd__nor2_1 _24384_ (.A(_04240_),
    .B(net929),
    .Y(_04243_));
 sky130_fd_sc_hd__nand2_1 _24385_ (.A(_04240_),
    .B(net929),
    .Y(_04244_));
 sky130_fd_sc_hd__or2b_1 _24386_ (.A(_04243_),
    .B_N(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__xnor2_1 _24387_ (.A(_04238_),
    .B(_04245_),
    .Y(_04246_));
 sky130_fd_sc_hd__o21a_1 _24388_ (.A1(_04162_),
    .A2(_04164_),
    .B1(_04121_),
    .X(_04247_));
 sky130_fd_sc_hd__a21o_1 _24389_ (.A1(_04162_),
    .A2(_04164_),
    .B1(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__xnor2_1 _24390_ (.A(net588),
    .B(net587),
    .Y(_04249_));
 sky130_fd_sc_hd__xnor2_1 _24391_ (.A(_04197_),
    .B(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__inv_2 _24392_ (.A(\pid_q.curr_error[10] ),
    .Y(_04251_));
 sky130_fd_sc_hd__o21ba_1 _24393_ (.A1(_04251_),
    .A2(_04180_),
    .B1_N(\pid_q.prev_error[10] ),
    .X(_04252_));
 sky130_fd_sc_hd__a21o_1 _24394_ (.A1(_04251_),
    .A2(_04180_),
    .B1(_04252_),
    .X(_04253_));
 sky130_fd_sc_hd__xnor2_1 _24395_ (.A(\pid_q.prev_error[11] ),
    .B(\pid_q.curr_error[11] ),
    .Y(_04254_));
 sky130_fd_sc_hd__nand2_1 _24396_ (.A(_04253_),
    .B(_04254_),
    .Y(_04255_));
 sky130_fd_sc_hd__or2_1 _24397_ (.A(_04253_),
    .B(_04254_),
    .X(_04256_));
 sky130_fd_sc_hd__and3_1 _24398_ (.A(net7506),
    .B(_04255_),
    .C(_04256_),
    .X(_04257_));
 sky130_fd_sc_hd__a221o_1 _24399_ (.A1(net7522),
    .A2(_04191_),
    .B1(net292),
    .B2(net7465),
    .C1(net374),
    .X(_04258_));
 sky130_fd_sc_hd__a22o_1 _24400_ (.A1(net9077),
    .A2(net3757),
    .B1(net2433),
    .B2(_04258_),
    .X(_00676_));
 sky130_fd_sc_hd__a21o_1 _24401_ (.A1(\pid_q.prev_int[11] ),
    .A2(_04189_),
    .B1(net5177),
    .X(_04259_));
 sky130_fd_sc_hd__or2_1 _24402_ (.A(\pid_q.prev_int[11] ),
    .B(_04189_),
    .X(_04260_));
 sky130_fd_sc_hd__nand2_1 _24403_ (.A(_04259_),
    .B(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__xor2_1 _24404_ (.A(net5175),
    .B(\pid_q.prev_int[12] ),
    .X(_04262_));
 sky130_fd_sc_hd__xnor2_1 _24405_ (.A(_04261_),
    .B(_04262_),
    .Y(_04263_));
 sky130_fd_sc_hd__nand2_1 _24406_ (.A(net588),
    .B(net587),
    .Y(_04264_));
 sky130_fd_sc_hd__nor2_1 _24407_ (.A(net588),
    .B(net587),
    .Y(_04265_));
 sky130_fd_sc_hd__a311o_1 _24408_ (.A1(net376),
    .A2(_04192_),
    .A3(_04193_),
    .B1(_04265_),
    .C1(_04196_),
    .X(_04266_));
 sky130_fd_sc_hd__nand2_1 _24409_ (.A(_04264_),
    .B(_04266_),
    .Y(_04267_));
 sky130_fd_sc_hd__a21oi_2 _24410_ (.A1(_04238_),
    .A2(_04244_),
    .B1(_04243_),
    .Y(_04268_));
 sky130_fd_sc_hd__a21o_1 _24411_ (.A1(_04222_),
    .A2(_04225_),
    .B1(_04221_),
    .X(_04269_));
 sky130_fd_sc_hd__o21a_1 _24412_ (.A1(_04222_),
    .A2(_04225_),
    .B1(_04269_),
    .X(_04270_));
 sky130_fd_sc_hd__o21a_1 _24413_ (.A1(net2019),
    .A2(net1652),
    .B1(_04213_),
    .X(_04271_));
 sky130_fd_sc_hd__a21oi_2 _24414_ (.A1(net2019),
    .A2(net1652),
    .B1(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__and3_1 _24415_ (.A(net4537),
    .B(net4555),
    .C(net3054),
    .X(_04273_));
 sky130_fd_sc_hd__xnor2_1 _24416_ (.A(net4791),
    .B(_04273_),
    .Y(_04274_));
 sky130_fd_sc_hd__a21oi_1 _24417_ (.A1(net4798),
    .A2(_04209_),
    .B1(_04273_),
    .Y(_04275_));
 sky130_fd_sc_hd__mux2_1 _24418_ (.A0(_04274_),
    .A1(_04275_),
    .S(net4581),
    .X(_04276_));
 sky130_fd_sc_hd__and3b_1 _24419_ (.A_N(net4589),
    .B(net4791),
    .C(_04230_),
    .X(_04277_));
 sky130_fd_sc_hd__xnor2_1 _24420_ (.A(_04276_),
    .B(_04277_),
    .Y(_04278_));
 sky130_fd_sc_hd__xnor2_2 _24421_ (.A(_04272_),
    .B(_04278_),
    .Y(_04279_));
 sky130_fd_sc_hd__nand2_1 _24422_ (.A(net2409),
    .B(net2404),
    .Y(_04280_));
 sky130_fd_sc_hd__o21ai_1 _24423_ (.A1(net2020),
    .A2(net2404),
    .B1(_04280_),
    .Y(_04281_));
 sky130_fd_sc_hd__a21o_1 _24424_ (.A1(net4994),
    .A2(_04216_),
    .B1(_04214_),
    .X(_04282_));
 sky130_fd_sc_hd__nand2_1 _24425_ (.A(net4485),
    .B(_04282_),
    .Y(_04283_));
 sky130_fd_sc_hd__xor2_4 _24426_ (.A(net1651),
    .B(net1650),
    .X(_04284_));
 sky130_fd_sc_hd__o21a_1 _24427_ (.A1(_04206_),
    .A2(_04211_),
    .B1(_04204_),
    .X(_04285_));
 sky130_fd_sc_hd__a21o_1 _24428_ (.A1(_04206_),
    .A2(_04211_),
    .B1(_04285_),
    .X(_04286_));
 sky130_fd_sc_hd__nand2_1 _24429_ (.A(net4872),
    .B(net4504),
    .Y(_04287_));
 sky130_fd_sc_hd__or3_1 _24430_ (.A(net4895),
    .B(net4504),
    .C(_04200_),
    .X(_04288_));
 sky130_fd_sc_hd__o21a_1 _24431_ (.A1(net4490),
    .A2(_04287_),
    .B1(_04288_),
    .X(_04289_));
 sky130_fd_sc_hd__inv_2 _24432_ (.A(net4872),
    .Y(_04290_));
 sky130_fd_sc_hd__nand2_1 _24433_ (.A(net4896),
    .B(net3745),
    .Y(_04291_));
 sky130_fd_sc_hd__a21o_1 _24434_ (.A1(net4872),
    .A2(net3745),
    .B1(net3753),
    .X(_04292_));
 sky130_fd_sc_hd__a22o_1 _24435_ (.A1(net3753),
    .A2(_04287_),
    .B1(_04292_),
    .B2(net4515),
    .X(_04293_));
 sky130_fd_sc_hd__a32o_1 _24436_ (.A1(net4918),
    .A2(_04290_),
    .A3(_04291_),
    .B1(_04293_),
    .B2(net4896),
    .X(_04294_));
 sky130_fd_sc_hd__nand2_1 _24437_ (.A(net4493),
    .B(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__inv_2 _24438_ (.A(net4515),
    .Y(_04296_));
 sky130_fd_sc_hd__a211o_1 _24439_ (.A1(_04296_),
    .A2(net4918),
    .B1(net4896),
    .C1(_04287_),
    .X(_04297_));
 sky130_fd_sc_hd__o211a_1 _24440_ (.A1(net4515),
    .A2(_04289_),
    .B1(_04295_),
    .C1(_04297_),
    .X(_04298_));
 sky130_fd_sc_hd__nand2_1 _24441_ (.A(net4544),
    .B(net4824),
    .Y(_04299_));
 sky130_fd_sc_hd__nand2_1 _24442_ (.A(net4516),
    .B(net4844),
    .Y(_04300_));
 sky130_fd_sc_hd__xor2_1 _24443_ (.A(_04299_),
    .B(_04300_),
    .X(_04301_));
 sky130_fd_sc_hd__and3_1 _24444_ (.A(net4565),
    .B(net4808),
    .C(_04301_),
    .X(_04302_));
 sky130_fd_sc_hd__a21oi_1 _24445_ (.A1(net4555),
    .A2(net4808),
    .B1(_04301_),
    .Y(_04303_));
 sky130_fd_sc_hd__or2_1 _24446_ (.A(_04302_),
    .B(_04303_),
    .X(_04304_));
 sky130_fd_sc_hd__xnor2_2 _24447_ (.A(_04298_),
    .B(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__xor2_2 _24448_ (.A(_04286_),
    .B(_04305_),
    .X(_04306_));
 sky130_fd_sc_hd__xor2_2 _24449_ (.A(_04284_),
    .B(_04306_),
    .X(_04307_));
 sky130_fd_sc_hd__xnor2_1 _24450_ (.A(_04279_),
    .B(_04307_),
    .Y(_04308_));
 sky130_fd_sc_hd__xnor2_1 _24451_ (.A(_04270_),
    .B(_04308_),
    .Y(_04309_));
 sky130_fd_sc_hd__o21a_1 _24452_ (.A1(_04229_),
    .A2(_04233_),
    .B1(_04234_),
    .X(_04310_));
 sky130_fd_sc_hd__a21o_1 _24453_ (.A1(_04229_),
    .A2(_04233_),
    .B1(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__o21ba_1 _24454_ (.A1(_04227_),
    .A2(net1012),
    .B1_N(_04199_),
    .X(_04312_));
 sky130_fd_sc_hd__a21o_1 _24455_ (.A1(_04227_),
    .A2(net1012),
    .B1(_04312_),
    .X(_04313_));
 sky130_fd_sc_hd__nand2b_2 _24456_ (.A_N(net928),
    .B(_04313_),
    .Y(_04314_));
 sky130_fd_sc_hd__or2b_2 _24457_ (.A(_04313_),
    .B_N(net928),
    .X(_04315_));
 sky130_fd_sc_hd__nand2_1 _24458_ (.A(_04314_),
    .B(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__xnor2_1 _24459_ (.A(net792),
    .B(_04316_),
    .Y(_04317_));
 sky130_fd_sc_hd__xnor2_1 _24460_ (.A(_04268_),
    .B(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hd__xnor2_1 _24461_ (.A(_04267_),
    .B(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__inv_2 _24462_ (.A(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__nand2_1 _24463_ (.A(\pid_q.prev_error[12] ),
    .B(net5167),
    .Y(_04321_));
 sky130_fd_sc_hd__or2_1 _24464_ (.A(\pid_q.prev_error[12] ),
    .B(net5167),
    .X(_04322_));
 sky130_fd_sc_hd__nand2_1 _24465_ (.A(_04321_),
    .B(_04322_),
    .Y(_04323_));
 sky130_fd_sc_hd__o21ba_1 _24466_ (.A1(\pid_q.prev_error[11] ),
    .A2(\pid_q.curr_error[11] ),
    .B1_N(_04253_),
    .X(_04324_));
 sky130_fd_sc_hd__a21oi_1 _24467_ (.A1(\pid_q.prev_error[11] ),
    .A2(\pid_q.curr_error[11] ),
    .B1(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__xnor2_1 _24468_ (.A(_04323_),
    .B(_04325_),
    .Y(_04326_));
 sky130_fd_sc_hd__nor2_1 _24469_ (.A(net4001),
    .B(_04326_),
    .Y(_04327_));
 sky130_fd_sc_hd__a221o_1 _24470_ (.A1(net7522),
    .A2(_04263_),
    .B1(net236),
    .B2(net7465),
    .C1(net290),
    .X(_04328_));
 sky130_fd_sc_hd__a22o_1 _24471_ (.A1(net5175),
    .A2(net3757),
    .B1(net2433),
    .B2(_04328_),
    .X(_00677_));
 sky130_fd_sc_hd__inv_2 _24472_ (.A(net2433),
    .Y(_04329_));
 sky130_fd_sc_hd__inv_2 _24473_ (.A(net7524),
    .Y(_04330_));
 sky130_fd_sc_hd__nand2_1 _24474_ (.A(net5173),
    .B(\pid_q.prev_int[13] ),
    .Y(_04331_));
 sky130_fd_sc_hd__or2_1 _24475_ (.A(net5173),
    .B(\pid_q.prev_int[13] ),
    .X(_04332_));
 sky130_fd_sc_hd__nand2_1 _24476_ (.A(_04331_),
    .B(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__or2_1 _24477_ (.A(net5175),
    .B(\pid_q.prev_int[12] ),
    .X(_04334_));
 sky130_fd_sc_hd__and2_1 _24478_ (.A(net5175),
    .B(\pid_q.prev_int[12] ),
    .X(_04335_));
 sky130_fd_sc_hd__a31oi_2 _24479_ (.A1(_04259_),
    .A2(_04260_),
    .A3(_04334_),
    .B1(_04335_),
    .Y(_04336_));
 sky130_fd_sc_hd__xnor2_1 _24480_ (.A(_04333_),
    .B(_04336_),
    .Y(_04337_));
 sky130_fd_sc_hd__xor2_1 _24481_ (.A(net1650),
    .B(_04306_),
    .X(_04338_));
 sky130_fd_sc_hd__o21ai_2 _24482_ (.A1(net1651),
    .A2(_04338_),
    .B1(net2018),
    .Y(_04339_));
 sky130_fd_sc_hd__o21ai_1 _24483_ (.A1(net4485),
    .A2(_04202_),
    .B1(_04288_),
    .Y(_04340_));
 sky130_fd_sc_hd__a2bb2o_1 _24484_ (.A1_N(_04200_),
    .A2_N(_04202_),
    .B1(_04340_),
    .B2(net4515),
    .X(_04341_));
 sky130_fd_sc_hd__a2bb2o_2 _24485_ (.A1_N(_04298_),
    .A2_N(_04304_),
    .B1(_04341_),
    .B2(net4873),
    .X(_04342_));
 sky130_fd_sc_hd__nand2_2 _24486_ (.A(net4523),
    .B(net4825),
    .Y(_04343_));
 sky130_fd_sc_hd__nand2_1 _24487_ (.A(net4545),
    .B(net4809),
    .Y(_04344_));
 sky130_fd_sc_hd__nand2_1 _24488_ (.A(net4848),
    .B(net4505),
    .Y(_04345_));
 sky130_fd_sc_hd__xor2_1 _24489_ (.A(_04344_),
    .B(_04345_),
    .X(_04346_));
 sky130_fd_sc_hd__xnor2_2 _24490_ (.A(_04343_),
    .B(_04346_),
    .Y(_04347_));
 sky130_fd_sc_hd__a21o_1 _24491_ (.A1(_03197_),
    .A2(net4499),
    .B1(net3756),
    .X(_04348_));
 sky130_fd_sc_hd__nand2_1 _24492_ (.A(_04291_),
    .B(net3037),
    .Y(_04349_));
 sky130_fd_sc_hd__or2_1 _24493_ (.A(net4894),
    .B(net4871),
    .X(_04350_));
 sky130_fd_sc_hd__o21ai_1 _24494_ (.A1(net4919),
    .A2(_04350_),
    .B1(net4491),
    .Y(_04351_));
 sky130_fd_sc_hd__a21o_1 _24495_ (.A1(net4871),
    .A2(_04349_),
    .B1(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__xnor2_2 _24496_ (.A(_04347_),
    .B(_04352_),
    .Y(_04353_));
 sky130_fd_sc_hd__xnor2_2 _24497_ (.A(_04342_),
    .B(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__xnor2_2 _24498_ (.A(_04284_),
    .B(_04354_),
    .Y(_04355_));
 sky130_fd_sc_hd__o21a_1 _24499_ (.A1(_04286_),
    .A2(_04305_),
    .B1(net1650),
    .X(_04356_));
 sky130_fd_sc_hd__a21o_1 _24500_ (.A1(_04286_),
    .A2(_04305_),
    .B1(_04356_),
    .X(_04357_));
 sky130_fd_sc_hd__inv_2 _24501_ (.A(net4555),
    .Y(_04358_));
 sky130_fd_sc_hd__a32o_1 _24502_ (.A1(net4516),
    .A2(net4537),
    .A3(net3054),
    .B1(net4793),
    .B2(_04358_),
    .X(_04359_));
 sky130_fd_sc_hd__or4b_1 _24503_ (.A(_04296_),
    .B(net4551),
    .C(net2406),
    .D_N(net4539),
    .X(_04360_));
 sky130_fd_sc_hd__o21ai_2 _24504_ (.A1(_04302_),
    .A2(_04359_),
    .B1(net2017),
    .Y(_04361_));
 sky130_fd_sc_hd__or3b_1 _24505_ (.A(net4582),
    .B(net3045),
    .C_N(_04273_),
    .X(_04362_));
 sky130_fd_sc_hd__xor2_1 _24506_ (.A(_04361_),
    .B(_04362_),
    .X(_04363_));
 sky130_fd_sc_hd__xnor2_2 _24507_ (.A(_04357_),
    .B(_04363_),
    .Y(_04364_));
 sky130_fd_sc_hd__xor2_1 _24508_ (.A(_04355_),
    .B(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__xnor2_2 _24509_ (.A(_04339_),
    .B(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__o21ba_1 _24510_ (.A1(_04272_),
    .A2(_04276_),
    .B1_N(_04277_),
    .X(_04367_));
 sky130_fd_sc_hd__a21oi_2 _24511_ (.A1(_04272_),
    .A2(_04276_),
    .B1(_04367_),
    .Y(_04368_));
 sky130_fd_sc_hd__o21a_1 _24512_ (.A1(_04279_),
    .A2(_04307_),
    .B1(_04270_),
    .X(_04369_));
 sky130_fd_sc_hd__a21o_1 _24513_ (.A1(_04279_),
    .A2(_04307_),
    .B1(_04369_),
    .X(_04370_));
 sky130_fd_sc_hd__xnor2_1 _24514_ (.A(_04368_),
    .B(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__xnor2_2 _24515_ (.A(_04366_),
    .B(_04371_),
    .Y(_04372_));
 sky130_fd_sc_hd__inv_2 _24516_ (.A(_04372_),
    .Y(_04373_));
 sky130_fd_sc_hd__or2_1 _24517_ (.A(_04268_),
    .B(net792),
    .X(_04374_));
 sky130_fd_sc_hd__nand2_1 _24518_ (.A(_04268_),
    .B(net792),
    .Y(_04375_));
 sky130_fd_sc_hd__a21bo_1 _24519_ (.A1(net792),
    .A2(_04315_),
    .B1_N(_04314_),
    .X(_04376_));
 sky130_fd_sc_hd__inv_2 _24520_ (.A(net792),
    .Y(_04377_));
 sky130_fd_sc_hd__o2bb2a_1 _24521_ (.A1_N(_04268_),
    .A2_N(_04376_),
    .B1(_04314_),
    .B2(_04377_),
    .X(_04378_));
 sky130_fd_sc_hd__o22a_1 _24522_ (.A1(net792),
    .A2(_04315_),
    .B1(_04376_),
    .B2(_04268_),
    .X(_04379_));
 sky130_fd_sc_hd__mux2_1 _24523_ (.A0(_04378_),
    .A1(_04379_),
    .S(_04267_),
    .X(_04380_));
 sky130_fd_sc_hd__o221a_1 _24524_ (.A1(_04315_),
    .A2(_04374_),
    .B1(_04375_),
    .B2(_04314_),
    .C1(_04380_),
    .X(_04381_));
 sky130_fd_sc_hd__xnor2_1 _24525_ (.A(_04373_),
    .B(_04381_),
    .Y(_04382_));
 sky130_fd_sc_hd__inv_2 _24526_ (.A(net7463),
    .Y(_04383_));
 sky130_fd_sc_hd__a21bo_1 _24527_ (.A1(_04321_),
    .A2(_04325_),
    .B1_N(_04322_),
    .X(_04384_));
 sky130_fd_sc_hd__xnor2_1 _24528_ (.A(\pid_q.prev_error[13] ),
    .B(net5166),
    .Y(_04385_));
 sky130_fd_sc_hd__and2_1 _24529_ (.A(net328),
    .B(_04385_),
    .X(_04386_));
 sky130_fd_sc_hd__nor2_1 _24530_ (.A(net328),
    .B(_04385_),
    .Y(_04387_));
 sky130_fd_sc_hd__or3_1 _24531_ (.A(net4001),
    .B(_04386_),
    .C(_04387_),
    .X(_04388_));
 sky130_fd_sc_hd__o221a_1 _24532_ (.A1(_04330_),
    .A2(_04337_),
    .B1(net200),
    .B2(_04383_),
    .C1(net265),
    .X(_04389_));
 sky130_fd_sc_hd__a2bb2o_1 _24533_ (.A1_N(_04329_),
    .A2_N(_04389_),
    .B1(net9066),
    .B2(_02867_),
    .X(_00678_));
 sky130_fd_sc_hd__a21boi_1 _24534_ (.A1(_04331_),
    .A2(_04336_),
    .B1_N(_04332_),
    .Y(_04390_));
 sky130_fd_sc_hd__xnor2_1 _24535_ (.A(net5170),
    .B(\pid_q.prev_int[14] ),
    .Y(_04391_));
 sky130_fd_sc_hd__xnor2_1 _24536_ (.A(_04390_),
    .B(_04391_),
    .Y(_04392_));
 sky130_fd_sc_hd__nand2_1 _24537_ (.A(_04314_),
    .B(_04372_),
    .Y(_04393_));
 sky130_fd_sc_hd__a22o_1 _24538_ (.A1(_04315_),
    .A2(_04373_),
    .B1(_04393_),
    .B2(net792),
    .X(_04394_));
 sky130_fd_sc_hd__a221o_1 _24539_ (.A1(_04373_),
    .A2(_04376_),
    .B1(_04394_),
    .B2(_04268_),
    .C1(_04266_),
    .X(_04395_));
 sky130_fd_sc_hd__a21bo_1 _24540_ (.A1(_04264_),
    .A2(_04374_),
    .B1_N(_04375_),
    .X(_04396_));
 sky130_fd_sc_hd__nor2_1 _24541_ (.A(_04314_),
    .B(_04372_),
    .Y(_04397_));
 sky130_fd_sc_hd__nand2_1 _24542_ (.A(_04372_),
    .B(_04375_),
    .Y(_04398_));
 sky130_fd_sc_hd__a22o_1 _24543_ (.A1(_04373_),
    .A2(_04374_),
    .B1(_04398_),
    .B2(_04264_),
    .X(_04399_));
 sky130_fd_sc_hd__and2_1 _24544_ (.A(_04315_),
    .B(_04399_),
    .X(_04400_));
 sky130_fd_sc_hd__a211o_1 _24545_ (.A1(_04393_),
    .A2(_04396_),
    .B1(_04397_),
    .C1(_04400_),
    .X(_04401_));
 sky130_fd_sc_hd__nand2_1 _24546_ (.A(_04395_),
    .B(_04401_),
    .Y(_04402_));
 sky130_fd_sc_hd__and2_1 _24547_ (.A(net1649),
    .B(_04354_),
    .X(_04403_));
 sky130_fd_sc_hd__nor2_1 _24548_ (.A(net1649),
    .B(_04354_),
    .Y(_04404_));
 sky130_fd_sc_hd__o31a_1 _24549_ (.A1(net1651),
    .A2(_04403_),
    .A3(_04404_),
    .B1(net2018),
    .X(_04405_));
 sky130_fd_sc_hd__o21a_1 _24550_ (.A1(_04357_),
    .A2(_04361_),
    .B1(_04362_),
    .X(_04406_));
 sky130_fd_sc_hd__a21o_1 _24551_ (.A1(_04357_),
    .A2(_04361_),
    .B1(_04406_),
    .X(_04407_));
 sky130_fd_sc_hd__nor2_1 _24552_ (.A(_04405_),
    .B(_04407_),
    .Y(_04408_));
 sky130_fd_sc_hd__nand2_1 _24553_ (.A(_04405_),
    .B(_04407_),
    .Y(_04409_));
 sky130_fd_sc_hd__and2b_1 _24554_ (.A_N(_04408_),
    .B(_04409_),
    .X(_04410_));
 sky130_fd_sc_hd__o21a_1 _24555_ (.A1(_04355_),
    .A2(_04364_),
    .B1(_04339_),
    .X(_04411_));
 sky130_fd_sc_hd__a21oi_1 _24556_ (.A1(_04355_),
    .A2(_04364_),
    .B1(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__a21bo_1 _24557_ (.A1(_04342_),
    .A2(_04353_),
    .B1_N(net1649),
    .X(_04413_));
 sky130_fd_sc_hd__o21a_1 _24558_ (.A1(_04342_),
    .A2(_04353_),
    .B1(_04413_),
    .X(_04414_));
 sky130_fd_sc_hd__inv_2 _24559_ (.A(net4809),
    .Y(_04415_));
 sky130_fd_sc_hd__a21oi_1 _24560_ (.A1(_04415_),
    .A2(_04343_),
    .B1(_04345_),
    .Y(_04416_));
 sky130_fd_sc_hd__a31o_1 _24561_ (.A1(net4523),
    .A2(net4825),
    .A3(net4809),
    .B1(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__nand2_1 _24562_ (.A(net4545),
    .B(_04417_),
    .Y(_04418_));
 sky130_fd_sc_hd__nor2_1 _24563_ (.A(_04343_),
    .B(_04345_),
    .Y(_04419_));
 sky130_fd_sc_hd__or3_1 _24564_ (.A(net4538),
    .B(net3046),
    .C(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__o311a_1 _24565_ (.A1(net4794),
    .A2(_04343_),
    .A3(_04345_),
    .B1(_04418_),
    .C1(_04420_),
    .X(_04421_));
 sky130_fd_sc_hd__xor2_1 _24566_ (.A(net2016),
    .B(_04421_),
    .X(_04422_));
 sky130_fd_sc_hd__xnor2_2 _24567_ (.A(_04414_),
    .B(_04422_),
    .Y(_04423_));
 sky130_fd_sc_hd__nand2_1 _24568_ (.A(net4823),
    .B(net4506),
    .Y(_04424_));
 sky130_fd_sc_hd__nand2_1 _24569_ (.A(net4514),
    .B(net4807),
    .Y(_04425_));
 sky130_fd_sc_hd__nand2_1 _24570_ (.A(net4843),
    .B(net4487),
    .Y(_04426_));
 sky130_fd_sc_hd__xnor2_1 _24571_ (.A(_04425_),
    .B(_04426_),
    .Y(_04427_));
 sky130_fd_sc_hd__xnor2_2 _24572_ (.A(_04424_),
    .B(_04427_),
    .Y(_04428_));
 sky130_fd_sc_hd__a31o_1 _24573_ (.A1(net4919),
    .A2(net4894),
    .A3(net4871),
    .B1(_04351_),
    .X(_04429_));
 sky130_fd_sc_hd__xor2_1 _24574_ (.A(_04428_),
    .B(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__xnor2_1 _24575_ (.A(net4918),
    .B(net4896),
    .Y(_04431_));
 sky130_fd_sc_hd__a21o_1 _24576_ (.A1(net4894),
    .A2(net4871),
    .B1(_04347_),
    .X(_04432_));
 sky130_fd_sc_hd__o311a_1 _24577_ (.A1(_04290_),
    .A2(net4506),
    .A3(_04431_),
    .B1(_04432_),
    .C1(net4491),
    .X(_04433_));
 sky130_fd_sc_hd__a21o_1 _24578_ (.A1(_04347_),
    .A2(_04350_),
    .B1(net4919),
    .X(_04434_));
 sky130_fd_sc_hd__and3_1 _24579_ (.A(_04430_),
    .B(_04433_),
    .C(_04434_),
    .X(_04435_));
 sky130_fd_sc_hd__a21o_1 _24580_ (.A1(_04433_),
    .A2(_04434_),
    .B1(_04430_),
    .X(_04436_));
 sky130_fd_sc_hd__or2b_1 _24581_ (.A(_04435_),
    .B_N(_04436_),
    .X(_04437_));
 sky130_fd_sc_hd__xnor2_2 _24582_ (.A(_04284_),
    .B(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__xor2_1 _24583_ (.A(_04423_),
    .B(_04438_),
    .X(_04439_));
 sky130_fd_sc_hd__xnor2_1 _24584_ (.A(_04412_),
    .B(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__xnor2_2 _24585_ (.A(_04410_),
    .B(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__o21ba_1 _24586_ (.A1(_04368_),
    .A2(_04370_),
    .B1_N(_04366_),
    .X(_04442_));
 sky130_fd_sc_hd__a21o_1 _24587_ (.A1(_04368_),
    .A2(_04370_),
    .B1(_04442_),
    .X(_04443_));
 sky130_fd_sc_hd__xnor2_1 _24588_ (.A(_04441_),
    .B(net631),
    .Y(_04444_));
 sky130_fd_sc_hd__xor2_1 _24589_ (.A(net263),
    .B(_04444_),
    .X(_04445_));
 sky130_fd_sc_hd__and2_1 _24590_ (.A(\pid_q.prev_error[14] ),
    .B(\pid_q.curr_error[14] ),
    .X(_04446_));
 sky130_fd_sc_hd__or2_1 _24591_ (.A(\pid_q.prev_error[14] ),
    .B(\pid_q.curr_error[14] ),
    .X(_04447_));
 sky130_fd_sc_hd__or2b_1 _24592_ (.A(_04446_),
    .B_N(_04447_),
    .X(_04448_));
 sky130_fd_sc_hd__nor2_1 _24593_ (.A(\pid_q.prev_error[13] ),
    .B(net5166),
    .Y(_04449_));
 sky130_fd_sc_hd__nand2_1 _24594_ (.A(\pid_q.prev_error[13] ),
    .B(net5166),
    .Y(_04450_));
 sky130_fd_sc_hd__o21ai_2 _24595_ (.A1(net328),
    .A2(_04449_),
    .B1(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__xor2_1 _24596_ (.A(_04448_),
    .B(_04451_),
    .X(_04452_));
 sky130_fd_sc_hd__nor2_1 _24597_ (.A(_09581_),
    .B(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__a221o_1 _24598_ (.A1(net7522),
    .A2(_04392_),
    .B1(net234),
    .B2(net7465),
    .C1(net230),
    .X(_04454_));
 sky130_fd_sc_hd__a22o_1 _24599_ (.A1(net5170),
    .A2(_02866_),
    .B1(net2433),
    .B2(_04454_),
    .X(_00679_));
 sky130_fd_sc_hd__xor2_1 _24600_ (.A(net5169),
    .B(\pid_q.prev_int[15] ),
    .X(_04455_));
 sky130_fd_sc_hd__and2_1 _24601_ (.A(net5170),
    .B(\pid_q.prev_int[14] ),
    .X(_04456_));
 sky130_fd_sc_hd__or2_1 _24602_ (.A(net5170),
    .B(\pid_q.prev_int[14] ),
    .X(_04457_));
 sky130_fd_sc_hd__o21a_1 _24603_ (.A1(_04390_),
    .A2(_04456_),
    .B1(_04457_),
    .X(_04458_));
 sky130_fd_sc_hd__xnor2_1 _24604_ (.A(_04455_),
    .B(_04458_),
    .Y(_04459_));
 sky130_fd_sc_hd__nand2_1 _24605_ (.A(_04408_),
    .B(_04438_),
    .Y(_04460_));
 sky130_fd_sc_hd__nor2_1 _24606_ (.A(_04409_),
    .B(_04438_),
    .Y(_04461_));
 sky130_fd_sc_hd__nand2_1 _24607_ (.A(_04423_),
    .B(_04461_),
    .Y(_04462_));
 sky130_fd_sc_hd__a21oi_1 _24608_ (.A1(_04409_),
    .A2(_04438_),
    .B1(_04408_),
    .Y(_04463_));
 sky130_fd_sc_hd__o21a_1 _24609_ (.A1(_04423_),
    .A2(_04463_),
    .B1(_04460_),
    .X(_04464_));
 sky130_fd_sc_hd__a21oi_1 _24610_ (.A1(_04423_),
    .A2(_04463_),
    .B1(_04461_),
    .Y(_04465_));
 sky130_fd_sc_hd__mux2_1 _24611_ (.A0(_04464_),
    .A1(_04465_),
    .S(_04412_),
    .X(_04466_));
 sky130_fd_sc_hd__o211a_1 _24612_ (.A1(_04423_),
    .A2(_04460_),
    .B1(_04462_),
    .C1(_04466_),
    .X(_04467_));
 sky130_fd_sc_hd__mux2_1 _24613_ (.A0(net1651),
    .A1(net2018),
    .S(net1649),
    .X(_04468_));
 sky130_fd_sc_hd__nor2_1 _24614_ (.A(net1649),
    .B(_04436_),
    .Y(_04469_));
 sky130_fd_sc_hd__a31o_1 _24615_ (.A1(net1651),
    .A2(net1649),
    .A3(_04435_),
    .B1(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__nand2_1 _24616_ (.A(net2018),
    .B(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__or2_1 _24617_ (.A(net2018),
    .B(net1649),
    .X(_04472_));
 sky130_fd_sc_hd__mux2_1 _24618_ (.A0(net1651),
    .A1(_04472_),
    .S(_04436_),
    .X(_04473_));
 sky130_fd_sc_hd__o211a_1 _24619_ (.A1(_04435_),
    .A2(_04468_),
    .B1(_04471_),
    .C1(_04473_),
    .X(_04474_));
 sky130_fd_sc_hd__inv_2 _24620_ (.A(net4843),
    .Y(_04475_));
 sky130_fd_sc_hd__o31a_1 _24621_ (.A1(net4539),
    .A2(_04475_),
    .A3(_04424_),
    .B1(net4514),
    .X(_04476_));
 sky130_fd_sc_hd__or2_1 _24622_ (.A(net3047),
    .B(_04476_),
    .X(_04477_));
 sky130_fd_sc_hd__nand2_1 _24623_ (.A(net4503),
    .B(net4807),
    .Y(_04478_));
 sky130_fd_sc_hd__o32a_1 _24624_ (.A1(net4823),
    .A2(net4498),
    .A3(_04426_),
    .B1(_04478_),
    .B2(net4490),
    .X(_04479_));
 sky130_fd_sc_hd__a211o_1 _24625_ (.A1(_04296_),
    .A2(net4842),
    .B1(net4823),
    .C1(_04478_),
    .X(_04480_));
 sky130_fd_sc_hd__a211o_1 _24626_ (.A1(net4823),
    .A2(net3745),
    .B1(net4807),
    .C1(_04475_),
    .X(_04481_));
 sky130_fd_sc_hd__a21o_1 _24627_ (.A1(net3745),
    .A2(net4807),
    .B1(_04475_),
    .X(_04482_));
 sky130_fd_sc_hd__a22o_1 _24628_ (.A1(net4514),
    .A2(_04482_),
    .B1(_04478_),
    .B2(_04475_),
    .X(_04483_));
 sky130_fd_sc_hd__nand2_1 _24629_ (.A(net4823),
    .B(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__a21o_1 _24630_ (.A1(_04481_),
    .A2(_04484_),
    .B1(_03705_),
    .X(_04485_));
 sky130_fd_sc_hd__o211a_1 _24631_ (.A1(net4514),
    .A2(_04479_),
    .B1(_04480_),
    .C1(_04485_),
    .X(_04486_));
 sky130_fd_sc_hd__xnor2_1 _24632_ (.A(_04477_),
    .B(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__a21o_1 _24633_ (.A1(net4894),
    .A2(net4871),
    .B1(_04428_),
    .X(_04488_));
 sky130_fd_sc_hd__a22o_1 _24634_ (.A1(_04350_),
    .A2(_04428_),
    .B1(_04488_),
    .B2(net4919),
    .X(_04489_));
 sky130_fd_sc_hd__nand2_1 _24635_ (.A(net4491),
    .B(_04489_),
    .Y(_04490_));
 sky130_fd_sc_hd__xnor2_1 _24636_ (.A(_04487_),
    .B(_04490_),
    .Y(_04491_));
 sky130_fd_sc_hd__xnor2_1 _24637_ (.A(_04474_),
    .B(_04491_),
    .Y(_04492_));
 sky130_fd_sc_hd__or2b_1 _24638_ (.A(_04421_),
    .B_N(_04414_),
    .X(_04493_));
 sky130_fd_sc_hd__and2b_1 _24639_ (.A_N(_04414_),
    .B(_04421_),
    .X(_04494_));
 sky130_fd_sc_hd__a21o_1 _24640_ (.A1(net2016),
    .A2(_04493_),
    .B1(_04494_),
    .X(_04495_));
 sky130_fd_sc_hd__xnor2_1 _24641_ (.A(_04492_),
    .B(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__xnor2_1 _24642_ (.A(_04467_),
    .B(_04496_),
    .Y(_04497_));
 sky130_fd_sc_hd__nor2_1 _24643_ (.A(_04441_),
    .B(net631),
    .Y(_04498_));
 sky130_fd_sc_hd__nand2_1 _24644_ (.A(_04441_),
    .B(net631),
    .Y(_04499_));
 sky130_fd_sc_hd__o21a_1 _24645_ (.A1(net263),
    .A2(_04498_),
    .B1(_04499_),
    .X(_04500_));
 sky130_fd_sc_hd__xor2_1 _24646_ (.A(net509),
    .B(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__xnor2_1 _24647_ (.A(\pid_q.prev_error[15] ),
    .B(\pid_q.curr_error[15] ),
    .Y(_04502_));
 sky130_fd_sc_hd__o21a_1 _24648_ (.A1(_04446_),
    .A2(_04451_),
    .B1(_04447_),
    .X(_04503_));
 sky130_fd_sc_hd__xnor2_1 _24649_ (.A(net3731),
    .B(_04503_),
    .Y(_04504_));
 sky130_fd_sc_hd__nand2_1 _24650_ (.A(net7496),
    .B(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__o221a_1 _24651_ (.A1(_04330_),
    .A2(_04459_),
    .B1(_04501_),
    .B2(_04383_),
    .C1(net195),
    .X(_04506_));
 sky130_fd_sc_hd__a2bb2o_1 _24652_ (.A1_N(_04329_),
    .A2_N(_04506_),
    .B1(net9015),
    .B2(_02867_),
    .X(_00680_));
 sky130_fd_sc_hd__a21o_1 _24653_ (.A1(net7477),
    .A2(net8862),
    .B1(net2146),
    .X(_04507_));
 sky130_fd_sc_hd__buf_1 _24654_ (.A(net1647),
    .X(_04508_));
 sky130_fd_sc_hd__a21oi_1 _24655_ (.A1(net7477),
    .A2(net8874),
    .B1(net2146),
    .Y(_04509_));
 sky130_fd_sc_hd__buf_1 _24656_ (.A(net1645),
    .X(_04510_));
 sky130_fd_sc_hd__and3_1 _24657_ (.A(\pid_q.curr_error[0] ),
    .B(_00011_),
    .C(net1374),
    .X(_04511_));
 sky130_fd_sc_hd__a21o_1 _24658_ (.A1(net9177),
    .A2(net1378),
    .B1(_04511_),
    .X(_00681_));
 sky130_fd_sc_hd__and3_1 _24659_ (.A(net5168),
    .B(_00011_),
    .C(net1374),
    .X(_04512_));
 sky130_fd_sc_hd__a21o_1 _24660_ (.A1(net9228),
    .A2(net1378),
    .B1(_04512_),
    .X(_00682_));
 sky130_fd_sc_hd__and3_1 _24661_ (.A(\pid_q.curr_error[2] ),
    .B(net2382),
    .C(net1372),
    .X(_04513_));
 sky130_fd_sc_hd__a21o_1 _24662_ (.A1(net9178),
    .A2(net1377),
    .B1(_04513_),
    .X(_00683_));
 sky130_fd_sc_hd__and3_1 _24663_ (.A(\pid_q.curr_error[3] ),
    .B(net2382),
    .C(net1372),
    .X(_04514_));
 sky130_fd_sc_hd__a21o_1 _24664_ (.A1(net9175),
    .A2(net1377),
    .B1(_04514_),
    .X(_00684_));
 sky130_fd_sc_hd__and3_1 _24665_ (.A(\pid_q.curr_error[4] ),
    .B(net2382),
    .C(net1372),
    .X(_04515_));
 sky130_fd_sc_hd__a21o_1 _24666_ (.A1(net9139),
    .A2(net1375),
    .B1(_04515_),
    .X(_00685_));
 sky130_fd_sc_hd__and3_1 _24667_ (.A(\pid_q.curr_error[5] ),
    .B(net2383),
    .C(net1373),
    .X(_04516_));
 sky130_fd_sc_hd__a21o_1 _24668_ (.A1(net9144),
    .A2(net1375),
    .B1(_04516_),
    .X(_00686_));
 sky130_fd_sc_hd__and3_1 _24669_ (.A(\pid_q.curr_error[6] ),
    .B(net2383),
    .C(net1373),
    .X(_04517_));
 sky130_fd_sc_hd__a21o_1 _24670_ (.A1(net9145),
    .A2(net1376),
    .B1(_04517_),
    .X(_00687_));
 sky130_fd_sc_hd__and3_1 _24671_ (.A(\pid_q.curr_error[7] ),
    .B(net2384),
    .C(net1373),
    .X(_04518_));
 sky130_fd_sc_hd__a21o_1 _24672_ (.A1(net9123),
    .A2(net1376),
    .B1(_04518_),
    .X(_00688_));
 sky130_fd_sc_hd__and3_1 _24673_ (.A(\pid_q.curr_error[8] ),
    .B(_00011_),
    .C(net1374),
    .X(_04519_));
 sky130_fd_sc_hd__a21o_1 _24674_ (.A1(net9142),
    .A2(net1378),
    .B1(_04519_),
    .X(_00689_));
 sky130_fd_sc_hd__and3_1 _24675_ (.A(\pid_q.curr_error[9] ),
    .B(net3019),
    .C(_04510_),
    .X(_04520_));
 sky130_fd_sc_hd__a21o_1 _24676_ (.A1(net9133),
    .A2(_04508_),
    .B1(_04520_),
    .X(_00690_));
 sky130_fd_sc_hd__and3_1 _24677_ (.A(\pid_q.curr_error[10] ),
    .B(net3020),
    .C(net1645),
    .X(_04521_));
 sky130_fd_sc_hd__a21o_1 _24678_ (.A1(net9127),
    .A2(net1648),
    .B1(_04521_),
    .X(_00691_));
 sky130_fd_sc_hd__and3_1 _24679_ (.A(\pid_q.curr_error[11] ),
    .B(net3021),
    .C(net1646),
    .X(_04522_));
 sky130_fd_sc_hd__a21o_1 _24680_ (.A1(net9184),
    .A2(net1647),
    .B1(_04522_),
    .X(_00692_));
 sky130_fd_sc_hd__and3_1 _24681_ (.A(net5167),
    .B(net3021),
    .C(net1646),
    .X(_04523_));
 sky130_fd_sc_hd__a21o_1 _24682_ (.A1(net9032),
    .A2(net1647),
    .B1(_04523_),
    .X(_00693_));
 sky130_fd_sc_hd__and3_1 _24683_ (.A(net5166),
    .B(net3021),
    .C(_04509_),
    .X(_04524_));
 sky130_fd_sc_hd__a21o_1 _24684_ (.A1(net9179),
    .A2(_04507_),
    .B1(_04524_),
    .X(_00694_));
 sky130_fd_sc_hd__and3_1 _24685_ (.A(\pid_q.curr_error[14] ),
    .B(net3021),
    .C(_04509_),
    .X(_04525_));
 sky130_fd_sc_hd__a21o_1 _24686_ (.A1(net9067),
    .A2(_04507_),
    .B1(_04525_),
    .X(_00695_));
 sky130_fd_sc_hd__and3_1 _24687_ (.A(\pid_q.curr_error[15] ),
    .B(net3020),
    .C(net1646),
    .X(_04526_));
 sky130_fd_sc_hd__a21o_1 _24688_ (.A1(net9107),
    .A2(net1648),
    .B1(_04526_),
    .X(_00696_));
 sky130_fd_sc_hd__o21a_1 _24689_ (.A1(net7475),
    .A2(net3269),
    .B1(net8875),
    .X(_04527_));
 sky130_fd_sc_hd__or2_1 _24690_ (.A(net3715),
    .B(_04527_),
    .X(_04528_));
 sky130_fd_sc_hd__buf_1 _24691_ (.A(_04528_),
    .X(_04529_));
 sky130_fd_sc_hd__buf_1 _24692_ (.A(net1643),
    .X(_04530_));
 sky130_fd_sc_hd__inv_2 _24693_ (.A(net7490),
    .Y(_04531_));
 sky130_fd_sc_hd__xnor2_1 _24694_ (.A(net8034),
    .B(net4265),
    .Y(_04532_));
 sky130_fd_sc_hd__nor2_1 _24695_ (.A(net3727),
    .B(net3034),
    .Y(_04533_));
 sky130_fd_sc_hd__or2_1 _24696_ (.A(net4310),
    .B(net3269),
    .X(_04534_));
 sky130_fd_sc_hd__nor2_1 _24697_ (.A(net7501),
    .B(_04534_),
    .Y(_04535_));
 sky130_fd_sc_hd__a22o_1 _24698_ (.A1(\pid_q.curr_error[0] ),
    .A2(net1370),
    .B1(_04533_),
    .B2(net2015),
    .X(_00697_));
 sky130_fd_sc_hd__or2b_1 _24699_ (.A(net8034),
    .B_N(net5307),
    .X(_04536_));
 sky130_fd_sc_hd__xnor2_1 _24700_ (.A(net5299),
    .B(_04536_),
    .Y(_04537_));
 sky130_fd_sc_hd__nand2_1 _24701_ (.A(net1621),
    .B(_04537_),
    .Y(_04538_));
 sky130_fd_sc_hd__xnor2_1 _24702_ (.A(net8028),
    .B(_04538_),
    .Y(_04539_));
 sky130_fd_sc_hd__nor2_2 _24703_ (.A(net4310),
    .B(net3269),
    .Y(_04540_));
 sky130_fd_sc_hd__and3_1 _24704_ (.A(net7488),
    .B(net4000),
    .C(_04540_),
    .X(_04541_));
 sky130_fd_sc_hd__buf_1 _24705_ (.A(_04541_),
    .X(_04542_));
 sky130_fd_sc_hd__a22o_1 _24706_ (.A1(net9055),
    .A2(_04530_),
    .B1(net1011),
    .B2(net1642),
    .X(_00698_));
 sky130_fd_sc_hd__buf_1 _24707_ (.A(net1642),
    .X(_04543_));
 sky130_fd_sc_hd__or2b_1 _24708_ (.A(net8028),
    .B_N(net5299),
    .X(_04544_));
 sky130_fd_sc_hd__and2b_1 _24709_ (.A_N(net5299),
    .B(net8028),
    .X(_04545_));
 sky130_fd_sc_hd__a21o_1 _24710_ (.A1(_04536_),
    .A2(_04544_),
    .B1(_04545_),
    .X(_04546_));
 sky130_fd_sc_hd__xnor2_1 _24711_ (.A(net5290),
    .B(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__nand2_1 _24712_ (.A(net1621),
    .B(_04547_),
    .Y(_04548_));
 sky130_fd_sc_hd__xnor2_1 _24713_ (.A(net8023),
    .B(net1158),
    .Y(_04549_));
 sky130_fd_sc_hd__a22o_1 _24714_ (.A1(\pid_q.curr_error[2] ),
    .A2(net1368),
    .B1(net1365),
    .B2(net1010),
    .X(_00699_));
 sky130_fd_sc_hd__a21bo_1 _24715_ (.A1(net8022),
    .A2(_04546_),
    .B1_N(net5290),
    .X(_04550_));
 sky130_fd_sc_hd__or2_1 _24716_ (.A(net8022),
    .B(_04546_),
    .X(_04551_));
 sky130_fd_sc_hd__a21o_1 _24717_ (.A1(_04550_),
    .A2(_04551_),
    .B1(net4232),
    .X(_04552_));
 sky130_fd_sc_hd__xor2_1 _24718_ (.A(net8017),
    .B(net4268),
    .X(_04553_));
 sky130_fd_sc_hd__xnor2_1 _24719_ (.A(_04552_),
    .B(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__a22o_1 _24720_ (.A1(\pid_q.curr_error[3] ),
    .A2(net1368),
    .B1(net1365),
    .B2(net1640),
    .X(_00700_));
 sky130_fd_sc_hd__inv_2 _24721_ (.A(net5283),
    .Y(_04555_));
 sky130_fd_sc_hd__a21o_1 _24722_ (.A1(net8017),
    .A2(_04552_),
    .B1(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__a211o_1 _24723_ (.A1(_04550_),
    .A2(_04551_),
    .B1(net8017),
    .C1(net4232),
    .X(_04557_));
 sky130_fd_sc_hd__a21oi_1 _24724_ (.A1(_04556_),
    .A2(_04557_),
    .B1(net5273),
    .Y(_04558_));
 sky130_fd_sc_hd__and3_1 _24725_ (.A(net5273),
    .B(_04556_),
    .C(_04557_),
    .X(_04559_));
 sky130_fd_sc_hd__o21a_1 _24726_ (.A1(_04558_),
    .A2(_04559_),
    .B1(net1988),
    .X(_04560_));
 sky130_fd_sc_hd__xor2_1 _24727_ (.A(net8012),
    .B(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__a22o_1 _24728_ (.A1(\pid_q.curr_error[4] ),
    .A2(net1368),
    .B1(net1365),
    .B2(_04561_),
    .X(_00701_));
 sky130_fd_sc_hd__inv_2 _24729_ (.A(net5273),
    .Y(_04562_));
 sky130_fd_sc_hd__a21o_1 _24730_ (.A1(net8012),
    .A2(_04557_),
    .B1(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__a221o_1 _24731_ (.A1(_04562_),
    .A2(net8012),
    .B1(_04552_),
    .B2(net8017),
    .C1(_04555_),
    .X(_04564_));
 sky130_fd_sc_hd__a21o_1 _24732_ (.A1(_04563_),
    .A2(_04564_),
    .B1(net4232),
    .X(_04565_));
 sky130_fd_sc_hd__or2_1 _24733_ (.A(net8012),
    .B(_04557_),
    .X(_04566_));
 sky130_fd_sc_hd__and2_1 _24734_ (.A(_04565_),
    .B(_04566_),
    .X(_04567_));
 sky130_fd_sc_hd__xor2_1 _24735_ (.A(net8007),
    .B(net4272),
    .X(_04568_));
 sky130_fd_sc_hd__xnor2_1 _24736_ (.A(_04567_),
    .B(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__a22o_1 _24737_ (.A1(\pid_q.curr_error[5] ),
    .A2(net1371),
    .B1(net1365),
    .B2(net1009),
    .X(_00702_));
 sky130_fd_sc_hd__inv_2 _24738_ (.A(net5265),
    .Y(_04570_));
 sky130_fd_sc_hd__and3_1 _24739_ (.A(net8007),
    .B(_04565_),
    .C(_04566_),
    .X(_04571_));
 sky130_fd_sc_hd__or2_1 _24740_ (.A(net8007),
    .B(_04567_),
    .X(_04572_));
 sky130_fd_sc_hd__o21a_1 _24741_ (.A1(_04570_),
    .A2(_04571_),
    .B1(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__xnor2_1 _24742_ (.A(net5259),
    .B(_04573_),
    .Y(_04574_));
 sky130_fd_sc_hd__nand2_1 _24743_ (.A(net1988),
    .B(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__xnor2_1 _24744_ (.A(net8002),
    .B(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hd__a22o_1 _24745_ (.A1(\pid_q.curr_error[6] ),
    .A2(net1371),
    .B1(net1366),
    .B2(net738),
    .X(_00703_));
 sky130_fd_sc_hd__inv_2 _24746_ (.A(net5259),
    .Y(_04577_));
 sky130_fd_sc_hd__a21o_1 _24747_ (.A1(net8002),
    .A2(_04572_),
    .B1(_04577_),
    .X(_04578_));
 sky130_fd_sc_hd__a211o_1 _24748_ (.A1(_04577_),
    .A2(net8002),
    .B1(_04571_),
    .C1(_04570_),
    .X(_04579_));
 sky130_fd_sc_hd__a21o_1 _24749_ (.A1(_04578_),
    .A2(_04579_),
    .B1(net4232),
    .X(_04580_));
 sky130_fd_sc_hd__or2_1 _24750_ (.A(net8002),
    .B(_04572_),
    .X(_04581_));
 sky130_fd_sc_hd__nand2_1 _24751_ (.A(_04580_),
    .B(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__nand2_1 _24752_ (.A(net5254),
    .B(net3031),
    .Y(_04583_));
 sky130_fd_sc_hd__xor2_1 _24753_ (.A(net7996),
    .B(net2009),
    .X(_04584_));
 sky130_fd_sc_hd__xnor2_1 _24754_ (.A(_04582_),
    .B(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__a22o_1 _24755_ (.A1(\pid_q.curr_error[7] ),
    .A2(net1369),
    .B1(net1366),
    .B2(net737),
    .X(_00704_));
 sky130_fd_sc_hd__a21o_1 _24756_ (.A1(_04580_),
    .A2(_04581_),
    .B1(net7996),
    .X(_04586_));
 sky130_fd_sc_hd__a31o_1 _24757_ (.A1(net7996),
    .A2(_04580_),
    .A3(_04581_),
    .B1(net2009),
    .X(_04587_));
 sky130_fd_sc_hd__and2_1 _24758_ (.A(_04586_),
    .B(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__nand2_1 _24759_ (.A(net5245),
    .B(net2390),
    .Y(_04589_));
 sky130_fd_sc_hd__xnor2_1 _24760_ (.A(net7990),
    .B(net1638),
    .Y(_04590_));
 sky130_fd_sc_hd__xnor2_1 _24761_ (.A(_04588_),
    .B(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__a22o_1 _24762_ (.A1(\pid_q.curr_error[8] ),
    .A2(net1368),
    .B1(net1367),
    .B2(net690),
    .X(_00705_));
 sky130_fd_sc_hd__a31o_1 _24763_ (.A1(net7990),
    .A2(_04586_),
    .A3(_04587_),
    .B1(net1638),
    .X(_04592_));
 sky130_fd_sc_hd__o21ai_2 _24764_ (.A1(net7990),
    .A2(_04588_),
    .B1(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__xnor2_1 _24765_ (.A(net7985),
    .B(net4256),
    .Y(_04594_));
 sky130_fd_sc_hd__xnor2_1 _24766_ (.A(_04593_),
    .B(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__a22o_1 _24767_ (.A1(\pid_q.curr_error[9] ),
    .A2(net1370),
    .B1(net1367),
    .B2(net629),
    .X(_00706_));
 sky130_fd_sc_hd__inv_2 _24768_ (.A(net7985),
    .Y(_04596_));
 sky130_fd_sc_hd__o21ai_1 _24769_ (.A1(_04596_),
    .A2(_04593_),
    .B1(net5235),
    .Y(_04597_));
 sky130_fd_sc_hd__nand2_1 _24770_ (.A(_04596_),
    .B(_04593_),
    .Y(_04598_));
 sky130_fd_sc_hd__a21oi_1 _24771_ (.A1(_04597_),
    .A2(_04598_),
    .B1(net5220),
    .Y(_04599_));
 sky130_fd_sc_hd__and3_1 _24772_ (.A(net5220),
    .B(_04597_),
    .C(_04598_),
    .X(_04600_));
 sky130_fd_sc_hd__o21ai_1 _24773_ (.A1(_04599_),
    .A2(_04600_),
    .B1(net1988),
    .Y(_04601_));
 sky130_fd_sc_hd__xor2_1 _24774_ (.A(net7980),
    .B(_04601_),
    .X(_04602_));
 sky130_fd_sc_hd__inv_2 _24775_ (.A(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__a32o_1 _24776_ (.A1(net7479),
    .A2(_04535_),
    .A3(net457),
    .B1(net9193),
    .B2(_04529_),
    .X(_00707_));
 sky130_fd_sc_hd__and2b_1 _24777_ (.A_N(net5228),
    .B(net7980),
    .X(_04604_));
 sky130_fd_sc_hd__nand2_1 _24778_ (.A(net7980),
    .B(_04598_),
    .Y(_04605_));
 sky130_fd_sc_hd__a2bb2o_1 _24779_ (.A1_N(_04604_),
    .A2_N(_04597_),
    .B1(net5220),
    .B2(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__a2bb2o_1 _24780_ (.A1_N(net7980),
    .A2_N(_04598_),
    .B1(_04606_),
    .B2(net2385),
    .X(_04607_));
 sky130_fd_sc_hd__inv_2 _24781_ (.A(net7974),
    .Y(_04608_));
 sky130_fd_sc_hd__nand2_1 _24782_ (.A(net5214),
    .B(net2390),
    .Y(_04609_));
 sky130_fd_sc_hd__xnor2_1 _24783_ (.A(_04608_),
    .B(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__xnor2_1 _24784_ (.A(_04607_),
    .B(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__a22o_1 _24785_ (.A1(\pid_q.curr_error[11] ),
    .A2(net1643),
    .B1(_04543_),
    .B2(net455),
    .X(_00708_));
 sky130_fd_sc_hd__a21bo_1 _24786_ (.A1(_04608_),
    .A2(_04607_),
    .B1_N(_04609_),
    .X(_04612_));
 sky130_fd_sc_hd__o21a_1 _24787_ (.A1(_04608_),
    .A2(_04607_),
    .B1(_04612_),
    .X(_04613_));
 sky130_fd_sc_hd__inv_2 _24788_ (.A(net7967),
    .Y(_04614_));
 sky130_fd_sc_hd__nand2_1 _24789_ (.A(net5206),
    .B(net1987),
    .Y(_04615_));
 sky130_fd_sc_hd__xnor2_1 _24790_ (.A(_04614_),
    .B(_04615_),
    .Y(_04616_));
 sky130_fd_sc_hd__xnor2_1 _24791_ (.A(_04613_),
    .B(_04616_),
    .Y(_04617_));
 sky130_fd_sc_hd__a22o_1 _24792_ (.A1(net5167),
    .A2(net1643),
    .B1(_04543_),
    .B2(net372),
    .X(_00709_));
 sky130_fd_sc_hd__inv_2 _24793_ (.A(net5198),
    .Y(_04618_));
 sky130_fd_sc_hd__o21ai_1 _24794_ (.A1(_04614_),
    .A2(_04613_),
    .B1(net5206),
    .Y(_04619_));
 sky130_fd_sc_hd__nand2_1 _24795_ (.A(_04614_),
    .B(_04613_),
    .Y(_04620_));
 sky130_fd_sc_hd__and3_1 _24796_ (.A(_04618_),
    .B(_04619_),
    .C(_04620_),
    .X(_04621_));
 sky130_fd_sc_hd__a21oi_1 _24797_ (.A1(_04619_),
    .A2(_04620_),
    .B1(_04618_),
    .Y(_04622_));
 sky130_fd_sc_hd__or3_1 _24798_ (.A(net2883),
    .B(_04621_),
    .C(_04622_),
    .X(_04623_));
 sky130_fd_sc_hd__xor2_1 _24799_ (.A(net7961),
    .B(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__inv_2 _24800_ (.A(net259),
    .Y(_04625_));
 sky130_fd_sc_hd__a22o_1 _24801_ (.A1(net8983),
    .A2(net1644),
    .B1(_04542_),
    .B2(_04625_),
    .X(_00710_));
 sky130_fd_sc_hd__a211o_1 _24802_ (.A1(net7961),
    .A2(_04620_),
    .B1(_06533_),
    .C1(_04618_),
    .X(_04626_));
 sky130_fd_sc_hd__a211o_1 _24803_ (.A1(_04618_),
    .A2(net7961),
    .B1(_06533_),
    .C1(_04619_),
    .X(_04627_));
 sky130_fd_sc_hd__o211a_1 _24804_ (.A1(net7961),
    .A2(_04620_),
    .B1(_04626_),
    .C1(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__nand2_1 _24805_ (.A(net5194),
    .B(net2385),
    .Y(_04629_));
 sky130_fd_sc_hd__xor2_1 _24806_ (.A(net7955),
    .B(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__xnor2_1 _24807_ (.A(_04628_),
    .B(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__inv_2 _24808_ (.A(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__a22o_1 _24809_ (.A1(net9151),
    .A2(net1644),
    .B1(_04542_),
    .B2(net227),
    .X(_00711_));
 sky130_fd_sc_hd__or2_1 _24810_ (.A(net7955),
    .B(_04628_),
    .X(_04633_));
 sky130_fd_sc_hd__a21o_1 _24811_ (.A1(net5189),
    .A2(_04633_),
    .B1(net5194),
    .X(_04634_));
 sky130_fd_sc_hd__nand2_1 _24812_ (.A(net5194),
    .B(net5189),
    .Y(_04635_));
 sky130_fd_sc_hd__nand2_1 _24813_ (.A(net7955),
    .B(_04628_),
    .Y(_04636_));
 sky130_fd_sc_hd__mux2_1 _24814_ (.A0(net5189),
    .A1(_04635_),
    .S(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__a21oi_1 _24815_ (.A1(net5189),
    .A2(net1989),
    .B1(_04633_),
    .Y(_04638_));
 sky130_fd_sc_hd__a31oi_1 _24816_ (.A1(net1626),
    .A2(_04634_),
    .A3(_04637_),
    .B1(_04638_),
    .Y(_04639_));
 sky130_fd_sc_hd__xnor2_1 _24817_ (.A(net7949),
    .B(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__a22o_1 _24818_ (.A1(net9164),
    .A2(net1644),
    .B1(_04542_),
    .B2(net175),
    .X(_00712_));
 sky130_fd_sc_hd__clkbuf_1 _24819_ (.A(net2403),
    .X(_04641_));
 sky130_fd_sc_hd__buf_2 _24820_ (.A(net2008),
    .X(_04642_));
 sky130_fd_sc_hd__clkbuf_1 _24821_ (.A(_04540_),
    .X(_04643_));
 sky130_fd_sc_hd__or2_1 _24822_ (.A(_03313_),
    .B(_04533_),
    .X(_04644_));
 sky130_fd_sc_hd__a22o_1 _24823_ (.A1(net5156),
    .A2(_04642_),
    .B1(net2000),
    .B2(_04644_),
    .X(_00713_));
 sky130_fd_sc_hd__a21o_1 _24824_ (.A1(net7482),
    .A2(net1011),
    .B1(net2419),
    .X(_04645_));
 sky130_fd_sc_hd__a22o_1 _24825_ (.A1(net5117),
    .A2(_04642_),
    .B1(net2000),
    .B2(net927),
    .X(_00714_));
 sky130_fd_sc_hd__a21o_1 _24826_ (.A1(net7480),
    .A2(net1010),
    .B1(net2416),
    .X(_04646_));
 sky130_fd_sc_hd__a22o_1 _24827_ (.A1(net5091),
    .A2(_04642_),
    .B1(net2000),
    .B2(net926),
    .X(_00715_));
 sky130_fd_sc_hd__a21o_1 _24828_ (.A1(net7480),
    .A2(net1640),
    .B1(_03575_),
    .X(_04647_));
 sky130_fd_sc_hd__a22o_1 _24829_ (.A1(net5072),
    .A2(_04642_),
    .B1(net2000),
    .B2(net1363),
    .X(_00716_));
 sky130_fd_sc_hd__a21o_1 _24830_ (.A1(net7480),
    .A2(_04561_),
    .B1(net1383),
    .X(_04648_));
 sky130_fd_sc_hd__a22o_1 _24831_ (.A1(net5043),
    .A2(_04642_),
    .B1(net2000),
    .B2(net924),
    .X(_00717_));
 sky130_fd_sc_hd__a21o_1 _24832_ (.A1(net7484),
    .A2(net1009),
    .B1(net1017),
    .X(_04649_));
 sky130_fd_sc_hd__a22o_1 _24833_ (.A1(net5021),
    .A2(_04642_),
    .B1(net2000),
    .B2(net922),
    .X(_00718_));
 sky130_fd_sc_hd__a21o_1 _24834_ (.A1(net7481),
    .A2(net738),
    .B1(net854),
    .X(_04650_));
 sky130_fd_sc_hd__a22o_1 _24835_ (.A1(net4988),
    .A2(_04642_),
    .B1(net2001),
    .B2(net688),
    .X(_00719_));
 sky130_fd_sc_hd__a21o_1 _24836_ (.A1(net7481),
    .A2(net737),
    .B1(_03952_),
    .X(_04651_));
 sky130_fd_sc_hd__a22o_1 _24837_ (.A1(net4956),
    .A2(_04642_),
    .B1(net2001),
    .B2(net686),
    .X(_00720_));
 sky130_fd_sc_hd__a21o_1 _24838_ (.A1(net7482),
    .A2(net690),
    .B1(_04035_),
    .X(_04652_));
 sky130_fd_sc_hd__a22o_1 _24839_ (.A1(net4933),
    .A2(net2008),
    .B1(net2001),
    .B2(net586),
    .X(_00721_));
 sky130_fd_sc_hd__a21o_1 _24840_ (.A1(net7482),
    .A2(net629),
    .B1(_04115_),
    .X(_04653_));
 sky130_fd_sc_hd__a22o_1 _24841_ (.A1(net4916),
    .A2(net2008),
    .B1(net2001),
    .B2(net508),
    .X(_00722_));
 sky130_fd_sc_hd__a21oi_1 _24842_ (.A1(net7479),
    .A2(net457),
    .B1(_04184_),
    .Y(_04654_));
 sky130_fd_sc_hd__a2bb2o_1 _24843_ (.A1_N(_04534_),
    .A2_N(_04654_),
    .B1(net4897),
    .B2(_04642_),
    .X(_00723_));
 sky130_fd_sc_hd__a21o_1 _24844_ (.A1(net7485),
    .A2(net455),
    .B1(_04257_),
    .X(_04655_));
 sky130_fd_sc_hd__a22o_1 _24845_ (.A1(net4874),
    .A2(net2007),
    .B1(_04540_),
    .B2(net327),
    .X(_00724_));
 sky130_fd_sc_hd__a21o_1 _24846_ (.A1(net7486),
    .A2(net372),
    .B1(_04327_),
    .X(_04656_));
 sky130_fd_sc_hd__a22o_1 _24847_ (.A1(net4841),
    .A2(net2007),
    .B1(_04540_),
    .B2(net258),
    .X(_00725_));
 sky130_fd_sc_hd__o21a_1 _24848_ (.A1(net3727),
    .A2(net259),
    .B1(net264),
    .X(_04657_));
 sky130_fd_sc_hd__a2bb2o_1 _24849_ (.A1_N(_04534_),
    .A2_N(_04657_),
    .B1(net4821),
    .B2(_04642_),
    .X(_00726_));
 sky130_fd_sc_hd__and3_1 _24850_ (.A(net7488),
    .B(_04540_),
    .C(net227),
    .X(_04658_));
 sky130_fd_sc_hd__a221o_1 _24851_ (.A1(net4806),
    .A2(net2007),
    .B1(_04540_),
    .B2(net231),
    .C1(_04658_),
    .X(_00727_));
 sky130_fd_sc_hd__a32o_1 _24852_ (.A1(net7502),
    .A2(_04504_),
    .A3(_04540_),
    .B1(net2007),
    .B2(net4787),
    .X(_04659_));
 sky130_fd_sc_hd__a31o_1 _24853_ (.A1(net7488),
    .A2(_04540_),
    .A3(net175),
    .B1(_04659_),
    .X(_00728_));
 sky130_fd_sc_hd__a22o_1 _24854_ (.A1(\pid_q.ki[0] ),
    .A2(net3022),
    .B1(net3007),
    .B2(\pid_q.kp[0] ),
    .X(_04660_));
 sky130_fd_sc_hd__mux2_1 _24855_ (.A0(_04660_),
    .A1(net4779),
    .S(net2003),
    .X(_04661_));
 sky130_fd_sc_hd__clkbuf_1 _24856_ (.A(_04661_),
    .X(_00729_));
 sky130_fd_sc_hd__a22o_1 _24857_ (.A1(\pid_q.ki[1] ),
    .A2(net3022),
    .B1(net3007),
    .B2(\pid_q.kp[1] ),
    .X(_04662_));
 sky130_fd_sc_hd__mux2_1 _24858_ (.A0(_04662_),
    .A1(net4767),
    .S(net2003),
    .X(_04663_));
 sky130_fd_sc_hd__clkbuf_1 _24859_ (.A(_04663_),
    .X(_00730_));
 sky130_fd_sc_hd__clkbuf_1 _24860_ (.A(net3710),
    .X(_04664_));
 sky130_fd_sc_hd__a22o_1 _24861_ (.A1(\pid_q.ki[2] ),
    .A2(net2397),
    .B1(net3009),
    .B2(\pid_q.kp[2] ),
    .X(_04665_));
 sky130_fd_sc_hd__mux2_1 _24862_ (.A0(net1999),
    .A1(net4744),
    .S(net2002),
    .X(_04666_));
 sky130_fd_sc_hd__clkbuf_1 _24863_ (.A(_04666_),
    .X(_00731_));
 sky130_fd_sc_hd__a22o_1 _24864_ (.A1(\pid_q.ki[3] ),
    .A2(net2398),
    .B1(net3008),
    .B2(\pid_q.kp[3] ),
    .X(_04667_));
 sky130_fd_sc_hd__clkbuf_1 _24865_ (.A(net2399),
    .X(_04668_));
 sky130_fd_sc_hd__mux2_1 _24866_ (.A0(_04667_),
    .A1(net4724),
    .S(net1997),
    .X(_04669_));
 sky130_fd_sc_hd__clkbuf_1 _24867_ (.A(_04669_),
    .X(_00732_));
 sky130_fd_sc_hd__a22o_1 _24868_ (.A1(\pid_q.ki[4] ),
    .A2(net2398),
    .B1(_00008_),
    .B2(\pid_q.kp[4] ),
    .X(_04670_));
 sky130_fd_sc_hd__mux2_1 _24869_ (.A0(_04670_),
    .A1(net4707),
    .S(net1996),
    .X(_04671_));
 sky130_fd_sc_hd__clkbuf_1 _24870_ (.A(_04671_),
    .X(_00733_));
 sky130_fd_sc_hd__a22o_1 _24871_ (.A1(net4481),
    .A2(net2397),
    .B1(net3009),
    .B2(net4478),
    .X(_04672_));
 sky130_fd_sc_hd__mux2_1 _24872_ (.A0(_04672_),
    .A1(net4687),
    .S(net1996),
    .X(_04673_));
 sky130_fd_sc_hd__clkbuf_1 _24873_ (.A(_04673_),
    .X(_00734_));
 sky130_fd_sc_hd__a22o_1 _24874_ (.A1(\pid_q.ki[6] ),
    .A2(net2397),
    .B1(net3009),
    .B2(\pid_q.kp[6] ),
    .X(_04674_));
 sky130_fd_sc_hd__mux2_1 _24875_ (.A0(_04674_),
    .A1(net4646),
    .S(net1996),
    .X(_04675_));
 sky130_fd_sc_hd__clkbuf_1 _24876_ (.A(_04675_),
    .X(_00735_));
 sky130_fd_sc_hd__a22o_1 _24877_ (.A1(\pid_q.ki[7] ),
    .A2(net2397),
    .B1(net3009),
    .B2(\pid_q.kp[7] ),
    .X(_04676_));
 sky130_fd_sc_hd__mux2_1 _24878_ (.A0(_04676_),
    .A1(net4630),
    .S(net1996),
    .X(_04677_));
 sky130_fd_sc_hd__clkbuf_1 _24879_ (.A(_04677_),
    .X(_00736_));
 sky130_fd_sc_hd__a22o_1 _24880_ (.A1(\pid_q.ki[8] ),
    .A2(net2397),
    .B1(net3009),
    .B2(\pid_q.kp[8] ),
    .X(_04678_));
 sky130_fd_sc_hd__mux2_1 _24881_ (.A0(_04678_),
    .A1(net4602),
    .S(net1996),
    .X(_04679_));
 sky130_fd_sc_hd__clkbuf_1 _24882_ (.A(_04679_),
    .X(_00737_));
 sky130_fd_sc_hd__a22o_1 _24883_ (.A1(net4479),
    .A2(net2397),
    .B1(net3699),
    .B2(net4476),
    .X(_04680_));
 sky130_fd_sc_hd__mux2_1 _24884_ (.A0(_04680_),
    .A1(net4594),
    .S(net1996),
    .X(_04681_));
 sky130_fd_sc_hd__clkbuf_1 _24885_ (.A(_04681_),
    .X(_00738_));
 sky130_fd_sc_hd__a22o_1 _24886_ (.A1(\pid_q.ki[10] ),
    .A2(net2398),
    .B1(net3700),
    .B2(\pid_q.kp[10] ),
    .X(_04682_));
 sky130_fd_sc_hd__mux2_1 _24887_ (.A0(_04682_),
    .A1(net4570),
    .S(net1997),
    .X(_04683_));
 sky130_fd_sc_hd__clkbuf_1 _24888_ (.A(_04683_),
    .X(_00739_));
 sky130_fd_sc_hd__a22o_1 _24889_ (.A1(\pid_q.ki[11] ),
    .A2(net2398),
    .B1(net3700),
    .B2(\pid_q.kp[11] ),
    .X(_04684_));
 sky130_fd_sc_hd__mux2_1 _24890_ (.A0(_04684_),
    .A1(net4556),
    .S(net1997),
    .X(_04685_));
 sky130_fd_sc_hd__clkbuf_1 _24891_ (.A(_04685_),
    .X(_00740_));
 sky130_fd_sc_hd__a22o_1 _24892_ (.A1(\pid_q.ki[12] ),
    .A2(net3710),
    .B1(net3700),
    .B2(\pid_q.kp[12] ),
    .X(_04686_));
 sky130_fd_sc_hd__mux2_1 _24893_ (.A0(_04686_),
    .A1(\pid_q.mult0.a[12] ),
    .S(net1998),
    .X(_04687_));
 sky130_fd_sc_hd__clkbuf_1 _24894_ (.A(_04687_),
    .X(_00741_));
 sky130_fd_sc_hd__a22o_1 _24895_ (.A1(\pid_q.ki[13] ),
    .A2(net3711),
    .B1(net3701),
    .B2(\pid_q.kp[13] ),
    .X(_04688_));
 sky130_fd_sc_hd__mux2_1 _24896_ (.A0(_04688_),
    .A1(net4525),
    .S(net2399),
    .X(_04689_));
 sky130_fd_sc_hd__clkbuf_1 _24897_ (.A(_04689_),
    .X(_00742_));
 sky130_fd_sc_hd__a22o_1 _24898_ (.A1(\pid_q.ki[14] ),
    .A2(net3711),
    .B1(net3701),
    .B2(\pid_q.kp[14] ),
    .X(_04690_));
 sky130_fd_sc_hd__mux2_1 _24899_ (.A0(_04690_),
    .A1(net4507),
    .S(net2399),
    .X(_04691_));
 sky130_fd_sc_hd__clkbuf_1 _24900_ (.A(_04691_),
    .X(_00743_));
 sky130_fd_sc_hd__a22o_1 _24901_ (.A1(\pid_q.ki[15] ),
    .A2(net3711),
    .B1(net3701),
    .B2(net4475),
    .X(_04692_));
 sky130_fd_sc_hd__mux2_1 _24902_ (.A0(_04692_),
    .A1(net4492),
    .S(net2399),
    .X(_04693_));
 sky130_fd_sc_hd__clkbuf_1 _24903_ (.A(_04693_),
    .X(_00744_));
 sky130_fd_sc_hd__and2b_1 _24904_ (.A_N(net8871),
    .B(net130),
    .X(_04694_));
 sky130_fd_sc_hd__or4_1 _24905_ (.A(net129),
    .B(net8885),
    .C(net116),
    .D(net119),
    .X(_04695_));
 sky130_fd_sc_hd__or4_1 _24906_ (.A(net115),
    .B(net118),
    .C(net117),
    .D(net120),
    .X(_04696_));
 sky130_fd_sc_hd__or4_1 _24907_ (.A(net8869),
    .B(net121),
    .C(net123),
    .D(net126),
    .X(_04697_));
 sky130_fd_sc_hd__or4_1 _24908_ (.A(net122),
    .B(net125),
    .C(net124),
    .D(net8886),
    .X(_04698_));
 sky130_fd_sc_hd__or4_1 _24909_ (.A(_04695_),
    .B(_04696_),
    .C(_04697_),
    .D(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__inv_2 _24910_ (.A(_04699_),
    .Y(_04700_));
 sky130_fd_sc_hd__a22o_1 _24911_ (.A1(net3730),
    .A2(net2011),
    .B1(_04700_),
    .B2(net114),
    .X(_04701_));
 sky130_fd_sc_hd__buf_1 _24912_ (.A(net1636),
    .X(_04702_));
 sky130_fd_sc_hd__mux2_1 _24913_ (.A0(\pid_q.ki[0] ),
    .A1(_04694_),
    .S(_04702_),
    .X(_04703_));
 sky130_fd_sc_hd__clkbuf_1 _24914_ (.A(_04703_),
    .X(_00745_));
 sky130_fd_sc_hd__and2b_1 _24915_ (.A_N(net8870),
    .B(net137),
    .X(_04704_));
 sky130_fd_sc_hd__mux2_1 _24916_ (.A0(\pid_q.ki[1] ),
    .A1(_04704_),
    .S(_04702_),
    .X(_04705_));
 sky130_fd_sc_hd__clkbuf_1 _24917_ (.A(_04705_),
    .X(_00746_));
 sky130_fd_sc_hd__and2b_1 _24918_ (.A_N(net8867),
    .B(net138),
    .X(_04706_));
 sky130_fd_sc_hd__mux2_1 _24919_ (.A0(\pid_q.ki[2] ),
    .A1(_04706_),
    .S(net1360),
    .X(_04707_));
 sky130_fd_sc_hd__clkbuf_1 _24920_ (.A(_04707_),
    .X(_00747_));
 sky130_fd_sc_hd__and2b_1 _24921_ (.A_N(net8866),
    .B(net139),
    .X(_04708_));
 sky130_fd_sc_hd__mux2_1 _24922_ (.A0(\pid_q.ki[3] ),
    .A1(_04708_),
    .S(net1362),
    .X(_04709_));
 sky130_fd_sc_hd__clkbuf_1 _24923_ (.A(_04709_),
    .X(_00748_));
 sky130_fd_sc_hd__and2b_1 _24924_ (.A_N(net8868),
    .B(net140),
    .X(_04710_));
 sky130_fd_sc_hd__mux2_1 _24925_ (.A0(\pid_q.ki[4] ),
    .A1(_04710_),
    .S(net1362),
    .X(_04711_));
 sky130_fd_sc_hd__clkbuf_1 _24926_ (.A(_04711_),
    .X(_00749_));
 sky130_fd_sc_hd__and2b_1 _24927_ (.A_N(net8867),
    .B(net141),
    .X(_04712_));
 sky130_fd_sc_hd__mux2_1 _24928_ (.A0(\pid_q.ki[5] ),
    .A1(_04712_),
    .S(net1360),
    .X(_04713_));
 sky130_fd_sc_hd__clkbuf_1 _24929_ (.A(_04713_),
    .X(_00750_));
 sky130_fd_sc_hd__and2b_1 _24930_ (.A_N(net8867),
    .B(net142),
    .X(_04714_));
 sky130_fd_sc_hd__mux2_1 _24931_ (.A0(\pid_q.ki[6] ),
    .A1(_04714_),
    .S(net1361),
    .X(_04715_));
 sky130_fd_sc_hd__clkbuf_1 _24932_ (.A(_04715_),
    .X(_00751_));
 sky130_fd_sc_hd__and2b_1 _24933_ (.A_N(net8868),
    .B(net143),
    .X(_04716_));
 sky130_fd_sc_hd__mux2_1 _24934_ (.A0(\pid_q.ki[7] ),
    .A1(_04716_),
    .S(net1361),
    .X(_04717_));
 sky130_fd_sc_hd__clkbuf_1 _24935_ (.A(_04717_),
    .X(_00752_));
 sky130_fd_sc_hd__and2b_1 _24936_ (.A_N(net8868),
    .B(net144),
    .X(_04718_));
 sky130_fd_sc_hd__mux2_1 _24937_ (.A0(\pid_q.ki[8] ),
    .A1(_04718_),
    .S(net1361),
    .X(_04719_));
 sky130_fd_sc_hd__clkbuf_1 _24938_ (.A(_04719_),
    .X(_00753_));
 sky130_fd_sc_hd__and2b_1 _24939_ (.A_N(net8867),
    .B(net145),
    .X(_04720_));
 sky130_fd_sc_hd__mux2_1 _24940_ (.A0(\pid_q.ki[9] ),
    .A1(_04720_),
    .S(net1360),
    .X(_04721_));
 sky130_fd_sc_hd__clkbuf_1 _24941_ (.A(_04721_),
    .X(_00754_));
 sky130_fd_sc_hd__and2b_1 _24942_ (.A_N(net8866),
    .B(net8882),
    .X(_04722_));
 sky130_fd_sc_hd__mux2_1 _24943_ (.A0(\pid_q.ki[10] ),
    .A1(_04722_),
    .S(net1636),
    .X(_04723_));
 sky130_fd_sc_hd__clkbuf_1 _24944_ (.A(_04723_),
    .X(_00755_));
 sky130_fd_sc_hd__and2b_1 _24945_ (.A_N(net8866),
    .B(net132),
    .X(_04724_));
 sky130_fd_sc_hd__mux2_1 _24946_ (.A0(\pid_q.ki[11] ),
    .A1(_04724_),
    .S(net1636),
    .X(_04725_));
 sky130_fd_sc_hd__clkbuf_1 _24947_ (.A(_04725_),
    .X(_00756_));
 sky130_fd_sc_hd__and2b_1 _24948_ (.A_N(net8870),
    .B(net133),
    .X(_04726_));
 sky130_fd_sc_hd__mux2_1 _24949_ (.A0(\pid_q.ki[12] ),
    .A1(_04726_),
    .S(net1636),
    .X(_04727_));
 sky130_fd_sc_hd__clkbuf_1 _24950_ (.A(_04727_),
    .X(_00757_));
 sky130_fd_sc_hd__and2b_1 _24951_ (.A_N(net8871),
    .B(net8881),
    .X(_04728_));
 sky130_fd_sc_hd__mux2_1 _24952_ (.A0(\pid_q.ki[13] ),
    .A1(_04728_),
    .S(net1637),
    .X(_04729_));
 sky130_fd_sc_hd__clkbuf_1 _24953_ (.A(_04729_),
    .X(_00758_));
 sky130_fd_sc_hd__and2b_1 _24954_ (.A_N(net8871),
    .B(net135),
    .X(_04730_));
 sky130_fd_sc_hd__mux2_1 _24955_ (.A0(\pid_q.ki[14] ),
    .A1(_04730_),
    .S(net1637),
    .X(_04731_));
 sky130_fd_sc_hd__clkbuf_1 _24956_ (.A(_04731_),
    .X(_00759_));
 sky130_fd_sc_hd__and2b_1 _24957_ (.A_N(net8869),
    .B(net136),
    .X(_04732_));
 sky130_fd_sc_hd__mux2_1 _24958_ (.A0(\pid_q.ki[15] ),
    .A1(_04732_),
    .S(_04701_),
    .X(_04733_));
 sky130_fd_sc_hd__clkbuf_1 _24959_ (.A(_04733_),
    .X(_00760_));
 sky130_fd_sc_hd__a2bb2o_1 _24960_ (.A1_N(_04699_),
    .A2_N(net114),
    .B1(net3730),
    .B2(net2011),
    .X(_04734_));
 sky130_fd_sc_hd__buf_1 _24961_ (.A(net1635),
    .X(_04735_));
 sky130_fd_sc_hd__mux2_1 _24962_ (.A0(\pid_q.kp[0] ),
    .A1(_04694_),
    .S(_04735_),
    .X(_04736_));
 sky130_fd_sc_hd__clkbuf_1 _24963_ (.A(_04736_),
    .X(_00761_));
 sky130_fd_sc_hd__mux2_1 _24964_ (.A0(\pid_q.kp[1] ),
    .A1(_04704_),
    .S(_04735_),
    .X(_04737_));
 sky130_fd_sc_hd__clkbuf_1 _24965_ (.A(_04737_),
    .X(_00762_));
 sky130_fd_sc_hd__mux2_1 _24966_ (.A0(\pid_q.kp[2] ),
    .A1(_04706_),
    .S(net1357),
    .X(_04738_));
 sky130_fd_sc_hd__clkbuf_1 _24967_ (.A(_04738_),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _24968_ (.A0(\pid_q.kp[3] ),
    .A1(_04708_),
    .S(net1359),
    .X(_04739_));
 sky130_fd_sc_hd__clkbuf_1 _24969_ (.A(_04739_),
    .X(_00764_));
 sky130_fd_sc_hd__mux2_1 _24970_ (.A0(\pid_q.kp[4] ),
    .A1(_04710_),
    .S(net1359),
    .X(_04740_));
 sky130_fd_sc_hd__clkbuf_1 _24971_ (.A(_04740_),
    .X(_00765_));
 sky130_fd_sc_hd__mux2_1 _24972_ (.A0(\pid_q.kp[5] ),
    .A1(_04712_),
    .S(net1357),
    .X(_04741_));
 sky130_fd_sc_hd__clkbuf_1 _24973_ (.A(_04741_),
    .X(_00766_));
 sky130_fd_sc_hd__mux2_1 _24974_ (.A0(\pid_q.kp[6] ),
    .A1(_04714_),
    .S(net1358),
    .X(_04742_));
 sky130_fd_sc_hd__clkbuf_1 _24975_ (.A(_04742_),
    .X(_00767_));
 sky130_fd_sc_hd__mux2_1 _24976_ (.A0(\pid_q.kp[7] ),
    .A1(_04716_),
    .S(net1358),
    .X(_04743_));
 sky130_fd_sc_hd__clkbuf_1 _24977_ (.A(_04743_),
    .X(_00768_));
 sky130_fd_sc_hd__mux2_1 _24978_ (.A0(\pid_q.kp[8] ),
    .A1(_04718_),
    .S(net1358),
    .X(_04744_));
 sky130_fd_sc_hd__clkbuf_1 _24979_ (.A(_04744_),
    .X(_00769_));
 sky130_fd_sc_hd__mux2_1 _24980_ (.A0(\pid_q.kp[9] ),
    .A1(_04720_),
    .S(net1357),
    .X(_04745_));
 sky130_fd_sc_hd__clkbuf_1 _24981_ (.A(_04745_),
    .X(_00770_));
 sky130_fd_sc_hd__mux2_1 _24982_ (.A0(\pid_q.kp[10] ),
    .A1(_04722_),
    .S(net1634),
    .X(_04746_));
 sky130_fd_sc_hd__clkbuf_1 _24983_ (.A(_04746_),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_1 _24984_ (.A0(\pid_q.kp[11] ),
    .A1(_04724_),
    .S(net1634),
    .X(_04747_));
 sky130_fd_sc_hd__clkbuf_1 _24985_ (.A(_04747_),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _24986_ (.A0(\pid_q.kp[12] ),
    .A1(_04726_),
    .S(net1634),
    .X(_04748_));
 sky130_fd_sc_hd__clkbuf_1 _24987_ (.A(_04748_),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_1 _24988_ (.A0(\pid_q.kp[13] ),
    .A1(_04728_),
    .S(_04734_),
    .X(_04749_));
 sky130_fd_sc_hd__clkbuf_1 _24989_ (.A(_04749_),
    .X(_00774_));
 sky130_fd_sc_hd__mux2_1 _24990_ (.A0(\pid_q.kp[14] ),
    .A1(_04730_),
    .S(net1635),
    .X(_04750_));
 sky130_fd_sc_hd__clkbuf_1 _24991_ (.A(_04750_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _24992_ (.A0(net4475),
    .A1(_04732_),
    .S(_04734_),
    .X(_04751_));
 sky130_fd_sc_hd__clkbuf_1 _24993_ (.A(_04751_),
    .X(_00776_));
 sky130_fd_sc_hd__clkbuf_1 _24994_ (.A(net2147),
    .X(_04752_));
 sky130_fd_sc_hd__nor3b_1 _24995_ (.A(net7483),
    .B(net3270),
    .C_N(net8874),
    .Y(_04753_));
 sky130_fd_sc_hd__xor2_1 _24996_ (.A(\pid_q.out[0] ),
    .B(net5183),
    .X(_04754_));
 sky130_fd_sc_hd__a22o_1 _24997_ (.A1(net7498),
    .A2(net543),
    .B1(_04754_),
    .B2(net7472),
    .X(_04755_));
 sky130_fd_sc_hd__a22o_1 _24998_ (.A1(net9163),
    .A2(net1632),
    .B1(net2395),
    .B2(_04755_),
    .X(_00777_));
 sky130_fd_sc_hd__xor2_1 _24999_ (.A(\pid_q.out[1] ),
    .B(net5181),
    .X(_04756_));
 sky130_fd_sc_hd__a21o_1 _25000_ (.A1(net4474),
    .A2(net5183),
    .B1(_04756_),
    .X(_04757_));
 sky130_fd_sc_hd__nand3_1 _25001_ (.A(net4474),
    .B(net5183),
    .C(_04756_),
    .Y(_04758_));
 sky130_fd_sc_hd__a32o_1 _25002_ (.A1(net7472),
    .A2(_04757_),
    .A3(_04758_),
    .B1(net7498),
    .B2(net538),
    .X(_04759_));
 sky130_fd_sc_hd__a22o_1 _25003_ (.A1(\pid_q.out[1] ),
    .A2(net1631),
    .B1(net2394),
    .B2(_04759_),
    .X(_00778_));
 sky130_fd_sc_hd__or2_1 _25004_ (.A(\pid_q.out[1] ),
    .B(net5181),
    .X(_04760_));
 sky130_fd_sc_hd__a22o_1 _25005_ (.A1(net4474),
    .A2(net5183),
    .B1(\pid_q.out[1] ),
    .B2(net5181),
    .X(_04761_));
 sky130_fd_sc_hd__and2_1 _25006_ (.A(_04760_),
    .B(_04761_),
    .X(_04762_));
 sky130_fd_sc_hd__xor2_1 _25007_ (.A(net4466),
    .B(net5179),
    .X(_04763_));
 sky130_fd_sc_hd__or2_1 _25008_ (.A(_04762_),
    .B(_04763_),
    .X(_04764_));
 sky130_fd_sc_hd__nand2_1 _25009_ (.A(_04762_),
    .B(_04763_),
    .Y(_04765_));
 sky130_fd_sc_hd__a32o_1 _25010_ (.A1(net7472),
    .A2(_04764_),
    .A3(_04765_),
    .B1(net7498),
    .B2(net512),
    .X(_04766_));
 sky130_fd_sc_hd__a22o_1 _25011_ (.A1(net4466),
    .A2(net1631),
    .B1(net2394),
    .B2(_04766_),
    .X(_00779_));
 sky130_fd_sc_hd__a31o_1 _25012_ (.A1(net5179),
    .A2(_04760_),
    .A3(_04761_),
    .B1(net4466),
    .X(_04767_));
 sky130_fd_sc_hd__o21ai_2 _25013_ (.A1(net5179),
    .A2(_04762_),
    .B1(_04767_),
    .Y(_04768_));
 sky130_fd_sc_hd__xnor2_1 _25014_ (.A(net4462),
    .B(\pid_q.curr_int[3] ),
    .Y(_04769_));
 sky130_fd_sc_hd__nand2_1 _25015_ (.A(_04768_),
    .B(_04769_),
    .Y(_04770_));
 sky130_fd_sc_hd__or2_1 _25016_ (.A(_04768_),
    .B(_04769_),
    .X(_04771_));
 sky130_fd_sc_hd__a32o_1 _25017_ (.A1(net7471),
    .A2(_04770_),
    .A3(_04771_),
    .B1(net7497),
    .B2(net467),
    .X(_04772_));
 sky130_fd_sc_hd__a22o_1 _25018_ (.A1(net4462),
    .A2(net1631),
    .B1(net2394),
    .B2(_04772_),
    .X(_00780_));
 sky130_fd_sc_hd__o21ba_1 _25019_ (.A1(_03578_),
    .A2(_04768_),
    .B1_N(net4462),
    .X(_04773_));
 sky130_fd_sc_hd__a21o_1 _25020_ (.A1(_03578_),
    .A2(_04768_),
    .B1(_04773_),
    .X(_04774_));
 sky130_fd_sc_hd__xnor2_1 _25021_ (.A(net4457),
    .B(\pid_q.curr_int[4] ),
    .Y(_04775_));
 sky130_fd_sc_hd__nand2_1 _25022_ (.A(_04774_),
    .B(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__or2_1 _25023_ (.A(_04774_),
    .B(_04775_),
    .X(_04777_));
 sky130_fd_sc_hd__a32o_1 _25024_ (.A1(net7471),
    .A2(_04776_),
    .A3(_04777_),
    .B1(net7497),
    .B2(net462),
    .X(_04778_));
 sky130_fd_sc_hd__a22o_1 _25025_ (.A1(net4457),
    .A2(net1631),
    .B1(net2394),
    .B2(_04778_),
    .X(_00781_));
 sky130_fd_sc_hd__and2_1 _25026_ (.A(net7512),
    .B(net2396),
    .X(_04779_));
 sky130_fd_sc_hd__clkbuf_1 _25027_ (.A(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__o21ba_1 _25028_ (.A1(_03671_),
    .A2(_04774_),
    .B1_N(net4457),
    .X(_04781_));
 sky130_fd_sc_hd__a21o_1 _25029_ (.A1(_03671_),
    .A2(_04774_),
    .B1(_04781_),
    .X(_04782_));
 sky130_fd_sc_hd__xnor2_1 _25030_ (.A(net3739),
    .B(net1157),
    .Y(_04783_));
 sky130_fd_sc_hd__and2_1 _25031_ (.A(net7473),
    .B(net2396),
    .X(_04784_));
 sky130_fd_sc_hd__clkbuf_1 _25032_ (.A(_04784_),
    .X(_04785_));
 sky130_fd_sc_hd__a21o_1 _25033_ (.A1(_04783_),
    .A2(net1628),
    .B1(net2147),
    .X(_04786_));
 sky130_fd_sc_hd__nand2_1 _25034_ (.A(net7473),
    .B(net2396),
    .Y(_04787_));
 sky130_fd_sc_hd__nor3_1 _25035_ (.A(\pid_q.out[5] ),
    .B(_04783_),
    .C(net1995),
    .Y(_04788_));
 sky130_fd_sc_hd__a221o_1 _25036_ (.A1(net405),
    .A2(net1630),
    .B1(_04786_),
    .B2(net9166),
    .C1(_04788_),
    .X(_00782_));
 sky130_fd_sc_hd__o21ba_1 _25037_ (.A1(net3739),
    .A2(net1157),
    .B1_N(\pid_q.out[5] ),
    .X(_04789_));
 sky130_fd_sc_hd__a21o_1 _25038_ (.A1(net3739),
    .A2(net1157),
    .B1(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__xnor2_1 _25039_ (.A(net3738),
    .B(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__a21o_1 _25040_ (.A1(net1628),
    .A2(_04791_),
    .B1(net2147),
    .X(_04792_));
 sky130_fd_sc_hd__nor3_1 _25041_ (.A(\pid_q.out[6] ),
    .B(net1995),
    .C(_04791_),
    .Y(_04793_));
 sky130_fd_sc_hd__a221o_1 _25042_ (.A1(net331),
    .A2(net1630),
    .B1(_04792_),
    .B2(net9174),
    .C1(_04793_),
    .X(_00783_));
 sky130_fd_sc_hd__o21ba_1 _25043_ (.A1(net3738),
    .A2(_04790_),
    .B1_N(\pid_q.out[6] ),
    .X(_04794_));
 sky130_fd_sc_hd__a21o_1 _25044_ (.A1(net3738),
    .A2(_04790_),
    .B1(_04794_),
    .X(_04795_));
 sky130_fd_sc_hd__xnor2_1 _25045_ (.A(\pid_q.out[7] ),
    .B(net5178),
    .Y(_04796_));
 sky130_fd_sc_hd__nand2_1 _25046_ (.A(_04795_),
    .B(_04796_),
    .Y(_04797_));
 sky130_fd_sc_hd__or2_1 _25047_ (.A(_04795_),
    .B(_04796_),
    .X(_04798_));
 sky130_fd_sc_hd__a32o_1 _25048_ (.A1(net7473),
    .A2(_04797_),
    .A3(_04798_),
    .B1(net7512),
    .B2(net329),
    .X(_04799_));
 sky130_fd_sc_hd__a22o_1 _25049_ (.A1(net9229),
    .A2(net1632),
    .B1(net2395),
    .B2(_04799_),
    .X(_00784_));
 sky130_fd_sc_hd__a21bo_1 _25050_ (.A1(_03955_),
    .A2(_04795_),
    .B1_N(\pid_q.out[7] ),
    .X(_04800_));
 sky130_fd_sc_hd__o21a_1 _25051_ (.A1(_03955_),
    .A2(_04795_),
    .B1(_04800_),
    .X(_04801_));
 sky130_fd_sc_hd__xnor2_1 _25052_ (.A(net3737),
    .B(net685),
    .Y(_04802_));
 sky130_fd_sc_hd__a21o_1 _25053_ (.A1(net1628),
    .A2(_04802_),
    .B1(net2147),
    .X(_04803_));
 sky130_fd_sc_hd__nor3_1 _25054_ (.A(\pid_q.out[8] ),
    .B(net1995),
    .C(_04802_),
    .Y(_04804_));
 sky130_fd_sc_hd__a221o_1 _25055_ (.A1(net239),
    .A2(net1630),
    .B1(_04803_),
    .B2(net9173),
    .C1(_04804_),
    .X(_00785_));
 sky130_fd_sc_hd__o21ba_1 _25056_ (.A1(net3737),
    .A2(net685),
    .B1_N(\pid_q.out[8] ),
    .X(_04805_));
 sky130_fd_sc_hd__a21o_1 _25057_ (.A1(net3737),
    .A2(net685),
    .B1(_04805_),
    .X(_04806_));
 sky130_fd_sc_hd__xnor2_1 _25058_ (.A(net3732),
    .B(_04806_),
    .Y(_04807_));
 sky130_fd_sc_hd__a21o_1 _25059_ (.A1(net1628),
    .A2(_04807_),
    .B1(net2147),
    .X(_04808_));
 sky130_fd_sc_hd__nor3_1 _25060_ (.A(net4430),
    .B(net1995),
    .C(_04807_),
    .Y(_04809_));
 sky130_fd_sc_hd__a221o_1 _25061_ (.A1(net266),
    .A2(net1630),
    .B1(_04808_),
    .B2(net4430),
    .C1(_04809_),
    .X(_00786_));
 sky130_fd_sc_hd__o21ba_1 _25062_ (.A1(net3732),
    .A2(_04806_),
    .B1_N(net4430),
    .X(_04810_));
 sky130_fd_sc_hd__a21o_1 _25063_ (.A1(net3732),
    .A2(_04806_),
    .B1(_04810_),
    .X(_04811_));
 sky130_fd_sc_hd__xnor2_1 _25064_ (.A(net3734),
    .B(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__a21o_1 _25065_ (.A1(net1627),
    .A2(_04812_),
    .B1(net2148),
    .X(_04813_));
 sky130_fd_sc_hd__or2_1 _25066_ (.A(net510),
    .B(net238),
    .X(_04814_));
 sky130_fd_sc_hd__nor3_1 _25067_ (.A(net4424),
    .B(net1994),
    .C(_04812_),
    .Y(_04815_));
 sky130_fd_sc_hd__a221o_1 _25068_ (.A1(net4424),
    .A2(_04813_),
    .B1(net193),
    .B2(net1629),
    .C1(_04815_),
    .X(_00787_));
 sky130_fd_sc_hd__a21bo_1 _25069_ (.A1(net3734),
    .A2(_04811_),
    .B1_N(net4424),
    .X(_04816_));
 sky130_fd_sc_hd__o21a_1 _25070_ (.A1(net3734),
    .A2(_04811_),
    .B1(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__xor2_1 _25071_ (.A(net4418),
    .B(net5176),
    .X(_04818_));
 sky130_fd_sc_hd__nand2_1 _25072_ (.A(_04817_),
    .B(_04818_),
    .Y(_04819_));
 sky130_fd_sc_hd__or2_1 _25073_ (.A(_04817_),
    .B(_04818_),
    .X(_04820_));
 sky130_fd_sc_hd__a21oi_1 _25074_ (.A1(_04819_),
    .A2(_04820_),
    .B1(net1994),
    .Y(_04821_));
 sky130_fd_sc_hd__a221o_1 _25075_ (.A1(net4418),
    .A2(net1633),
    .B1(net291),
    .B2(net1629),
    .C1(_04821_),
    .X(_00788_));
 sky130_fd_sc_hd__inv_2 _25076_ (.A(net5176),
    .Y(_04822_));
 sky130_fd_sc_hd__o21ba_1 _25077_ (.A1(_04822_),
    .A2(_04817_),
    .B1_N(net4418),
    .X(_04823_));
 sky130_fd_sc_hd__a21oi_2 _25078_ (.A1(_04822_),
    .A2(_04817_),
    .B1(_04823_),
    .Y(_04824_));
 sky130_fd_sc_hd__xnor2_1 _25079_ (.A(net4406),
    .B(net5174),
    .Y(_04825_));
 sky130_fd_sc_hd__or2_1 _25080_ (.A(_04824_),
    .B(_04825_),
    .X(_04826_));
 sky130_fd_sc_hd__nand2_1 _25081_ (.A(_04824_),
    .B(_04825_),
    .Y(_04827_));
 sky130_fd_sc_hd__a21oi_1 _25082_ (.A1(_04826_),
    .A2(_04827_),
    .B1(net1994),
    .Y(_04828_));
 sky130_fd_sc_hd__a221o_1 _25083_ (.A1(net4406),
    .A2(net1633),
    .B1(net235),
    .B2(net1629),
    .C1(_04828_),
    .X(_00789_));
 sky130_fd_sc_hd__nand2_1 _25084_ (.A(net7499),
    .B(net2396),
    .Y(_04829_));
 sky130_fd_sc_hd__a21o_1 _25085_ (.A1(net5174),
    .A2(_04824_),
    .B1(net4406),
    .X(_04830_));
 sky130_fd_sc_hd__o21a_1 _25086_ (.A1(net5174),
    .A2(_04824_),
    .B1(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__xnor2_1 _25087_ (.A(net5172),
    .B(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__a21o_1 _25088_ (.A1(net1627),
    .A2(_04832_),
    .B1(net1633),
    .X(_04833_));
 sky130_fd_sc_hd__nand2_1 _25089_ (.A(net4401),
    .B(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__or3_1 _25090_ (.A(net4401),
    .B(_04787_),
    .C(_04832_),
    .X(_04835_));
 sky130_fd_sc_hd__o211ai_1 _25091_ (.A1(net198),
    .A2(_04829_),
    .B1(_04834_),
    .C1(_04835_),
    .Y(_00790_));
 sky130_fd_sc_hd__inv_2 _25092_ (.A(net5171),
    .Y(_04836_));
 sky130_fd_sc_hd__a221o_1 _25093_ (.A1(net4401),
    .A2(net5172),
    .B1(_04824_),
    .B2(net5174),
    .C1(net4406),
    .X(_04837_));
 sky130_fd_sc_hd__a211o_1 _25094_ (.A1(net4401),
    .A2(net5172),
    .B1(_04824_),
    .C1(net5174),
    .X(_04838_));
 sky130_fd_sc_hd__o211ai_2 _25095_ (.A1(net4401),
    .A2(net5172),
    .B1(_04837_),
    .C1(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__xnor2_1 _25096_ (.A(_04836_),
    .B(_04839_),
    .Y(_04840_));
 sky130_fd_sc_hd__inv_2 _25097_ (.A(net4400),
    .Y(_04841_));
 sky130_fd_sc_hd__a211o_1 _25098_ (.A1(net1627),
    .A2(_04840_),
    .B1(_04841_),
    .C1(net2148),
    .X(_04842_));
 sky130_fd_sc_hd__o21ai_1 _25099_ (.A1(net1994),
    .A2(_04840_),
    .B1(_04841_),
    .Y(_04843_));
 sky130_fd_sc_hd__a22o_1 _25100_ (.A1(net232),
    .A2(net1629),
    .B1(_04842_),
    .B2(_04843_),
    .X(_00791_));
 sky130_fd_sc_hd__a21bo_1 _25101_ (.A1(_04836_),
    .A2(_04839_),
    .B1_N(net4400),
    .X(_04844_));
 sky130_fd_sc_hd__o21a_1 _25102_ (.A1(_04836_),
    .A2(_04839_),
    .B1(_04844_),
    .X(_04845_));
 sky130_fd_sc_hd__xor2_1 _25103_ (.A(net4393),
    .B(net5169),
    .X(_04846_));
 sky130_fd_sc_hd__xnor2_1 _25104_ (.A(_04845_),
    .B(_04846_),
    .Y(_04847_));
 sky130_fd_sc_hd__nor2_1 _25105_ (.A(net196),
    .B(_04829_),
    .Y(_04848_));
 sky130_fd_sc_hd__a221o_1 _25106_ (.A1(net4393),
    .A2(net1633),
    .B1(net1627),
    .B2(_04847_),
    .C1(_04848_),
    .X(_00792_));
 sky130_fd_sc_hd__a21oi_2 _25107_ (.A1(net4297),
    .A2(net9248),
    .B1(net4308),
    .Y(_04849_));
 sky130_fd_sc_hd__buf_1 _25108_ (.A(net3033),
    .X(_04850_));
 sky130_fd_sc_hd__and4_1 _25109_ (.A(net8902),
    .B(net4300),
    .C(net4332),
    .D(net3762),
    .X(_04851_));
 sky130_fd_sc_hd__clkbuf_2 _25110_ (.A(_04851_),
    .X(_04852_));
 sky130_fd_sc_hd__buf_1 _25111_ (.A(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__a22o_1 _25112_ (.A1(net4392),
    .A2(net2392),
    .B1(net1992),
    .B2(net9206),
    .X(_00793_));
 sky130_fd_sc_hd__a22o_1 _25113_ (.A1(\pid_d.prev_int[1] ),
    .A2(net2392),
    .B1(net1992),
    .B2(net5985),
    .X(_00794_));
 sky130_fd_sc_hd__a22o_1 _25114_ (.A1(\pid_d.prev_int[2] ),
    .A2(net2392),
    .B1(net1992),
    .B2(net9079),
    .X(_00795_));
 sky130_fd_sc_hd__a22o_1 _25115_ (.A1(\pid_d.prev_int[3] ),
    .A2(net2392),
    .B1(net1992),
    .B2(\pid_d.curr_int[3] ),
    .X(_00796_));
 sky130_fd_sc_hd__a22o_1 _25116_ (.A1(net9209),
    .A2(net2393),
    .B1(net1993),
    .B2(\pid_d.curr_int[4] ),
    .X(_00797_));
 sky130_fd_sc_hd__a22o_1 _25117_ (.A1(net9236),
    .A2(net2393),
    .B1(net1993),
    .B2(\pid_d.curr_int[5] ),
    .X(_00798_));
 sky130_fd_sc_hd__a22o_1 _25118_ (.A1(\pid_d.prev_int[6] ),
    .A2(net2393),
    .B1(net1993),
    .B2(net9196),
    .X(_00799_));
 sky130_fd_sc_hd__a22o_1 _25119_ (.A1(net9215),
    .A2(net2393),
    .B1(net1993),
    .B2(net5978),
    .X(_00800_));
 sky130_fd_sc_hd__a22o_1 _25120_ (.A1(net9217),
    .A2(_04850_),
    .B1(_04853_),
    .B2(net5977),
    .X(_00801_));
 sky130_fd_sc_hd__a22o_1 _25121_ (.A1(net9205),
    .A2(_04850_),
    .B1(_04853_),
    .B2(net5976),
    .X(_00802_));
 sky130_fd_sc_hd__a22o_1 _25122_ (.A1(\pid_d.prev_int[10] ),
    .A2(net3033),
    .B1(_04852_),
    .B2(net9169),
    .X(_00803_));
 sky130_fd_sc_hd__a22o_1 _25123_ (.A1(net9224),
    .A2(net3033),
    .B1(_04852_),
    .B2(\pid_d.curr_int[11] ),
    .X(_00804_));
 sky130_fd_sc_hd__a22o_1 _25124_ (.A1(net4391),
    .A2(_04849_),
    .B1(net2391),
    .B2(net5975),
    .X(_00805_));
 sky130_fd_sc_hd__a22o_1 _25125_ (.A1(net9109),
    .A2(_04849_),
    .B1(net2391),
    .B2(\pid_d.curr_int[13] ),
    .X(_00806_));
 sky130_fd_sc_hd__a22o_1 _25126_ (.A1(\pid_d.prev_int[14] ),
    .A2(_04849_),
    .B1(net2391),
    .B2(\pid_d.curr_int[14] ),
    .X(_00807_));
 sky130_fd_sc_hd__a22o_1 _25127_ (.A1(net9134),
    .A2(_04849_),
    .B1(net2391),
    .B2(net5974),
    .X(_00808_));
 sky130_fd_sc_hd__dfrtp_1 _25128_ (.CLK(clknet_leaf_51_clk),
    .D(_00017_),
    .RESET_B(net8809),
    .Q(\svm0.tC[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25129_ (.CLK(clknet_leaf_52_clk),
    .D(_00018_),
    .RESET_B(net8805),
    .Q(\svm0.tC[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25130_ (.CLK(clknet_leaf_52_clk),
    .D(_00019_),
    .RESET_B(net8805),
    .Q(\svm0.tC[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25131_ (.CLK(clknet_leaf_52_clk),
    .D(_00020_),
    .RESET_B(net8805),
    .Q(\svm0.tC[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25132_ (.CLK(clknet_leaf_52_clk),
    .D(_00021_),
    .RESET_B(net8803),
    .Q(\svm0.tC[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25133_ (.CLK(clknet_leaf_52_clk),
    .D(_00022_),
    .RESET_B(net8803),
    .Q(\svm0.tC[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25134_ (.CLK(clknet_leaf_52_clk),
    .D(_00023_),
    .RESET_B(net8803),
    .Q(\svm0.tC[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25135_ (.CLK(clknet_leaf_52_clk),
    .D(_00024_),
    .RESET_B(net8806),
    .Q(\svm0.tC[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25136_ (.CLK(clknet_leaf_51_clk),
    .D(_00025_),
    .RESET_B(net8809),
    .Q(\svm0.tC[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25137_ (.CLK(clknet_leaf_51_clk),
    .D(_00026_),
    .RESET_B(net8809),
    .Q(\svm0.tC[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25138_ (.CLK(clknet_4_14__leaf_clk),
    .D(_00027_),
    .RESET_B(net8832),
    .Q(\svm0.tC[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25139_ (.CLK(clknet_leaf_51_clk),
    .D(_00028_),
    .RESET_B(net8810),
    .Q(\svm0.tC[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25140_ (.CLK(clknet_leaf_50_clk),
    .D(_00029_),
    .RESET_B(net8757),
    .Q(\svm0.tC[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25141_ (.CLK(clknet_leaf_50_clk),
    .D(_00030_),
    .RESET_B(net8757),
    .Q(\svm0.tC[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25142_ (.CLK(clknet_leaf_50_clk),
    .D(_00031_),
    .RESET_B(net8757),
    .Q(\svm0.tC[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25143_ (.CLK(clknet_leaf_48_clk),
    .D(_00032_),
    .RESET_B(net8762),
    .Q(\svm0.tC[15] ));
 sky130_fd_sc_hd__dfstp_1 _25144_ (.CLK(clknet_leaf_65_clk),
    .D(_00033_),
    .SET_B(net8655),
    .Q(net152));
 sky130_fd_sc_hd__dfrtp_1 _25145_ (.CLK(clknet_leaf_104_clk),
    .D(_00034_),
    .RESET_B(net8363),
    .Q(\cordic0.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25146_ (.CLK(clknet_leaf_41_clk),
    .D(_00035_),
    .RESET_B(net8767),
    .Q(\pid_q.target[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25147_ (.CLK(clknet_leaf_41_clk),
    .D(_00036_),
    .RESET_B(net8767),
    .Q(\pid_q.target[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25148_ (.CLK(clknet_leaf_41_clk),
    .D(_00037_),
    .RESET_B(net8767),
    .Q(\pid_q.target[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25149_ (.CLK(clknet_leaf_44_clk),
    .D(_00038_),
    .RESET_B(net8781),
    .Q(\pid_q.target[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25150_ (.CLK(clknet_leaf_41_clk),
    .D(_00039_),
    .RESET_B(net8767),
    .Q(\pid_q.target[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25151_ (.CLK(clknet_leaf_44_clk),
    .D(_00040_),
    .RESET_B(net8781),
    .Q(\pid_q.target[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25152_ (.CLK(clknet_leaf_41_clk),
    .D(_00041_),
    .RESET_B(net8767),
    .Q(\pid_q.target[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25153_ (.CLK(clknet_leaf_41_clk),
    .D(_00042_),
    .RESET_B(net8767),
    .Q(\pid_q.target[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25154_ (.CLK(clknet_leaf_41_clk),
    .D(_00043_),
    .RESET_B(net8767),
    .Q(\pid_q.target[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25155_ (.CLK(clknet_leaf_44_clk),
    .D(_00044_),
    .RESET_B(net8781),
    .Q(\pid_q.target[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25156_ (.CLK(clknet_leaf_44_clk),
    .D(_00045_),
    .RESET_B(net8781),
    .Q(\pid_q.target[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25157_ (.CLK(clknet_leaf_54_clk),
    .D(_00046_),
    .RESET_B(net8727),
    .Q(\pid_q.target[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25158_ (.CLK(clknet_leaf_54_clk),
    .D(_00047_),
    .RESET_B(net8727),
    .Q(\pid_q.target[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25159_ (.CLK(clknet_leaf_45_clk),
    .D(_00048_),
    .RESET_B(net8781),
    .Q(\pid_q.target[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25160_ (.CLK(clknet_leaf_44_clk),
    .D(_00049_),
    .RESET_B(net8785),
    .Q(\pid_q.target[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25161_ (.CLK(clknet_leaf_45_clk),
    .D(_00050_),
    .RESET_B(net8785),
    .Q(\pid_q.target[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25162_ (.CLK(clknet_leaf_54_clk),
    .D(_00051_),
    .RESET_B(net8730),
    .Q(\svm0.periodTop[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25163_ (.CLK(clknet_leaf_54_clk),
    .D(_00052_),
    .RESET_B(net8730),
    .Q(\svm0.periodTop[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25164_ (.CLK(clknet_leaf_54_clk),
    .D(_00053_),
    .RESET_B(net8730),
    .Q(\svm0.periodTop[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25165_ (.CLK(clknet_leaf_54_clk),
    .D(_00054_),
    .RESET_B(net8730),
    .Q(\svm0.periodTop[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25166_ (.CLK(clknet_leaf_55_clk),
    .D(_00055_),
    .RESET_B(net8728),
    .Q(\svm0.periodTop[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25167_ (.CLK(clknet_leaf_55_clk),
    .D(_00056_),
    .RESET_B(net8728),
    .Q(\svm0.periodTop[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25168_ (.CLK(clknet_leaf_55_clk),
    .D(_00057_),
    .RESET_B(net8728),
    .Q(\svm0.periodTop[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25169_ (.CLK(clknet_leaf_54_clk),
    .D(_00058_),
    .RESET_B(net8729),
    .Q(\svm0.periodTop[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25170_ (.CLK(clknet_leaf_54_clk),
    .D(_00059_),
    .RESET_B(net8730),
    .Q(\svm0.periodTop[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25171_ (.CLK(clknet_leaf_54_clk),
    .D(_00060_),
    .RESET_B(net8729),
    .Q(\svm0.periodTop[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25172_ (.CLK(clknet_leaf_55_clk),
    .D(_00061_),
    .RESET_B(net8728),
    .Q(\svm0.periodTop[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25173_ (.CLK(clknet_leaf_54_clk),
    .D(_00062_),
    .RESET_B(net8730),
    .Q(\svm0.periodTop[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25174_ (.CLK(clknet_leaf_54_clk),
    .D(_00063_),
    .RESET_B(net8730),
    .Q(\svm0.periodTop[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25175_ (.CLK(clknet_leaf_54_clk),
    .D(_00064_),
    .RESET_B(net8730),
    .Q(\svm0.periodTop[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25176_ (.CLK(clknet_leaf_54_clk),
    .D(_00065_),
    .RESET_B(net8729),
    .Q(\svm0.periodTop[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25177_ (.CLK(clknet_leaf_55_clk),
    .D(_00066_),
    .RESET_B(net8728),
    .Q(\svm0.periodTop[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25178_ (.CLK(clknet_leaf_72_clk),
    .D(_00067_),
    .RESET_B(net8469),
    .Q(\matmul0.a_in[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25179_ (.CLK(clknet_leaf_95_clk),
    .D(_00068_),
    .RESET_B(net8448),
    .Q(\matmul0.a_in[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25180_ (.CLK(clknet_leaf_68_clk),
    .D(_00069_),
    .RESET_B(net8452),
    .Q(\matmul0.a_in[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25181_ (.CLK(clknet_leaf_70_clk),
    .D(_00070_),
    .RESET_B(net8452),
    .Q(\matmul0.a_in[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25182_ (.CLK(clknet_leaf_68_clk),
    .D(_00071_),
    .RESET_B(net8450),
    .Q(\matmul0.a_in[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25183_ (.CLK(clknet_leaf_67_clk),
    .D(_00072_),
    .RESET_B(net8450),
    .Q(\matmul0.a_in[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25184_ (.CLK(clknet_leaf_72_clk),
    .D(_00073_),
    .RESET_B(net8470),
    .Q(\matmul0.a_in[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25185_ (.CLK(clknet_leaf_69_clk),
    .D(_00074_),
    .RESET_B(net8468),
    .Q(\matmul0.a_in[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25186_ (.CLK(clknet_leaf_72_clk),
    .D(_00075_),
    .RESET_B(net8662),
    .Q(\matmul0.a_in[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25187_ (.CLK(clknet_leaf_63_clk),
    .D(_00076_),
    .RESET_B(net8667),
    .Q(\matmul0.a_in[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25188_ (.CLK(clknet_leaf_62_clk),
    .D(_00077_),
    .RESET_B(net8671),
    .Q(\matmul0.a_in[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25189_ (.CLK(clknet_leaf_58_clk),
    .D(_00078_),
    .RESET_B(net8720),
    .Q(\matmul0.a_in[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25190_ (.CLK(clknet_leaf_57_clk),
    .D(_00079_),
    .RESET_B(net8711),
    .Q(\matmul0.a_in[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25191_ (.CLK(clknet_leaf_61_clk),
    .D(_00080_),
    .RESET_B(net8721),
    .Q(\matmul0.a_in[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25192_ (.CLK(clknet_leaf_58_clk),
    .D(_00081_),
    .RESET_B(net8721),
    .Q(\matmul0.a_in[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25193_ (.CLK(clknet_leaf_58_clk),
    .D(_00082_),
    .RESET_B(net8721),
    .Q(\matmul0.a_in[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25194_ (.CLK(clknet_leaf_63_clk),
    .D(_00083_),
    .RESET_B(net8665),
    .Q(\matmul0.b_in[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25195_ (.CLK(clknet_leaf_62_clk),
    .D(_00084_),
    .RESET_B(net8708),
    .Q(\matmul0.b_in[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25196_ (.CLK(clknet_leaf_63_clk),
    .D(_00085_),
    .RESET_B(net8665),
    .Q(\matmul0.b_in[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25197_ (.CLK(clknet_leaf_63_clk),
    .D(_00086_),
    .RESET_B(net8665),
    .Q(\matmul0.b_in[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25198_ (.CLK(clknet_leaf_73_clk),
    .D(_00087_),
    .RESET_B(net8474),
    .Q(\matmul0.b_in[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25199_ (.CLK(clknet_leaf_62_clk),
    .D(_00088_),
    .RESET_B(net8666),
    .Q(\matmul0.b_in[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25200_ (.CLK(clknet_leaf_58_clk),
    .D(_00089_),
    .RESET_B(net8710),
    .Q(\matmul0.b_in[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25201_ (.CLK(clknet_leaf_82_clk),
    .D(_00090_),
    .RESET_B(net8496),
    .Q(\matmul0.b_in[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25202_ (.CLK(clknet_leaf_81_clk),
    .D(_00091_),
    .RESET_B(net8495),
    .Q(\matmul0.b_in[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25203_ (.CLK(clknet_leaf_57_clk),
    .D(_00092_),
    .RESET_B(net8715),
    .Q(\matmul0.b_in[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25204_ (.CLK(clknet_leaf_57_clk),
    .D(_00093_),
    .RESET_B(net8715),
    .Q(\matmul0.b_in[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25205_ (.CLK(clknet_leaf_57_clk),
    .D(_00094_),
    .RESET_B(net8715),
    .Q(\matmul0.b_in[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25206_ (.CLK(clknet_leaf_82_clk),
    .D(_00095_),
    .RESET_B(net8709),
    .Q(\matmul0.b_in[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25207_ (.CLK(clknet_leaf_62_clk),
    .D(_00096_),
    .RESET_B(net8666),
    .Q(\matmul0.b_in[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25208_ (.CLK(clknet_leaf_61_clk),
    .D(_00097_),
    .RESET_B(net8671),
    .Q(\matmul0.b_in[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25209_ (.CLK(clknet_leaf_62_clk),
    .D(_00098_),
    .RESET_B(net8672),
    .Q(\matmul0.b_in[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25210_ (.CLK(clknet_leaf_64_clk),
    .D(_00099_),
    .RESET_B(net8670),
    .Q(\matmul0.op_in[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25211_ (.CLK(clknet_leaf_64_clk),
    .D(_00100_),
    .RESET_B(net8661),
    .Q(\matmul0.op_in[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25212_ (.CLK(clknet_leaf_61_clk),
    .D(_00101_),
    .RESET_B(net8717),
    .Q(\svm0.vC[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25213_ (.CLK(clknet_leaf_61_clk),
    .D(_00102_),
    .RESET_B(net8717),
    .Q(\svm0.vC[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25214_ (.CLK(clknet_leaf_61_clk),
    .D(_00103_),
    .RESET_B(net8717),
    .Q(\svm0.vC[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25215_ (.CLK(clknet_leaf_61_clk),
    .D(_00104_),
    .RESET_B(net8688),
    .Q(\svm0.vC[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25216_ (.CLK(clknet_leaf_59_clk),
    .D(_00105_),
    .RESET_B(net8732),
    .Q(\svm0.vC[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25217_ (.CLK(clknet_leaf_59_clk),
    .D(_00106_),
    .RESET_B(net8688),
    .Q(\svm0.vC[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25218_ (.CLK(clknet_leaf_59_clk),
    .D(_00107_),
    .RESET_B(net8689),
    .Q(\svm0.vC[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25219_ (.CLK(clknet_leaf_59_clk),
    .D(_00108_),
    .RESET_B(net8688),
    .Q(\svm0.vC[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25220_ (.CLK(clknet_leaf_59_clk),
    .D(_00109_),
    .RESET_B(net8693),
    .Q(\svm0.vC[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25221_ (.CLK(clknet_leaf_60_clk),
    .D(_00110_),
    .RESET_B(net8669),
    .Q(\svm0.vC[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25222_ (.CLK(clknet_leaf_59_clk),
    .D(_00111_),
    .RESET_B(net8693),
    .Q(\svm0.vC[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25223_ (.CLK(clknet_leaf_60_clk),
    .D(_00112_),
    .RESET_B(net8690),
    .Q(\svm0.vC[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25224_ (.CLK(clknet_leaf_59_clk),
    .D(_00113_),
    .RESET_B(net8693),
    .Q(\svm0.vC[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25225_ (.CLK(clknet_leaf_59_clk),
    .D(_00114_),
    .RESET_B(net8694),
    .Q(\svm0.vC[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25226_ (.CLK(clknet_leaf_59_clk),
    .D(_00115_),
    .RESET_B(net8694),
    .Q(\svm0.vC[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25227_ (.CLK(clknet_leaf_59_clk),
    .D(_00116_),
    .RESET_B(net8694),
    .Q(\svm0.vC[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25228_ (.CLK(clknet_leaf_66_clk),
    .D(_00117_),
    .RESET_B(net8647),
    .Q(cordic_done));
 sky130_fd_sc_hd__dfrtp_1 _25229_ (.CLK(clknet_leaf_66_clk),
    .D(_00118_),
    .RESET_B(net8647),
    .Q(clarke_done));
 sky130_fd_sc_hd__dfrtp_1 _25230_ (.CLK(clknet_leaf_65_clk),
    .D(_00119_),
    .RESET_B(net8655),
    .Q(\cordic0.in_valid ));
 sky130_fd_sc_hd__dfrtp_1 _25231_ (.CLK(clknet_leaf_64_clk),
    .D(_00120_),
    .RESET_B(net8661),
    .Q(\matmul0.start ));
 sky130_fd_sc_hd__dfrtp_1 _25232_ (.CLK(clknet_leaf_65_clk),
    .D(_00121_),
    .RESET_B(net8655),
    .Q(\pid_d.iterate_enable ));
 sky130_fd_sc_hd__dfstp_1 _25233_ (.CLK(clknet_leaf_23_clk),
    .D(_00016_),
    .SET_B(net8587),
    .Q(\pid_q.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25234_ (.CLK(clknet_leaf_23_clk),
    .D(_00007_),
    .RESET_B(net8582),
    .Q(\pid_q.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25235_ (.CLK(clknet_leaf_17_clk),
    .D(net3007),
    .RESET_B(net8631),
    .Q(\pid_q.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25236_ (.CLK(clknet_leaf_23_clk),
    .D(_00009_),
    .RESET_B(net8582),
    .Q(\pid_q.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25237_ (.CLK(clknet_leaf_23_clk),
    .D(_00010_),
    .RESET_B(net8582),
    .Q(\pid_q.state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25238_ (.CLK(clknet_leaf_32_clk),
    .D(net2384),
    .RESET_B(net8683),
    .Q(\pid_q.state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25239_ (.CLK(clknet_leaf_68_clk),
    .D(_00122_),
    .RESET_B(net8454),
    .Q(\matmul0.op[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25240_ (.CLK(clknet_leaf_69_clk),
    .D(_00123_),
    .RESET_B(net8468),
    .Q(\matmul0.op[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25241_ (.CLK(clknet_leaf_89_clk),
    .D(_00124_),
    .RESET_B(net8421),
    .Q(\matmul0.matmul_stage_inst.a[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25242_ (.CLK(clknet_leaf_86_clk),
    .D(_00125_),
    .RESET_B(net8531),
    .Q(\matmul0.matmul_stage_inst.a[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25243_ (.CLK(clknet_leaf_87_clk),
    .D(_00126_),
    .RESET_B(net8442),
    .Q(\matmul0.matmul_stage_inst.a[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25244_ (.CLK(clknet_leaf_89_clk),
    .D(_00127_),
    .RESET_B(net8443),
    .Q(\matmul0.matmul_stage_inst.a[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25245_ (.CLK(clknet_leaf_87_clk),
    .D(_00128_),
    .RESET_B(net8436),
    .Q(\matmul0.matmul_stage_inst.a[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25246_ (.CLK(clknet_leaf_88_clk),
    .D(_00129_),
    .RESET_B(net8443),
    .Q(\matmul0.matmul_stage_inst.a[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25247_ (.CLK(clknet_leaf_87_clk),
    .D(_00130_),
    .RESET_B(net8436),
    .Q(\matmul0.matmul_stage_inst.a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25248_ (.CLK(clknet_leaf_87_clk),
    .D(_00131_),
    .RESET_B(net8436),
    .Q(\matmul0.matmul_stage_inst.a[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25249_ (.CLK(clknet_leaf_87_clk),
    .D(_00132_),
    .RESET_B(net8442),
    .Q(\matmul0.matmul_stage_inst.a[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25250_ (.CLK(clknet_leaf_87_clk),
    .D(_00133_),
    .RESET_B(net8442),
    .Q(\matmul0.matmul_stage_inst.a[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25251_ (.CLK(clknet_leaf_88_clk),
    .D(_00134_),
    .RESET_B(net8431),
    .Q(\matmul0.matmul_stage_inst.a[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25252_ (.CLK(clknet_leaf_88_clk),
    .D(_00135_),
    .RESET_B(net8430),
    .Q(\matmul0.matmul_stage_inst.a[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25253_ (.CLK(clknet_leaf_88_clk),
    .D(_00136_),
    .RESET_B(net8431),
    .Q(\matmul0.matmul_stage_inst.a[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25254_ (.CLK(clknet_leaf_88_clk),
    .D(_00137_),
    .RESET_B(net8430),
    .Q(\matmul0.matmul_stage_inst.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25255_ (.CLK(clknet_leaf_77_clk),
    .D(_00138_),
    .RESET_B(net8437),
    .Q(\matmul0.matmul_stage_inst.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25256_ (.CLK(clknet_leaf_71_clk),
    .D(_00139_),
    .RESET_B(net8457),
    .Q(\matmul0.matmul_stage_inst.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25257_ (.CLK(clknet_leaf_70_clk),
    .D(_00140_),
    .RESET_B(net8457),
    .Q(\matmul0.matmul_stage_inst.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25258_ (.CLK(clknet_leaf_71_clk),
    .D(_00141_),
    .RESET_B(net8458),
    .Q(\matmul0.matmul_stage_inst.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25259_ (.CLK(clknet_leaf_71_clk),
    .D(_00142_),
    .RESET_B(net8457),
    .Q(\matmul0.matmul_stage_inst.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25260_ (.CLK(clknet_leaf_76_clk),
    .D(_00143_),
    .RESET_B(net8458),
    .Q(\matmul0.matmul_stage_inst.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25261_ (.CLK(clknet_leaf_75_clk),
    .D(_00144_),
    .RESET_B(net8458),
    .Q(\matmul0.matmul_stage_inst.b[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25262_ (.CLK(clknet_leaf_76_clk),
    .D(_00145_),
    .RESET_B(net8458),
    .Q(\matmul0.matmul_stage_inst.b[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25263_ (.CLK(clknet_leaf_77_clk),
    .D(_00146_),
    .RESET_B(net8437),
    .Q(\matmul0.matmul_stage_inst.b[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25264_ (.CLK(clknet_leaf_88_clk),
    .D(_00147_),
    .RESET_B(net8435),
    .Q(\matmul0.matmul_stage_inst.b[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25265_ (.CLK(clknet_leaf_88_clk),
    .D(_00148_),
    .RESET_B(net8435),
    .Q(\matmul0.matmul_stage_inst.b[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25266_ (.CLK(clknet_leaf_88_clk),
    .D(_00149_),
    .RESET_B(net8430),
    .Q(\matmul0.matmul_stage_inst.b[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25267_ (.CLK(clknet_leaf_77_clk),
    .D(_00150_),
    .RESET_B(net8440),
    .Q(\matmul0.matmul_stage_inst.b[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25268_ (.CLK(clknet_leaf_77_clk),
    .D(_00151_),
    .RESET_B(net8437),
    .Q(\matmul0.matmul_stage_inst.b[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25269_ (.CLK(clknet_leaf_88_clk),
    .D(_00152_),
    .RESET_B(net8421),
    .Q(\matmul0.matmul_stage_inst.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25270_ (.CLK(clknet_leaf_92_clk),
    .D(_00153_),
    .RESET_B(net8433),
    .Q(\matmul0.matmul_stage_inst.c[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25271_ (.CLK(clknet_leaf_88_clk),
    .D(_00154_),
    .RESET_B(net8438),
    .Q(\matmul0.matmul_stage_inst.c[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25272_ (.CLK(clknet_leaf_93_clk),
    .D(_00155_),
    .RESET_B(net8446),
    .Q(\matmul0.matmul_stage_inst.c[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25273_ (.CLK(clknet_leaf_93_clk),
    .D(_00156_),
    .RESET_B(net8449),
    .Q(\matmul0.matmul_stage_inst.c[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25274_ (.CLK(clknet_leaf_76_clk),
    .D(_00157_),
    .RESET_B(net8458),
    .Q(\matmul0.matmul_stage_inst.c[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25275_ (.CLK(clknet_leaf_93_clk),
    .D(_00158_),
    .RESET_B(net8447),
    .Q(\matmul0.matmul_stage_inst.c[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25276_ (.CLK(clknet_leaf_77_clk),
    .D(_00159_),
    .RESET_B(net8457),
    .Q(\matmul0.matmul_stage_inst.c[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25277_ (.CLK(clknet_leaf_71_clk),
    .D(_00160_),
    .RESET_B(net8457),
    .Q(\matmul0.matmul_stage_inst.c[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25278_ (.CLK(clknet_leaf_70_clk),
    .D(_00161_),
    .RESET_B(net8447),
    .Q(\matmul0.matmul_stage_inst.c[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25279_ (.CLK(clknet_leaf_92_clk),
    .D(_00162_),
    .RESET_B(net8434),
    .Q(\matmul0.matmul_stage_inst.c[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25280_ (.CLK(clknet_leaf_92_clk),
    .D(_00163_),
    .RESET_B(net8434),
    .Q(\matmul0.matmul_stage_inst.c[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25281_ (.CLK(clknet_leaf_92_clk),
    .D(_00164_),
    .RESET_B(net8428),
    .Q(\matmul0.matmul_stage_inst.c[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25282_ (.CLK(clknet_leaf_92_clk),
    .D(_00165_),
    .RESET_B(net8429),
    .Q(\matmul0.matmul_stage_inst.c[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25283_ (.CLK(clknet_leaf_77_clk),
    .D(_00166_),
    .RESET_B(net8440),
    .Q(\matmul0.matmul_stage_inst.c[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25284_ (.CLK(clknet_leaf_77_clk),
    .D(_00167_),
    .RESET_B(net8440),
    .Q(\matmul0.matmul_stage_inst.c[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25285_ (.CLK(clknet_leaf_89_clk),
    .D(_00168_),
    .RESET_B(net8421),
    .Q(\matmul0.matmul_stage_inst.d[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25286_ (.CLK(clknet_leaf_89_clk),
    .D(_00169_),
    .RESET_B(net8443),
    .Q(\matmul0.matmul_stage_inst.d[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25287_ (.CLK(clknet_leaf_88_clk),
    .D(_00170_),
    .RESET_B(net8444),
    .Q(\matmul0.matmul_stage_inst.d[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25288_ (.CLK(clknet_leaf_89_clk),
    .D(_00171_),
    .RESET_B(net8422),
    .Q(\matmul0.matmul_stage_inst.a[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25289_ (.CLK(clknet_leaf_89_clk),
    .D(_00172_),
    .RESET_B(net8422),
    .Q(\matmul0.matmul_stage_inst.d[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25290_ (.CLK(clknet_leaf_77_clk),
    .D(_00173_),
    .RESET_B(net8436),
    .Q(\matmul0.matmul_stage_inst.d[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25291_ (.CLK(clknet_leaf_88_clk),
    .D(_00174_),
    .RESET_B(net8420),
    .Q(\matmul0.matmul_stage_inst.d[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25292_ (.CLK(clknet_leaf_77_clk),
    .D(_00175_),
    .RESET_B(net8438),
    .Q(\matmul0.matmul_stage_inst.d[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25293_ (.CLK(clknet_leaf_88_clk),
    .D(_00176_),
    .RESET_B(net8435),
    .Q(\matmul0.matmul_stage_inst.d[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25294_ (.CLK(clknet_leaf_88_clk),
    .D(_00177_),
    .RESET_B(net8431),
    .Q(\matmul0.matmul_stage_inst.d[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25295_ (.CLK(clknet_leaf_89_clk),
    .D(_00178_),
    .RESET_B(net8420),
    .Q(\matmul0.matmul_stage_inst.d[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25296_ (.CLK(clknet_leaf_92_clk),
    .D(_00179_),
    .RESET_B(net8429),
    .Q(\matmul0.matmul_stage_inst.d[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25297_ (.CLK(clknet_leaf_92_clk),
    .D(_00180_),
    .RESET_B(net8429),
    .Q(\matmul0.matmul_stage_inst.d[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25298_ (.CLK(clknet_leaf_88_clk),
    .D(_00181_),
    .RESET_B(net8431),
    .Q(\matmul0.matmul_stage_inst.d[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25299_ (.CLK(clknet_leaf_88_clk),
    .D(_00182_),
    .RESET_B(net8444),
    .Q(\matmul0.matmul_stage_inst.a[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25300_ (.CLK(clknet_leaf_76_clk),
    .D(_00183_),
    .RESET_B(net8460),
    .Q(\matmul0.matmul_stage_inst.e[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25301_ (.CLK(clknet_leaf_70_clk),
    .D(_00184_),
    .RESET_B(net8447),
    .Q(\matmul0.matmul_stage_inst.e[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25302_ (.CLK(clknet_leaf_70_clk),
    .D(_00185_),
    .RESET_B(net8459),
    .Q(\matmul0.matmul_stage_inst.e[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25303_ (.CLK(clknet_leaf_70_clk),
    .D(_00186_),
    .RESET_B(net8459),
    .Q(\matmul0.matmul_stage_inst.e[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25304_ (.CLK(clknet_leaf_69_clk),
    .D(_00187_),
    .RESET_B(net8451),
    .Q(\matmul0.matmul_stage_inst.e[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25305_ (.CLK(clknet_leaf_69_clk),
    .D(_00188_),
    .RESET_B(net8451),
    .Q(\matmul0.matmul_stage_inst.e[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25306_ (.CLK(clknet_leaf_71_clk),
    .D(_00189_),
    .RESET_B(net8461),
    .Q(\matmul0.matmul_stage_inst.e[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25307_ (.CLK(clknet_leaf_71_clk),
    .D(_00190_),
    .RESET_B(net8461),
    .Q(\matmul0.matmul_stage_inst.e[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25308_ (.CLK(clknet_leaf_72_clk),
    .D(_00191_),
    .RESET_B(net8469),
    .Q(\matmul0.matmul_stage_inst.e[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25309_ (.CLK(clknet_leaf_76_clk),
    .D(_00192_),
    .RESET_B(net8462),
    .Q(\matmul0.matmul_stage_inst.e[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25310_ (.CLK(clknet_leaf_76_clk),
    .D(_00193_),
    .RESET_B(net8462),
    .Q(\matmul0.matmul_stage_inst.e[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25311_ (.CLK(clknet_leaf_79_clk),
    .D(_00194_),
    .RESET_B(net8490),
    .Q(\matmul0.matmul_stage_inst.e[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25312_ (.CLK(clknet_leaf_80_clk),
    .D(_00195_),
    .RESET_B(net8511),
    .Q(\matmul0.matmul_stage_inst.e[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25313_ (.CLK(clknet_leaf_78_clk),
    .D(_00196_),
    .RESET_B(net8511),
    .Q(\matmul0.matmul_stage_inst.e[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25314_ (.CLK(clknet_leaf_79_clk),
    .D(_00197_),
    .RESET_B(net8490),
    .Q(\matmul0.matmul_stage_inst.e[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25315_ (.CLK(clknet_leaf_80_clk),
    .D(_00198_),
    .RESET_B(net8489),
    .Q(\matmul0.matmul_stage_inst.e[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25316_ (.CLK(clknet_leaf_75_clk),
    .D(_00199_),
    .RESET_B(net8463),
    .Q(\matmul0.matmul_stage_inst.f[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25317_ (.CLK(clknet_leaf_78_clk),
    .D(_00200_),
    .RESET_B(net8439),
    .Q(\matmul0.matmul_stage_inst.f[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25318_ (.CLK(clknet_leaf_75_clk),
    .D(_00201_),
    .RESET_B(net8463),
    .Q(\matmul0.matmul_stage_inst.f[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25319_ (.CLK(clknet_leaf_78_clk),
    .D(_00202_),
    .RESET_B(net8439),
    .Q(\matmul0.matmul_stage_inst.f[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25320_ (.CLK(clknet_leaf_75_clk),
    .D(_00203_),
    .RESET_B(net8463),
    .Q(\matmul0.matmul_stage_inst.f[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25321_ (.CLK(clknet_leaf_74_clk),
    .D(_00204_),
    .RESET_B(net8464),
    .Q(\matmul0.matmul_stage_inst.f[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25322_ (.CLK(clknet_leaf_75_clk),
    .D(_00205_),
    .RESET_B(net8467),
    .Q(\matmul0.matmul_stage_inst.f[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25323_ (.CLK(clknet_leaf_74_clk),
    .D(_00206_),
    .RESET_B(net8464),
    .Q(\matmul0.matmul_stage_inst.f[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25324_ (.CLK(clknet_leaf_75_clk),
    .D(_00207_),
    .RESET_B(net8464),
    .Q(\matmul0.matmul_stage_inst.f[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25325_ (.CLK(clknet_leaf_79_clk),
    .D(_00208_),
    .RESET_B(net8491),
    .Q(\matmul0.matmul_stage_inst.f[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25326_ (.CLK(clknet_leaf_79_clk),
    .D(_00209_),
    .RESET_B(net8491),
    .Q(\matmul0.matmul_stage_inst.f[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25327_ (.CLK(clknet_leaf_80_clk),
    .D(_00210_),
    .RESET_B(net8491),
    .Q(\matmul0.matmul_stage_inst.f[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25328_ (.CLK(clknet_leaf_80_clk),
    .D(_00211_),
    .RESET_B(net8497),
    .Q(\matmul0.matmul_stage_inst.f[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25329_ (.CLK(clknet_leaf_80_clk),
    .D(_00212_),
    .RESET_B(net8464),
    .Q(\matmul0.matmul_stage_inst.f[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25330_ (.CLK(clknet_leaf_80_clk),
    .D(_00213_),
    .RESET_B(net8488),
    .Q(\matmul0.matmul_stage_inst.f[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25331_ (.CLK(clknet_leaf_76_clk),
    .D(_00214_),
    .RESET_B(net8462),
    .Q(\matmul0.matmul_stage_inst.f[15] ));
 sky130_fd_sc_hd__dfrtp_2 _25332_ (.CLK(clknet_leaf_82_clk),
    .D(_00215_),
    .RESET_B(net8503),
    .Q(\matmul0.matmul_stage_inst.mult1[0] ));
 sky130_fd_sc_hd__dfrtp_2 _25333_ (.CLK(clknet_leaf_82_clk),
    .D(_00216_),
    .RESET_B(net8503),
    .Q(\matmul0.matmul_stage_inst.mult1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25334_ (.CLK(clknet_leaf_82_clk),
    .D(_00217_),
    .RESET_B(net8502),
    .Q(\matmul0.matmul_stage_inst.mult1[2] ));
 sky130_fd_sc_hd__dfrtp_2 _25335_ (.CLK(clknet_leaf_83_clk),
    .D(_00218_),
    .RESET_B(net8502),
    .Q(\matmul0.matmul_stage_inst.mult1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25336_ (.CLK(clknet_leaf_84_clk),
    .D(_00219_),
    .RESET_B(net8507),
    .Q(\matmul0.matmul_stage_inst.mult1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25337_ (.CLK(clknet_leaf_83_clk),
    .D(_00220_),
    .RESET_B(net8507),
    .Q(\matmul0.matmul_stage_inst.mult1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25338_ (.CLK(clknet_leaf_84_clk),
    .D(_00221_),
    .RESET_B(net8506),
    .Q(\matmul0.matmul_stage_inst.mult1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25339_ (.CLK(clknet_leaf_85_clk),
    .D(_00222_),
    .RESET_B(net8506),
    .Q(\matmul0.matmul_stage_inst.mult1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25340_ (.CLK(clknet_leaf_56_clk),
    .D(_00223_),
    .RESET_B(net8723),
    .Q(\matmul0.matmul_stage_inst.mult1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25341_ (.CLK(clknet_leaf_56_clk),
    .D(_00224_),
    .RESET_B(net8723),
    .Q(\matmul0.matmul_stage_inst.mult1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25342_ (.CLK(clknet_leaf_83_clk),
    .D(_00225_),
    .RESET_B(net8714),
    .Q(\matmul0.matmul_stage_inst.mult1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25343_ (.CLK(clknet_leaf_56_clk),
    .D(_00226_),
    .RESET_B(net8714),
    .Q(\matmul0.matmul_stage_inst.mult1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25344_ (.CLK(clknet_leaf_73_clk),
    .D(_00227_),
    .RESET_B(net8471),
    .Q(\matmul0.matmul_stage_inst.mult1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25345_ (.CLK(clknet_leaf_72_clk),
    .D(_00228_),
    .RESET_B(net8472),
    .Q(\matmul0.matmul_stage_inst.mult1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25346_ (.CLK(clknet_leaf_72_clk),
    .D(_00229_),
    .RESET_B(net8470),
    .Q(\matmul0.matmul_stage_inst.mult1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25347_ (.CLK(clknet_leaf_72_clk),
    .D(_00230_),
    .RESET_B(net8477),
    .Q(\matmul0.matmul_stage_inst.mult1[15] ));
 sky130_fd_sc_hd__dfrtp_2 _25348_ (.CLK(clknet_leaf_82_clk),
    .D(_00231_),
    .RESET_B(net8503),
    .Q(\matmul0.matmul_stage_inst.mult2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25349_ (.CLK(clknet_leaf_82_clk),
    .D(_00232_),
    .RESET_B(net8503),
    .Q(\matmul0.matmul_stage_inst.mult2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25350_ (.CLK(clknet_leaf_83_clk),
    .D(_00233_),
    .RESET_B(net8502),
    .Q(\matmul0.matmul_stage_inst.mult2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25351_ (.CLK(clknet_leaf_83_clk),
    .D(_00234_),
    .RESET_B(net8502),
    .Q(\matmul0.matmul_stage_inst.mult2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25352_ (.CLK(clknet_leaf_84_clk),
    .D(_00235_),
    .RESET_B(net8507),
    .Q(\matmul0.matmul_stage_inst.mult2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25353_ (.CLK(clknet_leaf_83_clk),
    .D(_00236_),
    .RESET_B(net8507),
    .Q(\matmul0.matmul_stage_inst.mult2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25354_ (.CLK(clknet_leaf_84_clk),
    .D(_00237_),
    .RESET_B(net8506),
    .Q(\matmul0.matmul_stage_inst.mult2[6] ));
 sky130_fd_sc_hd__dfstp_1 _25355_ (.CLK(clknet_leaf_42_clk),
    .D(_00238_),
    .SET_B(net8771),
    .Q(\svm0.delta[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25356_ (.CLK(clknet_leaf_85_clk),
    .D(_00239_),
    .RESET_B(net8513),
    .Q(\matmul0.matmul_stage_inst.mult2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25357_ (.CLK(clknet_leaf_84_clk),
    .D(_00240_),
    .RESET_B(net8723),
    .Q(\matmul0.matmul_stage_inst.mult2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25358_ (.CLK(clknet_leaf_56_clk),
    .D(_00241_),
    .RESET_B(net8723),
    .Q(\matmul0.matmul_stage_inst.mult2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25359_ (.CLK(clknet_leaf_56_clk),
    .D(_00242_),
    .RESET_B(net8718),
    .Q(\matmul0.matmul_stage_inst.mult2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25360_ (.CLK(clknet_leaf_57_clk),
    .D(_00243_),
    .RESET_B(net8718),
    .Q(\matmul0.matmul_stage_inst.mult2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25361_ (.CLK(clknet_leaf_72_clk),
    .D(_00244_),
    .RESET_B(net8477),
    .Q(\matmul0.matmul_stage_inst.mult2[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25362_ (.CLK(clknet_leaf_72_clk),
    .D(_00245_),
    .RESET_B(net8472),
    .Q(\matmul0.matmul_stage_inst.mult2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25363_ (.CLK(clknet_leaf_72_clk),
    .D(_00246_),
    .RESET_B(net8478),
    .Q(\matmul0.matmul_stage_inst.mult2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25364_ (.CLK(clknet_leaf_72_clk),
    .D(_00247_),
    .RESET_B(net8477),
    .Q(\matmul0.matmul_stage_inst.mult2[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25365_ (.CLK(clknet_leaf_72_clk),
    .D(_00248_),
    .RESET_B(net8478),
    .Q(\matmul0.alpha_pass[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25366_ (.CLK(clknet_leaf_81_clk),
    .D(_00249_),
    .RESET_B(net8495),
    .Q(\matmul0.alpha_pass[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25367_ (.CLK(clknet_leaf_81_clk),
    .D(_00250_),
    .RESET_B(net8496),
    .Q(\matmul0.alpha_pass[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25368_ (.CLK(clknet_leaf_81_clk),
    .D(_00251_),
    .RESET_B(net8498),
    .Q(\matmul0.alpha_pass[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25369_ (.CLK(clknet_leaf_81_clk),
    .D(_00252_),
    .RESET_B(net8500),
    .Q(\matmul0.alpha_pass[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25370_ (.CLK(clknet_leaf_81_clk),
    .D(_00253_),
    .RESET_B(net8500),
    .Q(\matmul0.alpha_pass[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25371_ (.CLK(clknet_leaf_57_clk),
    .D(_00254_),
    .RESET_B(net8711),
    .Q(\matmul0.alpha_pass[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25372_ (.CLK(clknet_leaf_81_clk),
    .D(_00255_),
    .RESET_B(net8709),
    .Q(\matmul0.alpha_pass[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25373_ (.CLK(clknet_leaf_63_clk),
    .D(_00256_),
    .RESET_B(net8708),
    .Q(\matmul0.alpha_pass[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25374_ (.CLK(clknet_leaf_57_clk),
    .D(_00257_),
    .RESET_B(net8710),
    .Q(\matmul0.alpha_pass[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25375_ (.CLK(clknet_leaf_57_clk),
    .D(_00258_),
    .RESET_B(net8716),
    .Q(\matmul0.alpha_pass[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25376_ (.CLK(clknet_leaf_58_clk),
    .D(_00259_),
    .RESET_B(net8726),
    .Q(\matmul0.alpha_pass[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25377_ (.CLK(clknet_leaf_64_clk),
    .D(_00260_),
    .RESET_B(net8663),
    .Q(\matmul0.alpha_pass[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25378_ (.CLK(clknet_leaf_63_clk),
    .D(_00261_),
    .RESET_B(net8667),
    .Q(\matmul0.alpha_pass[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25379_ (.CLK(clknet_leaf_64_clk),
    .D(_00262_),
    .RESET_B(net8663),
    .Q(\matmul0.alpha_pass[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25380_ (.CLK(clknet_leaf_64_clk),
    .D(_00263_),
    .RESET_B(net8663),
    .Q(\matmul0.alpha_pass[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25381_ (.CLK(clknet_leaf_74_clk),
    .D(_00264_),
    .RESET_B(net8466),
    .Q(\matmul0.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25382_ (.CLK(clknet_leaf_74_clk),
    .D(_00265_),
    .RESET_B(net8473),
    .Q(\matmul0.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25383_ (.CLK(clknet_leaf_73_clk),
    .D(_00266_),
    .RESET_B(net8476),
    .Q(\matmul0.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25384_ (.CLK(clknet_leaf_74_clk),
    .D(_00267_),
    .RESET_B(net8473),
    .Q(\matmul0.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25385_ (.CLK(clknet_leaf_73_clk),
    .D(_00268_),
    .RESET_B(net8474),
    .Q(\matmul0.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25386_ (.CLK(clknet_leaf_74_clk),
    .D(_00269_),
    .RESET_B(net8466),
    .Q(\matmul0.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25387_ (.CLK(clknet_leaf_73_clk),
    .D(_00270_),
    .RESET_B(net8473),
    .Q(\matmul0.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25388_ (.CLK(clknet_leaf_80_clk),
    .D(_00271_),
    .RESET_B(net8498),
    .Q(\matmul0.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25389_ (.CLK(clknet_leaf_74_clk),
    .D(_00272_),
    .RESET_B(net8466),
    .Q(\matmul0.b[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25390_ (.CLK(clknet_leaf_83_clk),
    .D(_00273_),
    .RESET_B(net8493),
    .Q(\matmul0.b[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25391_ (.CLK(clknet_leaf_79_clk),
    .D(_00274_),
    .RESET_B(net8493),
    .Q(\matmul0.b[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25392_ (.CLK(clknet_leaf_82_clk),
    .D(_00275_),
    .RESET_B(net8508),
    .Q(\matmul0.b[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25393_ (.CLK(clknet_leaf_80_clk),
    .D(_00276_),
    .RESET_B(net8497),
    .Q(\matmul0.b[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25394_ (.CLK(clknet_leaf_74_clk),
    .D(_00277_),
    .RESET_B(net8466),
    .Q(\matmul0.b[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25395_ (.CLK(clknet_leaf_74_clk),
    .D(_00278_),
    .RESET_B(net8498),
    .Q(\matmul0.b[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25396_ (.CLK(clknet_leaf_76_clk),
    .D(_00279_),
    .RESET_B(net8460),
    .Q(\matmul0.b[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25397_ (.CLK(clknet_leaf_71_clk),
    .D(_00280_),
    .RESET_B(net8461),
    .Q(\matmul0.a[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25398_ (.CLK(clknet_leaf_70_clk),
    .D(_00281_),
    .RESET_B(net8448),
    .Q(\matmul0.a[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25399_ (.CLK(clknet_leaf_70_clk),
    .D(_00282_),
    .RESET_B(net8451),
    .Q(\matmul0.a[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25400_ (.CLK(clknet_leaf_69_clk),
    .D(_00283_),
    .RESET_B(net8484),
    .Q(\matmul0.a[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25401_ (.CLK(clknet_leaf_68_clk),
    .D(_00284_),
    .RESET_B(net8450),
    .Q(\matmul0.a[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25402_ (.CLK(clknet_leaf_69_clk),
    .D(_00285_),
    .RESET_B(net8450),
    .Q(\matmul0.a[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25403_ (.CLK(clknet_leaf_72_clk),
    .D(_00286_),
    .RESET_B(net8469),
    .Q(\matmul0.a[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25404_ (.CLK(clknet_leaf_72_clk),
    .D(_00287_),
    .RESET_B(net8468),
    .Q(\matmul0.a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25405_ (.CLK(clknet_leaf_72_clk),
    .D(_00288_),
    .RESET_B(net8469),
    .Q(\matmul0.a[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25406_ (.CLK(clknet_leaf_76_clk),
    .D(_00289_),
    .RESET_B(net8472),
    .Q(\matmul0.a[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25407_ (.CLK(clknet_leaf_72_clk),
    .D(_00290_),
    .RESET_B(net8465),
    .Q(\matmul0.a[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25408_ (.CLK(clknet_leaf_80_clk),
    .D(_00291_),
    .RESET_B(net8489),
    .Q(\matmul0.a[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25409_ (.CLK(clknet_leaf_80_clk),
    .D(_00292_),
    .RESET_B(net8489),
    .Q(\matmul0.a[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25410_ (.CLK(clknet_leaf_75_clk),
    .D(_00293_),
    .RESET_B(net8511),
    .Q(\matmul0.a[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25411_ (.CLK(clknet_leaf_80_clk),
    .D(_00294_),
    .RESET_B(net8494),
    .Q(\matmul0.a[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25412_ (.CLK(clknet_leaf_80_clk),
    .D(_00295_),
    .RESET_B(net8494),
    .Q(\matmul0.a[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25413_ (.CLK(clknet_leaf_90_clk),
    .D(_00296_),
    .RESET_B(net8420),
    .Q(\matmul0.cos[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25414_ (.CLK(clknet_leaf_86_clk),
    .D(_00297_),
    .RESET_B(net8531),
    .Q(\matmul0.cos[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25415_ (.CLK(clknet_leaf_89_clk),
    .D(_00298_),
    .RESET_B(net8424),
    .Q(\matmul0.cos[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25416_ (.CLK(clknet_leaf_89_clk),
    .D(_00299_),
    .RESET_B(net8422),
    .Q(\matmul0.cos[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25417_ (.CLK(clknet_leaf_86_clk),
    .D(_00300_),
    .RESET_B(net8531),
    .Q(\matmul0.cos[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25418_ (.CLK(clknet_leaf_91_clk),
    .D(_00301_),
    .RESET_B(net8428),
    .Q(\matmul0.cos[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25419_ (.CLK(clknet_leaf_90_clk),
    .D(_00302_),
    .RESET_B(net8424),
    .Q(\matmul0.cos[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25420_ (.CLK(clknet_leaf_98_clk),
    .D(_00303_),
    .RESET_B(net8382),
    .Q(\matmul0.cos[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25421_ (.CLK(clknet_leaf_99_clk),
    .D(_00304_),
    .RESET_B(net8382),
    .Q(\matmul0.cos[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25422_ (.CLK(clknet_leaf_99_clk),
    .D(_00305_),
    .RESET_B(net8382),
    .Q(\matmul0.cos[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25423_ (.CLK(clknet_leaf_90_clk),
    .D(_00306_),
    .RESET_B(net8424),
    .Q(\matmul0.cos[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25424_ (.CLK(clknet_leaf_91_clk),
    .D(_00307_),
    .RESET_B(net8427),
    .Q(\matmul0.cos[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25425_ (.CLK(clknet_leaf_91_clk),
    .D(_00308_),
    .RESET_B(net8428),
    .Q(\matmul0.cos[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25426_ (.CLK(clknet_leaf_91_clk),
    .D(_00309_),
    .RESET_B(net8427),
    .Q(\matmul0.cos[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25427_ (.CLK(clknet_leaf_98_clk),
    .D(_00310_),
    .RESET_B(net8380),
    .Q(\matmul0.sin[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25428_ (.CLK(clknet_leaf_97_clk),
    .D(_00311_),
    .RESET_B(net8380),
    .Q(\matmul0.sin[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25429_ (.CLK(clknet_leaf_98_clk),
    .D(_00312_),
    .RESET_B(net8384),
    .Q(\matmul0.sin[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25430_ (.CLK(clknet_leaf_97_clk),
    .D(_00313_),
    .RESET_B(net8399),
    .Q(\matmul0.sin[3] ));
 sky130_fd_sc_hd__dfrtp_2 _25431_ (.CLK(clknet_leaf_94_clk),
    .D(_00314_),
    .RESET_B(net8445),
    .Q(\matmul0.sin[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25432_ (.CLK(clknet_leaf_96_clk),
    .D(_00315_),
    .RESET_B(net8399),
    .Q(\matmul0.sin[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25433_ (.CLK(clknet_leaf_97_clk),
    .D(_00316_),
    .RESET_B(net8400),
    .Q(\matmul0.sin[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25434_ (.CLK(clknet_leaf_94_clk),
    .D(_00317_),
    .RESET_B(net8445),
    .Q(\matmul0.sin[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25435_ (.CLK(clknet_leaf_96_clk),
    .D(_00318_),
    .RESET_B(net8445),
    .Q(\matmul0.sin[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25436_ (.CLK(clknet_leaf_97_clk),
    .D(_00319_),
    .RESET_B(net8399),
    .Q(\matmul0.sin[9] ));
 sky130_fd_sc_hd__dfrtp_4 _25437_ (.CLK(clknet_leaf_98_clk),
    .D(_00320_),
    .RESET_B(net8384),
    .Q(\matmul0.sin[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25438_ (.CLK(clknet_leaf_94_clk),
    .D(_00321_),
    .RESET_B(net8426),
    .Q(\matmul0.sin[11] ));
 sky130_fd_sc_hd__dfrtp_2 _25439_ (.CLK(clknet_leaf_91_clk),
    .D(_00322_),
    .RESET_B(net8426),
    .Q(\matmul0.sin[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25440_ (.CLK(clknet_leaf_91_clk),
    .D(_00323_),
    .RESET_B(net8432),
    .Q(\matmul0.sin[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25441_ (.CLK(clknet_leaf_113_clk),
    .D(_00324_),
    .RESET_B(net8340),
    .Q(\cordic0.vec[1][0] ));
 sky130_fd_sc_hd__dfrtp_1 _25442_ (.CLK(clknet_leaf_113_clk),
    .D(_00325_),
    .RESET_B(net8338),
    .Q(\cordic0.vec[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _25443_ (.CLK(clknet_leaf_113_clk),
    .D(_00326_),
    .RESET_B(net8340),
    .Q(\cordic0.vec[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _25444_ (.CLK(clknet_leaf_114_clk),
    .D(_00327_),
    .RESET_B(net8333),
    .Q(\cordic0.vec[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _25445_ (.CLK(clknet_leaf_117_clk),
    .D(_00328_),
    .RESET_B(net8332),
    .Q(\cordic0.vec[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _25446_ (.CLK(clknet_4_1__leaf_clk),
    .D(_00329_),
    .RESET_B(net8334),
    .Q(\cordic0.vec[1][5] ));
 sky130_fd_sc_hd__dfrtp_1 _25447_ (.CLK(clknet_leaf_114_clk),
    .D(_00330_),
    .RESET_B(net8334),
    .Q(\cordic0.vec[1][6] ));
 sky130_fd_sc_hd__dfrtp_1 _25448_ (.CLK(clknet_leaf_113_clk),
    .D(_00331_),
    .RESET_B(net8340),
    .Q(\cordic0.vec[1][7] ));
 sky130_fd_sc_hd__dfrtp_1 _25449_ (.CLK(clknet_leaf_119_clk),
    .D(_00332_),
    .RESET_B(net8338),
    .Q(\cordic0.vec[1][8] ));
 sky130_fd_sc_hd__dfrtp_1 _25450_ (.CLK(clknet_leaf_112_clk),
    .D(_00333_),
    .RESET_B(net8341),
    .Q(\cordic0.vec[1][9] ));
 sky130_fd_sc_hd__dfrtp_1 _25451_ (.CLK(clknet_leaf_119_clk),
    .D(_00334_),
    .RESET_B(net8342),
    .Q(\cordic0.vec[1][10] ));
 sky130_fd_sc_hd__dfrtp_1 _25452_ (.CLK(clknet_leaf_112_clk),
    .D(_00335_),
    .RESET_B(net8341),
    .Q(\cordic0.vec[1][11] ));
 sky130_fd_sc_hd__dfrtp_1 _25453_ (.CLK(clknet_leaf_112_clk),
    .D(_00336_),
    .RESET_B(net8539),
    .Q(\cordic0.vec[1][12] ));
 sky130_fd_sc_hd__dfrtp_1 _25454_ (.CLK(clknet_leaf_112_clk),
    .D(_00337_),
    .RESET_B(net8362),
    .Q(\cordic0.vec[1][13] ));
 sky130_fd_sc_hd__dfrtp_1 _25455_ (.CLK(clknet_4_1__leaf_clk),
    .D(_00338_),
    .RESET_B(net8362),
    .Q(\cordic0.vec[1][14] ));
 sky130_fd_sc_hd__dfrtp_1 _25456_ (.CLK(clknet_leaf_100_clk),
    .D(_00339_),
    .RESET_B(net8368),
    .Q(\cordic0.vec[1][15] ));
 sky130_fd_sc_hd__dfrtp_1 _25457_ (.CLK(clknet_leaf_100_clk),
    .D(_00340_),
    .RESET_B(net8389),
    .Q(\cordic0.vec[1][16] ));
 sky130_fd_sc_hd__dfrtp_1 _25458_ (.CLK(clknet_leaf_100_clk),
    .D(_00341_),
    .RESET_B(net8389),
    .Q(\cordic0.vec[1][17] ));
 sky130_fd_sc_hd__dfstp_1 _25459_ (.CLK(clknet_leaf_66_clk),
    .D(_00013_),
    .SET_B(net8662),
    .Q(\matmul0.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25460_ (.CLK(clknet_leaf_66_clk),
    .D(net8977),
    .RESET_B(net8647),
    .Q(\matmul0.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25461_ (.CLK(clknet_leaf_68_clk),
    .D(_00001_),
    .RESET_B(net8454),
    .Q(\matmul0.matmul_stage_inst.start ));
 sky130_fd_sc_hd__dfrtp_1 _25462_ (.CLK(clknet_leaf_53_clk),
    .D(_00342_),
    .RESET_B(net8804),
    .Q(\svm0.tB[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25463_ (.CLK(clknet_leaf_53_clk),
    .D(_00343_),
    .RESET_B(net8807),
    .Q(\svm0.tB[1] ));
 sky130_fd_sc_hd__dfrtp_2 _25464_ (.CLK(clknet_leaf_53_clk),
    .D(_00344_),
    .RESET_B(net8807),
    .Q(\svm0.tB[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25465_ (.CLK(clknet_leaf_53_clk),
    .D(_00345_),
    .RESET_B(net8807),
    .Q(\svm0.tB[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25466_ (.CLK(clknet_leaf_52_clk),
    .D(_00346_),
    .RESET_B(net8807),
    .Q(\svm0.tB[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25467_ (.CLK(clknet_leaf_53_clk),
    .D(_00347_),
    .RESET_B(net8807),
    .Q(\svm0.tB[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25468_ (.CLK(clknet_leaf_52_clk),
    .D(_00348_),
    .RESET_B(net8806),
    .Q(\svm0.tB[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25469_ (.CLK(clknet_leaf_52_clk),
    .D(_00349_),
    .RESET_B(net8806),
    .Q(\svm0.tB[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25470_ (.CLK(clknet_leaf_51_clk),
    .D(_00350_),
    .RESET_B(net8811),
    .Q(\svm0.tB[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25471_ (.CLK(clknet_leaf_46_clk),
    .D(_00351_),
    .RESET_B(net8811),
    .Q(\svm0.tB[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25472_ (.CLK(clknet_leaf_48_clk),
    .D(_00352_),
    .RESET_B(net8761),
    .Q(\svm0.tB[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25473_ (.CLK(clknet_leaf_46_clk),
    .D(_00353_),
    .RESET_B(net8774),
    .Q(\svm0.tB[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25474_ (.CLK(clknet_leaf_47_clk),
    .D(_00354_),
    .RESET_B(net8776),
    .Q(\svm0.tB[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25475_ (.CLK(clknet_leaf_47_clk),
    .D(_00355_),
    .RESET_B(net8775),
    .Q(\svm0.tB[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25476_ (.CLK(clknet_leaf_48_clk),
    .D(_00356_),
    .RESET_B(net8762),
    .Q(\svm0.tB[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25477_ (.CLK(clknet_leaf_48_clk),
    .D(_00357_),
    .RESET_B(net8762),
    .Q(\svm0.tB[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25478_ (.CLK(clknet_leaf_46_clk),
    .D(_00358_),
    .RESET_B(net8787),
    .Q(\svm0.tA[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25479_ (.CLK(clknet_leaf_45_clk),
    .D(_00359_),
    .RESET_B(net8787),
    .Q(\svm0.tA[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25480_ (.CLK(clknet_leaf_52_clk),
    .D(_00360_),
    .RESET_B(net8787),
    .Q(\svm0.tA[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25481_ (.CLK(clknet_leaf_45_clk),
    .D(_00361_),
    .RESET_B(net8789),
    .Q(\svm0.tA[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25482_ (.CLK(clknet_leaf_45_clk),
    .D(_00362_),
    .RESET_B(net8789),
    .Q(\svm0.tA[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25483_ (.CLK(clknet_leaf_45_clk),
    .D(_00363_),
    .RESET_B(net8787),
    .Q(\svm0.tA[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25484_ (.CLK(clknet_leaf_45_clk),
    .D(_00364_),
    .RESET_B(net8788),
    .Q(\svm0.tA[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25485_ (.CLK(clknet_leaf_45_clk),
    .D(_00365_),
    .RESET_B(net8788),
    .Q(\svm0.tA[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25486_ (.CLK(clknet_leaf_46_clk),
    .D(_00366_),
    .RESET_B(net8780),
    .Q(\svm0.tA[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25487_ (.CLK(clknet_leaf_46_clk),
    .D(_00367_),
    .RESET_B(net8780),
    .Q(\svm0.tA[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25488_ (.CLK(clknet_leaf_48_clk),
    .D(_00368_),
    .RESET_B(net8761),
    .Q(\svm0.tA[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25489_ (.CLK(clknet_leaf_48_clk),
    .D(_00369_),
    .RESET_B(net8779),
    .Q(\svm0.tA[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25490_ (.CLK(clknet_leaf_47_clk),
    .D(_00370_),
    .RESET_B(net8778),
    .Q(\svm0.tA[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25491_ (.CLK(clknet_leaf_47_clk),
    .D(_00371_),
    .RESET_B(net8775),
    .Q(\svm0.tA[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25492_ (.CLK(clknet_leaf_48_clk),
    .D(_00372_),
    .RESET_B(net8759),
    .Q(\svm0.tA[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25493_ (.CLK(clknet_leaf_48_clk),
    .D(_00373_),
    .RESET_B(net8762),
    .Q(\svm0.tA[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25494_ (.CLK(clknet_leaf_44_clk),
    .D(_00374_),
    .RESET_B(net8786),
    .Q(\svm0.calc_ready ));
 sky130_fd_sc_hd__dfstp_1 _25495_ (.CLK(clknet_leaf_48_clk),
    .D(_00375_),
    .SET_B(net8759),
    .Q(\svm0.rising ));
 sky130_fd_sc_hd__dfrtp_1 _25496_ (.CLK(clknet_leaf_42_clk),
    .D(_00376_),
    .RESET_B(net8771),
    .Q(\svm0.delta[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25497_ (.CLK(clknet_leaf_42_clk),
    .D(_00377_),
    .RESET_B(net8768),
    .Q(\svm0.delta[2] ));
 sky130_fd_sc_hd__dfrtp_2 _25498_ (.CLK(clknet_leaf_42_clk),
    .D(_00378_),
    .RESET_B(net8782),
    .Q(\svm0.delta[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25499_ (.CLK(clknet_leaf_41_clk),
    .D(_00379_),
    .RESET_B(net8782),
    .Q(\svm0.delta[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25500_ (.CLK(clknet_leaf_41_clk),
    .D(_00380_),
    .RESET_B(net8768),
    .Q(\svm0.delta[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25501_ (.CLK(clknet_leaf_41_clk),
    .D(_00381_),
    .RESET_B(net8768),
    .Q(\svm0.delta[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25502_ (.CLK(clknet_leaf_41_clk),
    .D(_00382_),
    .RESET_B(net8772),
    .Q(\svm0.delta[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25503_ (.CLK(clknet_leaf_39_clk),
    .D(_00383_),
    .RESET_B(net8771),
    .Q(\svm0.delta[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25504_ (.CLK(clknet_leaf_39_clk),
    .D(_00384_),
    .RESET_B(net8770),
    .Q(\svm0.delta[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25505_ (.CLK(clknet_leaf_39_clk),
    .D(_00385_),
    .RESET_B(net8770),
    .Q(\svm0.delta[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25506_ (.CLK(clknet_leaf_39_clk),
    .D(_00386_),
    .RESET_B(net8770),
    .Q(\svm0.delta[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25507_ (.CLK(clknet_leaf_39_clk),
    .D(_00387_),
    .RESET_B(net8754),
    .Q(\svm0.delta[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25508_ (.CLK(clknet_leaf_39_clk),
    .D(_00388_),
    .RESET_B(net8754),
    .Q(\svm0.delta[13] ));
 sky130_fd_sc_hd__dfrtp_2 _25509_ (.CLK(clknet_leaf_36_clk),
    .D(_00389_),
    .RESET_B(net8754),
    .Q(\svm0.delta[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25510_ (.CLK(clknet_leaf_36_clk),
    .D(_00390_),
    .RESET_B(net8758),
    .Q(\svm0.delta[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25511_ (.CLK(clknet_leaf_42_clk),
    .D(_00391_),
    .RESET_B(net8777),
    .Q(\svm0.counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25512_ (.CLK(clknet_leaf_43_clk),
    .D(_00392_),
    .RESET_B(net8778),
    .Q(\svm0.counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25513_ (.CLK(clknet_leaf_43_clk),
    .D(_00393_),
    .RESET_B(net8783),
    .Q(\svm0.counter[2] ));
 sky130_fd_sc_hd__dfrtp_4 _25514_ (.CLK(clknet_leaf_43_clk),
    .D(_00394_),
    .RESET_B(net8783),
    .Q(\svm0.counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25515_ (.CLK(clknet_leaf_44_clk),
    .D(_00395_),
    .RESET_B(net8783),
    .Q(\svm0.counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25516_ (.CLK(clknet_leaf_44_clk),
    .D(_00396_),
    .RESET_B(net8785),
    .Q(\svm0.counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25517_ (.CLK(clknet_leaf_41_clk),
    .D(_00397_),
    .RESET_B(net8784),
    .Q(\svm0.counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25518_ (.CLK(clknet_leaf_44_clk),
    .D(_00398_),
    .RESET_B(net8785),
    .Q(\svm0.counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25519_ (.CLK(clknet_leaf_42_clk),
    .D(_00399_),
    .RESET_B(net8777),
    .Q(\svm0.counter[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25520_ (.CLK(clknet_leaf_42_clk),
    .D(_00400_),
    .RESET_B(net8773),
    .Q(\svm0.counter[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25521_ (.CLK(clknet_leaf_47_clk),
    .D(_00401_),
    .RESET_B(net8777),
    .Q(\svm0.counter[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25522_ (.CLK(clknet_leaf_47_clk),
    .D(_00402_),
    .RESET_B(net8777),
    .Q(\svm0.counter[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25523_ (.CLK(clknet_leaf_48_clk),
    .D(_00403_),
    .RESET_B(net8756),
    .Q(\svm0.counter[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25524_ (.CLK(clknet_leaf_48_clk),
    .D(_00404_),
    .RESET_B(net8759),
    .Q(\svm0.counter[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25525_ (.CLK(clknet_leaf_35_clk),
    .D(_00405_),
    .RESET_B(net8758),
    .Q(\svm0.counter[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25526_ (.CLK(clknet_leaf_35_clk),
    .D(_00406_),
    .RESET_B(net8758),
    .Q(\svm0.counter[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25527_ (.CLK(clknet_leaf_45_clk),
    .D(net9001),
    .RESET_B(net8788),
    .Q(net151));
 sky130_fd_sc_hd__dfrtp_1 _25528_ (.CLK(clknet_leaf_45_clk),
    .D(net8963),
    .RESET_B(net8791),
    .Q(net150));
 sky130_fd_sc_hd__dfrtp_1 _25529_ (.CLK(clknet_leaf_45_clk),
    .D(_00409_),
    .RESET_B(net8791),
    .Q(net149));
 sky130_fd_sc_hd__dfrtp_1 _25530_ (.CLK(clknet_leaf_35_clk),
    .D(_00410_),
    .RESET_B(net8764),
    .Q(\svm0.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _25531_ (.CLK(clknet_leaf_35_clk),
    .D(_00411_),
    .RESET_B(net8764),
    .Q(\svm0.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25532_ (.CLK(clknet_leaf_47_clk),
    .D(_00412_),
    .RESET_B(net8776),
    .Q(\svm0.state[2] ));
 sky130_fd_sc_hd__dfstp_1 _25533_ (.CLK(clknet_leaf_35_clk),
    .D(_00413_),
    .SET_B(net8765),
    .Q(\svm0.ready ));
 sky130_fd_sc_hd__dfrtp_1 _25534_ (.CLK(clknet_leaf_32_clk),
    .D(_00414_),
    .RESET_B(net8692),
    .Q(\pid_q.prev_int[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25535_ (.CLK(clknet_4_12__leaf_clk),
    .D(_00415_),
    .RESET_B(net8695),
    .Q(\pid_q.prev_int[1] ));
 sky130_fd_sc_hd__dfrtp_2 _25536_ (.CLK(clknet_leaf_33_clk),
    .D(_00416_),
    .RESET_B(net8687),
    .Q(\pid_q.prev_int[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25537_ (.CLK(clknet_leaf_33_clk),
    .D(_00417_),
    .RESET_B(net8691),
    .Q(\pid_q.prev_int[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25538_ (.CLK(clknet_leaf_33_clk),
    .D(_00418_),
    .RESET_B(net8687),
    .Q(\pid_q.prev_int[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25539_ (.CLK(clknet_leaf_32_clk),
    .D(_00419_),
    .RESET_B(net8682),
    .Q(\pid_q.prev_int[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25540_ (.CLK(clknet_leaf_32_clk),
    .D(_00420_),
    .RESET_B(net8683),
    .Q(\pid_q.prev_int[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25541_ (.CLK(clknet_leaf_33_clk),
    .D(_00421_),
    .RESET_B(net8674),
    .Q(\pid_q.prev_int[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25542_ (.CLK(clknet_leaf_29_clk),
    .D(_00422_),
    .RESET_B(net8674),
    .Q(\pid_q.prev_int[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25543_ (.CLK(clknet_leaf_32_clk),
    .D(_00423_),
    .RESET_B(net8679),
    .Q(\pid_q.prev_int[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25544_ (.CLK(clknet_leaf_30_clk),
    .D(net9203),
    .RESET_B(net8676),
    .Q(\pid_q.prev_int[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25545_ (.CLK(clknet_leaf_28_clk),
    .D(_00425_),
    .RESET_B(net8652),
    .Q(\pid_q.prev_int[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25546_ (.CLK(clknet_leaf_28_clk),
    .D(_00426_),
    .RESET_B(net8652),
    .Q(\pid_q.prev_int[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25547_ (.CLK(clknet_leaf_28_clk),
    .D(_00427_),
    .RESET_B(net8649),
    .Q(\pid_q.prev_int[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25548_ (.CLK(clknet_leaf_30_clk),
    .D(_00428_),
    .RESET_B(net8673),
    .Q(\pid_q.prev_int[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25549_ (.CLK(clknet_leaf_28_clk),
    .D(_00429_),
    .RESET_B(net8649),
    .Q(\pid_q.prev_int[15] ));
 sky130_fd_sc_hd__dfstp_1 _25550_ (.CLK(clknet_leaf_66_clk),
    .D(_00012_),
    .SET_B(net8647),
    .Q(\matmul0.matmul_stage_inst.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25551_ (.CLK(clknet_leaf_69_clk),
    .D(net6555),
    .RESET_B(net8452),
    .Q(\matmul0.matmul_stage_inst.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25552_ (.CLK(clknet_leaf_79_clk),
    .D(net6592),
    .RESET_B(net8490),
    .Q(\matmul0.matmul_stage_inst.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25553_ (.CLK(clknet_leaf_64_clk),
    .D(net6572),
    .RESET_B(net8662),
    .Q(\matmul0.done_pass ));
 sky130_fd_sc_hd__dfrtp_1 _25554_ (.CLK(clknet_leaf_78_clk),
    .D(net3003),
    .RESET_B(net8439),
    .Q(\matmul0.matmul_stage_inst.state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25555_ (.CLK(clknet_leaf_72_clk),
    .D(net6632),
    .RESET_B(net8468),
    .Q(\matmul0.matmul_stage_inst.state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25556_ (.CLK(clknet_leaf_77_clk),
    .D(net6619),
    .RESET_B(net8439),
    .Q(\matmul0.matmul_stage_inst.state[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25557_ (.CLK(clknet_leaf_117_clk),
    .D(_00430_),
    .RESET_B(net8332),
    .Q(\cordic0.gm0.iter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25558_ (.CLK(clknet_leaf_111_clk),
    .D(_00431_),
    .RESET_B(net8365),
    .Q(\cordic0.gm0.iter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25559_ (.CLK(clknet_leaf_115_clk),
    .D(_00432_),
    .RESET_B(net8335),
    .Q(\cordic0.gm0.iter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25560_ (.CLK(clknet_leaf_115_clk),
    .D(_00433_),
    .RESET_B(net8335),
    .Q(\cordic0.gm0.iter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25561_ (.CLK(clknet_leaf_115_clk),
    .D(_00434_),
    .RESET_B(net8336),
    .Q(\cordic0.gm0.iter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25562_ (.CLK(clknet_leaf_64_clk),
    .D(_00435_),
    .RESET_B(net8670),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25563_ (.CLK(clknet_leaf_64_clk),
    .D(_00436_),
    .RESET_B(net8664),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25564_ (.CLK(clknet_leaf_66_clk),
    .D(_00437_),
    .RESET_B(net8659),
    .Q(\state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25565_ (.CLK(clknet_leaf_100_clk),
    .D(_00438_),
    .RESET_B(net8390),
    .Q(\cordic0.out_valid ));
 sky130_fd_sc_hd__dfrtp_1 _25566_ (.CLK(clknet_leaf_98_clk),
    .D(_00439_),
    .RESET_B(net8387),
    .Q(\cordic0.sin[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25567_ (.CLK(clknet_leaf_98_clk),
    .D(_00440_),
    .RESET_B(net8381),
    .Q(\cordic0.sin[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25568_ (.CLK(clknet_leaf_98_clk),
    .D(_00441_),
    .RESET_B(net8383),
    .Q(\cordic0.sin[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25569_ (.CLK(clknet_leaf_99_clk),
    .D(_00442_),
    .RESET_B(net8387),
    .Q(\cordic0.sin[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25570_ (.CLK(clknet_leaf_97_clk),
    .D(_00443_),
    .RESET_B(net8398),
    .Q(\cordic0.sin[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25571_ (.CLK(clknet_leaf_98_clk),
    .D(_00444_),
    .RESET_B(net8381),
    .Q(\cordic0.sin[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25572_ (.CLK(clknet_leaf_97_clk),
    .D(_00445_),
    .RESET_B(net8398),
    .Q(\cordic0.sin[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25573_ (.CLK(clknet_leaf_97_clk),
    .D(_00446_),
    .RESET_B(net8398),
    .Q(\cordic0.sin[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25574_ (.CLK(clknet_leaf_97_clk),
    .D(_00447_),
    .RESET_B(net8398),
    .Q(\cordic0.sin[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25575_ (.CLK(clknet_leaf_97_clk),
    .D(_00448_),
    .RESET_B(net8398),
    .Q(\cordic0.sin[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25576_ (.CLK(clknet_leaf_97_clk),
    .D(_00449_),
    .RESET_B(net8385),
    .Q(\cordic0.sin[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25577_ (.CLK(clknet_leaf_98_clk),
    .D(_00450_),
    .RESET_B(net8383),
    .Q(\cordic0.sin[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25578_ (.CLK(clknet_leaf_98_clk),
    .D(_00451_),
    .RESET_B(net8383),
    .Q(\cordic0.sin[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25579_ (.CLK(clknet_leaf_98_clk),
    .D(_00452_),
    .RESET_B(net8384),
    .Q(\cordic0.sin[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25580_ (.CLK(clknet_leaf_90_clk),
    .D(_00453_),
    .RESET_B(net8425),
    .Q(\cordic0.cos[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25581_ (.CLK(clknet_leaf_86_clk),
    .D(_00454_),
    .RESET_B(net8531),
    .Q(\cordic0.cos[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25582_ (.CLK(clknet_leaf_86_clk),
    .D(_00455_),
    .RESET_B(net8532),
    .Q(\cordic0.cos[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25583_ (.CLK(clknet_leaf_90_clk),
    .D(_00456_),
    .RESET_B(net8422),
    .Q(\cordic0.cos[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25584_ (.CLK(clknet_leaf_86_clk),
    .D(_00457_),
    .RESET_B(net8532),
    .Q(\cordic0.cos[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25585_ (.CLK(clknet_leaf_91_clk),
    .D(_00458_),
    .RESET_B(net8428),
    .Q(\cordic0.cos[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25586_ (.CLK(clknet_leaf_90_clk),
    .D(_00459_),
    .RESET_B(net8425),
    .Q(\cordic0.cos[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25587_ (.CLK(clknet_leaf_99_clk),
    .D(_00460_),
    .RESET_B(net8382),
    .Q(\cordic0.cos[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25588_ (.CLK(clknet_leaf_99_clk),
    .D(_00461_),
    .RESET_B(net8381),
    .Q(\cordic0.cos[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25589_ (.CLK(clknet_leaf_99_clk),
    .D(_00462_),
    .RESET_B(net8382),
    .Q(\cordic0.cos[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25590_ (.CLK(clknet_leaf_91_clk),
    .D(_00463_),
    .RESET_B(net8425),
    .Q(\cordic0.cos[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25591_ (.CLK(clknet_leaf_91_clk),
    .D(_00464_),
    .RESET_B(net8423),
    .Q(\cordic0.cos[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25592_ (.CLK(clknet_leaf_91_clk),
    .D(_00465_),
    .RESET_B(net8428),
    .Q(\cordic0.cos[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25593_ (.CLK(clknet_leaf_91_clk),
    .D(_00466_),
    .RESET_B(net8427),
    .Q(\cordic0.cos[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25594_ (.CLK(clknet_leaf_106_clk),
    .D(_00467_),
    .RESET_B(net8356),
    .Q(\cordic0.slte0.opB[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25595_ (.CLK(clknet_leaf_106_clk),
    .D(_00468_),
    .RESET_B(net8355),
    .Q(\cordic0.slte0.opB[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25596_ (.CLK(clknet_leaf_106_clk),
    .D(_00469_),
    .RESET_B(net8355),
    .Q(\cordic0.slte0.opB[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25597_ (.CLK(clknet_leaf_105_clk),
    .D(_00470_),
    .RESET_B(net8354),
    .Q(\cordic0.slte0.opB[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25598_ (.CLK(clknet_leaf_105_clk),
    .D(_00471_),
    .RESET_B(net8354),
    .Q(\cordic0.slte0.opB[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25599_ (.CLK(clknet_leaf_105_clk),
    .D(_00472_),
    .RESET_B(net8354),
    .Q(\cordic0.slte0.opB[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25600_ (.CLK(clknet_leaf_105_clk),
    .D(_00473_),
    .RESET_B(net8358),
    .Q(\cordic0.slte0.opB[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25601_ (.CLK(clknet_leaf_105_clk),
    .D(_00474_),
    .RESET_B(net8358),
    .Q(\cordic0.slte0.opB[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25602_ (.CLK(clknet_leaf_106_clk),
    .D(_00475_),
    .RESET_B(net8355),
    .Q(\cordic0.slte0.opB[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25603_ (.CLK(clknet_leaf_109_clk),
    .D(_00476_),
    .RESET_B(net8345),
    .Q(\cordic0.slte0.opB[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25604_ (.CLK(clknet_leaf_108_clk),
    .D(_00477_),
    .RESET_B(net8344),
    .Q(\cordic0.slte0.opB[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25605_ (.CLK(clknet_leaf_109_clk),
    .D(_00478_),
    .RESET_B(net8344),
    .Q(\cordic0.slte0.opB[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25606_ (.CLK(clknet_leaf_109_clk),
    .D(_00479_),
    .RESET_B(net8345),
    .Q(\cordic0.slte0.opB[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25607_ (.CLK(clknet_leaf_109_clk),
    .D(_00480_),
    .RESET_B(net8344),
    .Q(\cordic0.slte0.opB[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25608_ (.CLK(clknet_leaf_105_clk),
    .D(_00481_),
    .RESET_B(net8358),
    .Q(\cordic0.domain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25609_ (.CLK(clknet_leaf_105_clk),
    .D(_00482_),
    .RESET_B(net8356),
    .Q(\cordic0.domain[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25610_ (.CLK(clknet_leaf_108_clk),
    .D(_00483_),
    .RESET_B(net8350),
    .Q(\cordic0.slte0.opA[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25611_ (.CLK(clknet_leaf_108_clk),
    .D(_00484_),
    .RESET_B(net8349),
    .Q(\cordic0.slte0.opA[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25612_ (.CLK(clknet_leaf_111_clk),
    .D(_00485_),
    .RESET_B(net8349),
    .Q(\cordic0.slte0.opA[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25613_ (.CLK(clknet_leaf_109_clk),
    .D(_00486_),
    .RESET_B(net8352),
    .Q(\cordic0.slte0.opA[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25614_ (.CLK(clknet_leaf_108_clk),
    .D(_00487_),
    .RESET_B(net8351),
    .Q(\cordic0.slte0.opA[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25615_ (.CLK(clknet_leaf_109_clk),
    .D(_00488_),
    .RESET_B(net8346),
    .Q(\cordic0.slte0.opA[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25616_ (.CLK(clknet_leaf_109_clk),
    .D(_00489_),
    .RESET_B(net8346),
    .Q(\cordic0.slte0.opA[6] ));
 sky130_fd_sc_hd__dfrtp_4 _25617_ (.CLK(clknet_leaf_110_clk),
    .D(_00490_),
    .RESET_B(net8343),
    .Q(\cordic0.slte0.opA[7] ));
 sky130_fd_sc_hd__dfrtp_2 _25618_ (.CLK(clknet_leaf_110_clk),
    .D(_00491_),
    .RESET_B(net8347),
    .Q(\cordic0.slte0.opA[8] ));
 sky130_fd_sc_hd__dfrtp_4 _25619_ (.CLK(clknet_leaf_110_clk),
    .D(_00492_),
    .RESET_B(net8347),
    .Q(\cordic0.slte0.opA[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25620_ (.CLK(clknet_leaf_116_clk),
    .D(_00493_),
    .RESET_B(net8329),
    .Q(\cordic0.slte0.opA[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25621_ (.CLK(clknet_leaf_116_clk),
    .D(_00494_),
    .RESET_B(net8329),
    .Q(\cordic0.slte0.opA[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25622_ (.CLK(clknet_leaf_115_clk),
    .D(_00495_),
    .RESET_B(net8330),
    .Q(\cordic0.slte0.opA[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25623_ (.CLK(clknet_leaf_116_clk),
    .D(_00496_),
    .RESET_B(net8329),
    .Q(\cordic0.slte0.opA[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25624_ (.CLK(clknet_leaf_117_clk),
    .D(_00497_),
    .RESET_B(net8331),
    .Q(\cordic0.slte0.opA[14] ));
 sky130_fd_sc_hd__dfrtp_2 _25625_ (.CLK(clknet_leaf_117_clk),
    .D(_00498_),
    .RESET_B(net8332),
    .Q(\cordic0.slte0.opA[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25626_ (.CLK(clknet_leaf_117_clk),
    .D(_00499_),
    .RESET_B(net8337),
    .Q(\cordic0.slte0.opA[16] ));
 sky130_fd_sc_hd__dfrtp_1 _25627_ (.CLK(clknet_leaf_117_clk),
    .D(_00500_),
    .RESET_B(net8331),
    .Q(\cordic0.slte0.opA[17] ));
 sky130_fd_sc_hd__dfstp_1 _25628_ (.CLK(clknet_leaf_104_clk),
    .D(_00501_),
    .SET_B(net8357),
    .Q(\cordic0.vec[0][0] ));
 sky130_fd_sc_hd__dfstp_1 _25629_ (.CLK(clknet_leaf_108_clk),
    .D(_00502_),
    .SET_B(net8350),
    .Q(\cordic0.vec[0][1] ));
 sky130_fd_sc_hd__dfstp_1 _25630_ (.CLK(clknet_leaf_108_clk),
    .D(_00503_),
    .SET_B(net8351),
    .Q(\cordic0.vec[0][2] ));
 sky130_fd_sc_hd__dfstp_1 _25631_ (.CLK(clknet_leaf_106_clk),
    .D(_00504_),
    .SET_B(net8353),
    .Q(\cordic0.vec[0][3] ));
 sky130_fd_sc_hd__dfstp_1 _25632_ (.CLK(clknet_4_2__leaf_clk),
    .D(_00505_),
    .SET_B(net8357),
    .Q(\cordic0.vec[0][4] ));
 sky130_fd_sc_hd__dfstp_1 _25633_ (.CLK(clknet_leaf_105_clk),
    .D(_00506_),
    .SET_B(net8356),
    .Q(\cordic0.vec[0][5] ));
 sky130_fd_sc_hd__dfstp_1 _25634_ (.CLK(clknet_leaf_104_clk),
    .D(_00507_),
    .SET_B(net8361),
    .Q(\cordic0.vec[0][6] ));
 sky130_fd_sc_hd__dfstp_1 _25635_ (.CLK(clknet_leaf_104_clk),
    .D(_00508_),
    .SET_B(net8361),
    .Q(\cordic0.vec[0][7] ));
 sky130_fd_sc_hd__dfstp_1 _25636_ (.CLK(clknet_leaf_104_clk),
    .D(_00509_),
    .SET_B(net8359),
    .Q(\cordic0.vec[0][8] ));
 sky130_fd_sc_hd__dfstp_1 _25637_ (.CLK(clknet_leaf_103_clk),
    .D(_00510_),
    .SET_B(net8375),
    .Q(\cordic0.vec[0][9] ));
 sky130_fd_sc_hd__dfstp_1 _25638_ (.CLK(clknet_leaf_103_clk),
    .D(_00511_),
    .SET_B(net8375),
    .Q(\cordic0.vec[0][10] ));
 sky130_fd_sc_hd__dfstp_1 _25639_ (.CLK(clknet_leaf_102_clk),
    .D(_00512_),
    .SET_B(net8364),
    .Q(\cordic0.vec[0][11] ));
 sky130_fd_sc_hd__dfstp_1 _25640_ (.CLK(clknet_leaf_102_clk),
    .D(_00513_),
    .SET_B(net8366),
    .Q(\cordic0.vec[0][12] ));
 sky130_fd_sc_hd__dfstp_1 _25641_ (.CLK(clknet_leaf_103_clk),
    .D(_00514_),
    .SET_B(net8376),
    .Q(\cordic0.vec[0][13] ));
 sky130_fd_sc_hd__dfstp_1 _25642_ (.CLK(clknet_leaf_102_clk),
    .D(_00515_),
    .SET_B(net8366),
    .Q(\cordic0.vec[0][14] ));
 sky130_fd_sc_hd__dfstp_1 _25643_ (.CLK(clknet_leaf_102_clk),
    .D(_00516_),
    .SET_B(net8366),
    .Q(\cordic0.vec[0][15] ));
 sky130_fd_sc_hd__dfrtp_1 _25644_ (.CLK(clknet_leaf_102_clk),
    .D(_00517_),
    .RESET_B(net8367),
    .Q(\cordic0.vec[0][16] ));
 sky130_fd_sc_hd__dfrtp_1 _25645_ (.CLK(clknet_leaf_100_clk),
    .D(_00518_),
    .RESET_B(net8390),
    .Q(\cordic0.vec[0][17] ));
 sky130_fd_sc_hd__dfrtp_1 _25646_ (.CLK(clknet_leaf_1_clk),
    .D(_00519_),
    .RESET_B(net8403),
    .Q(\pid_d.curr_int[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25647_ (.CLK(clknet_leaf_122_clk),
    .D(_00520_),
    .RESET_B(net8403),
    .Q(\pid_d.curr_int[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25648_ (.CLK(clknet_leaf_122_clk),
    .D(_00521_),
    .RESET_B(net8407),
    .Q(\pid_d.curr_int[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25649_ (.CLK(clknet_leaf_1_clk),
    .D(_00522_),
    .RESET_B(net8403),
    .Q(\pid_d.curr_int[3] ));
 sky130_fd_sc_hd__dfrtp_2 _25650_ (.CLK(clknet_leaf_1_clk),
    .D(_00523_),
    .RESET_B(net8403),
    .Q(\pid_d.curr_int[4] ));
 sky130_fd_sc_hd__dfrtp_2 _25651_ (.CLK(clknet_leaf_1_clk),
    .D(_00524_),
    .RESET_B(net8404),
    .Q(\pid_d.curr_int[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25652_ (.CLK(clknet_leaf_1_clk),
    .D(_00525_),
    .RESET_B(net8401),
    .Q(\pid_d.curr_int[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25653_ (.CLK(clknet_leaf_2_clk),
    .D(_00526_),
    .RESET_B(net8570),
    .Q(\pid_d.curr_int[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25654_ (.CLK(clknet_leaf_2_clk),
    .D(_00527_),
    .RESET_B(net8570),
    .Q(\pid_d.curr_int[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25655_ (.CLK(clknet_leaf_2_clk),
    .D(_00528_),
    .RESET_B(net8573),
    .Q(\pid_d.curr_int[9] ));
 sky130_fd_sc_hd__dfrtp_4 _25656_ (.CLK(clknet_leaf_2_clk),
    .D(_00529_),
    .RESET_B(net8573),
    .Q(\pid_d.curr_int[10] ));
 sky130_fd_sc_hd__dfrtp_4 _25657_ (.CLK(clknet_leaf_25_clk),
    .D(_00530_),
    .RESET_B(net8577),
    .Q(\pid_d.curr_int[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25658_ (.CLK(clknet_leaf_3_clk),
    .D(_00531_),
    .RESET_B(net8580),
    .Q(\pid_d.curr_int[12] ));
 sky130_fd_sc_hd__dfrtp_4 _25659_ (.CLK(clknet_leaf_25_clk),
    .D(_00532_),
    .RESET_B(net8579),
    .Q(\pid_d.curr_int[13] ));
 sky130_fd_sc_hd__dfrtp_4 _25660_ (.CLK(clknet_leaf_24_clk),
    .D(_00533_),
    .RESET_B(net8584),
    .Q(\pid_d.curr_int[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25661_ (.CLK(clknet_leaf_24_clk),
    .D(_00534_),
    .RESET_B(net8584),
    .Q(\pid_d.curr_int[15] ));
 sky130_fd_sc_hd__dfrtp_2 _25662_ (.CLK(clknet_leaf_121_clk),
    .D(_00535_),
    .RESET_B(net8406),
    .Q(\pid_d.prev_error[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25663_ (.CLK(clknet_leaf_121_clk),
    .D(_00536_),
    .RESET_B(net8396),
    .Q(\pid_d.prev_error[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25664_ (.CLK(clknet_leaf_121_clk),
    .D(_00537_),
    .RESET_B(net8396),
    .Q(\pid_d.prev_error[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25665_ (.CLK(clknet_leaf_121_clk),
    .D(_00538_),
    .RESET_B(net8396),
    .Q(\pid_d.prev_error[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25666_ (.CLK(clknet_leaf_120_clk),
    .D(_00539_),
    .RESET_B(net8397),
    .Q(\pid_d.prev_error[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25667_ (.CLK(clknet_leaf_120_clk),
    .D(_00540_),
    .RESET_B(net8397),
    .Q(\pid_d.prev_error[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25668_ (.CLK(clknet_leaf_120_clk),
    .D(_00541_),
    .RESET_B(net8394),
    .Q(\pid_d.prev_error[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25669_ (.CLK(clknet_leaf_5_clk),
    .D(_00542_),
    .RESET_B(net8565),
    .Q(\pid_d.prev_error[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25670_ (.CLK(clknet_leaf_5_clk),
    .D(_00543_),
    .RESET_B(net8565),
    .Q(\pid_d.prev_error[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25671_ (.CLK(clknet_leaf_4_clk),
    .D(_00544_),
    .RESET_B(net8568),
    .Q(\pid_d.prev_error[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25672_ (.CLK(clknet_leaf_4_clk),
    .D(_00545_),
    .RESET_B(net8567),
    .Q(\pid_d.prev_error[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25673_ (.CLK(clknet_leaf_4_clk),
    .D(_00546_),
    .RESET_B(net8563),
    .Q(\pid_d.prev_error[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25674_ (.CLK(clknet_leaf_4_clk),
    .D(_00547_),
    .RESET_B(net8563),
    .Q(\pid_d.prev_error[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25675_ (.CLK(clknet_leaf_4_clk),
    .D(_00548_),
    .RESET_B(net8561),
    .Q(\pid_d.prev_error[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25676_ (.CLK(clknet_leaf_6_clk),
    .D(_00549_),
    .RESET_B(net8561),
    .Q(\pid_d.prev_error[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25677_ (.CLK(clknet_leaf_4_clk),
    .D(_00550_),
    .RESET_B(net8563),
    .Q(\pid_d.prev_error[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25678_ (.CLK(clknet_leaf_0_clk),
    .D(_00551_),
    .RESET_B(net8405),
    .Q(\pid_d.curr_error[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25679_ (.CLK(clknet_leaf_1_clk),
    .D(_00552_),
    .RESET_B(net8405),
    .Q(\pid_d.curr_error[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25680_ (.CLK(clknet_leaf_0_clk),
    .D(_00553_),
    .RESET_B(net8409),
    .Q(\pid_d.curr_error[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25681_ (.CLK(clknet_leaf_0_clk),
    .D(_00554_),
    .RESET_B(net8409),
    .Q(\pid_d.curr_error[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25682_ (.CLK(clknet_leaf_120_clk),
    .D(_00555_),
    .RESET_B(net8395),
    .Q(\pid_d.curr_error[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25683_ (.CLK(clknet_leaf_0_clk),
    .D(_00556_),
    .RESET_B(net8409),
    .Q(\pid_d.curr_error[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25684_ (.CLK(clknet_leaf_0_clk),
    .D(_00557_),
    .RESET_B(net8571),
    .Q(\pid_d.curr_error[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25685_ (.CLK(clknet_leaf_5_clk),
    .D(_00558_),
    .RESET_B(net8566),
    .Q(\pid_d.curr_error[7] ));
 sky130_fd_sc_hd__dfrtp_2 _25686_ (.CLK(clknet_leaf_3_clk),
    .D(_00559_),
    .RESET_B(net8572),
    .Q(\pid_d.curr_error[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25687_ (.CLK(clknet_leaf_2_clk),
    .D(_00560_),
    .RESET_B(net8572),
    .Q(\pid_d.curr_error[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25688_ (.CLK(clknet_leaf_5_clk),
    .D(_00561_),
    .RESET_B(net8567),
    .Q(\pid_d.curr_error[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25689_ (.CLK(clknet_leaf_3_clk),
    .D(_00562_),
    .RESET_B(net8569),
    .Q(\pid_d.curr_error[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25690_ (.CLK(clknet_leaf_6_clk),
    .D(_00563_),
    .RESET_B(net8562),
    .Q(\pid_d.curr_error[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25691_ (.CLK(clknet_leaf_3_clk),
    .D(_00564_),
    .RESET_B(net8569),
    .Q(\pid_d.curr_error[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25692_ (.CLK(clknet_leaf_6_clk),
    .D(_00565_),
    .RESET_B(net8562),
    .Q(\pid_d.curr_error[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25693_ (.CLK(clknet_leaf_3_clk),
    .D(_00566_),
    .RESET_B(net8569),
    .Q(\pid_d.curr_error[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25694_ (.CLK(clknet_leaf_121_clk),
    .D(_00567_),
    .RESET_B(net8395),
    .Q(\pid_d.mult0.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25695_ (.CLK(clknet_leaf_0_clk),
    .D(_00568_),
    .RESET_B(net8406),
    .Q(\pid_d.mult0.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25696_ (.CLK(clknet_leaf_3_clk),
    .D(_00569_),
    .RESET_B(net8575),
    .Q(\pid_d.mult0.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25697_ (.CLK(clknet_leaf_120_clk),
    .D(_00570_),
    .RESET_B(net8395),
    .Q(\pid_d.mult0.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25698_ (.CLK(clknet_leaf_120_clk),
    .D(_00571_),
    .RESET_B(net8395),
    .Q(\pid_d.mult0.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25699_ (.CLK(clknet_leaf_0_clk),
    .D(_00572_),
    .RESET_B(net8409),
    .Q(\pid_d.mult0.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25700_ (.CLK(clknet_leaf_120_clk),
    .D(_00573_),
    .RESET_B(net8414),
    .Q(\pid_d.mult0.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25701_ (.CLK(clknet_leaf_5_clk),
    .D(_00574_),
    .RESET_B(net8566),
    .Q(\pid_d.mult0.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25702_ (.CLK(clknet_leaf_2_clk),
    .D(_00575_),
    .RESET_B(net8572),
    .Q(\pid_d.mult0.b[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25703_ (.CLK(clknet_leaf_2_clk),
    .D(_00576_),
    .RESET_B(net8572),
    .Q(\pid_d.mult0.b[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25704_ (.CLK(clknet_leaf_5_clk),
    .D(_00577_),
    .RESET_B(net8567),
    .Q(\pid_d.mult0.b[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25705_ (.CLK(clknet_leaf_3_clk),
    .D(_00578_),
    .RESET_B(net8580),
    .Q(\pid_d.mult0.b[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25706_ (.CLK(clknet_leaf_6_clk),
    .D(_00579_),
    .RESET_B(net8562),
    .Q(\pid_d.mult0.b[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25707_ (.CLK(clknet_leaf_6_clk),
    .D(_00580_),
    .RESET_B(net8561),
    .Q(\pid_d.mult0.b[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25708_ (.CLK(clknet_leaf_6_clk),
    .D(_00581_),
    .RESET_B(net8564),
    .Q(\pid_d.mult0.b[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25709_ (.CLK(clknet_leaf_4_clk),
    .D(_00582_),
    .RESET_B(net8562),
    .Q(\pid_d.mult0.b[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25710_ (.CLK(clknet_leaf_9_clk),
    .D(_00583_),
    .RESET_B(net8552),
    .Q(\pid_d.mult0.a[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25711_ (.CLK(clknet_leaf_9_clk),
    .D(_00584_),
    .RESET_B(net8552),
    .Q(\pid_d.mult0.a[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25712_ (.CLK(clknet_leaf_9_clk),
    .D(_00585_),
    .RESET_B(net8552),
    .Q(\pid_d.mult0.a[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25713_ (.CLK(clknet_leaf_9_clk),
    .D(_00586_),
    .RESET_B(net8552),
    .Q(\pid_d.mult0.a[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25714_ (.CLK(clknet_leaf_9_clk),
    .D(_00587_),
    .RESET_B(net8559),
    .Q(\pid_d.mult0.a[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25715_ (.CLK(clknet_leaf_9_clk),
    .D(_00588_),
    .RESET_B(net8559),
    .Q(\pid_d.mult0.a[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25716_ (.CLK(clknet_leaf_9_clk),
    .D(_00589_),
    .RESET_B(net8559),
    .Q(\pid_d.mult0.a[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25717_ (.CLK(clknet_leaf_9_clk),
    .D(_00590_),
    .RESET_B(net8555),
    .Q(\pid_d.mult0.a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25718_ (.CLK(clknet_leaf_12_clk),
    .D(_00591_),
    .RESET_B(net8605),
    .Q(\pid_d.mult0.a[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25719_ (.CLK(clknet_leaf_11_clk),
    .D(_00592_),
    .RESET_B(net8602),
    .Q(\pid_d.mult0.a[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25720_ (.CLK(clknet_leaf_11_clk),
    .D(_00593_),
    .RESET_B(net8603),
    .Q(\pid_d.mult0.a[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25721_ (.CLK(clknet_leaf_13_clk),
    .D(_00594_),
    .RESET_B(net8603),
    .Q(\pid_d.mult0.a[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25722_ (.CLK(clknet_4_5__leaf_clk),
    .D(_00595_),
    .RESET_B(net8609),
    .Q(\pid_d.mult0.a[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25723_ (.CLK(clknet_leaf_13_clk),
    .D(_00596_),
    .RESET_B(net8609),
    .Q(\pid_d.mult0.a[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25724_ (.CLK(clknet_leaf_11_clk),
    .D(_00597_),
    .RESET_B(net8603),
    .Q(\pid_d.mult0.a[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25725_ (.CLK(clknet_leaf_13_clk),
    .D(_00598_),
    .RESET_B(net8609),
    .Q(\pid_d.mult0.a[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25726_ (.CLK(clknet_leaf_8_clk),
    .D(_00599_),
    .RESET_B(net8553),
    .Q(\pid_d.ki[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25727_ (.CLK(clknet_leaf_8_clk),
    .D(_00600_),
    .RESET_B(net8553),
    .Q(\pid_d.ki[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25728_ (.CLK(clknet_leaf_8_clk),
    .D(_00601_),
    .RESET_B(net8551),
    .Q(\pid_d.ki[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25729_ (.CLK(clknet_leaf_8_clk),
    .D(_00602_),
    .RESET_B(net8553),
    .Q(\pid_d.ki[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25730_ (.CLK(clknet_leaf_8_clk),
    .D(_00603_),
    .RESET_B(net8554),
    .Q(\pid_d.ki[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25731_ (.CLK(clknet_leaf_9_clk),
    .D(_00604_),
    .RESET_B(net8560),
    .Q(\pid_d.ki[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25732_ (.CLK(clknet_leaf_9_clk),
    .D(_00605_),
    .RESET_B(net8560),
    .Q(\pid_d.ki[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25733_ (.CLK(clknet_leaf_10_clk),
    .D(_00606_),
    .RESET_B(net8555),
    .Q(\pid_d.ki[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25734_ (.CLK(clknet_leaf_12_clk),
    .D(_00607_),
    .RESET_B(net8605),
    .Q(\pid_d.ki[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25735_ (.CLK(clknet_leaf_11_clk),
    .D(_00608_),
    .RESET_B(net8602),
    .Q(\pid_d.ki[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25736_ (.CLK(clknet_leaf_12_clk),
    .D(_00609_),
    .RESET_B(net8604),
    .Q(\pid_d.ki[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25737_ (.CLK(clknet_leaf_12_clk),
    .D(_00610_),
    .RESET_B(net8822),
    .Q(\pid_d.ki[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25738_ (.CLK(clknet_leaf_13_clk),
    .D(_00611_),
    .RESET_B(net8614),
    .Q(\pid_d.ki[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25739_ (.CLK(clknet_leaf_13_clk),
    .D(_00612_),
    .RESET_B(net8608),
    .Q(\pid_d.ki[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25740_ (.CLK(clknet_leaf_13_clk),
    .D(_00613_),
    .RESET_B(net8604),
    .Q(\pid_d.ki[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25741_ (.CLK(clknet_leaf_13_clk),
    .D(_00614_),
    .RESET_B(net8608),
    .Q(\pid_d.ki[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25742_ (.CLK(clknet_leaf_8_clk),
    .D(_00615_),
    .RESET_B(net8554),
    .Q(\pid_d.kp[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25743_ (.CLK(clknet_leaf_8_clk),
    .D(_00616_),
    .RESET_B(net8553),
    .Q(\pid_d.kp[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25744_ (.CLK(clknet_leaf_8_clk),
    .D(_00617_),
    .RESET_B(net8554),
    .Q(\pid_d.kp[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25745_ (.CLK(clknet_leaf_8_clk),
    .D(_00618_),
    .RESET_B(net8553),
    .Q(\pid_d.kp[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25746_ (.CLK(clknet_leaf_8_clk),
    .D(_00619_),
    .RESET_B(net8554),
    .Q(\pid_d.kp[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25747_ (.CLK(clknet_leaf_9_clk),
    .D(_00620_),
    .RESET_B(net8560),
    .Q(\pid_d.kp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25748_ (.CLK(clknet_leaf_9_clk),
    .D(_00621_),
    .RESET_B(net8601),
    .Q(\pid_d.kp[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25749_ (.CLK(clknet_leaf_10_clk),
    .D(_00622_),
    .RESET_B(net8590),
    .Q(\pid_d.kp[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25750_ (.CLK(clknet_leaf_12_clk),
    .D(_00623_),
    .RESET_B(net8605),
    .Q(\pid_d.kp[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25751_ (.CLK(clknet_leaf_11_clk),
    .D(_00624_),
    .RESET_B(net8602),
    .Q(\pid_d.kp[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25752_ (.CLK(clknet_leaf_13_clk),
    .D(_00625_),
    .RESET_B(net8604),
    .Q(\pid_d.kp[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25753_ (.CLK(clknet_leaf_12_clk),
    .D(_00626_),
    .RESET_B(net8604),
    .Q(\pid_d.kp[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25754_ (.CLK(clknet_leaf_13_clk),
    .D(_00627_),
    .RESET_B(net8614),
    .Q(\pid_d.kp[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25755_ (.CLK(clknet_leaf_13_clk),
    .D(_00628_),
    .RESET_B(net8608),
    .Q(\pid_d.kp[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25756_ (.CLK(clknet_leaf_13_clk),
    .D(_00629_),
    .RESET_B(net8606),
    .Q(\pid_d.kp[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25757_ (.CLK(clknet_leaf_13_clk),
    .D(_00630_),
    .RESET_B(net8608),
    .Q(\pid_d.kp[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25758_ (.CLK(clknet_leaf_27_clk),
    .D(_00631_),
    .RESET_B(net8645),
    .Q(\pid_d.out_valid ));
 sky130_fd_sc_hd__dfrtp_2 _25759_ (.CLK(clknet_leaf_95_clk),
    .D(_00632_),
    .RESET_B(net8402),
    .Q(\pid_d.out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25760_ (.CLK(clknet_leaf_95_clk),
    .D(_00633_),
    .RESET_B(net8455),
    .Q(\pid_d.out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25761_ (.CLK(clknet_leaf_95_clk),
    .D(_00634_),
    .RESET_B(net8455),
    .Q(\pid_d.out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _25762_ (.CLK(clknet_leaf_95_clk),
    .D(_00635_),
    .RESET_B(net8455),
    .Q(\pid_d.out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _25763_ (.CLK(clknet_leaf_67_clk),
    .D(_00636_),
    .RESET_B(net8455),
    .Q(\pid_d.out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25764_ (.CLK(clknet_leaf_67_clk),
    .D(_00637_),
    .RESET_B(net8456),
    .Q(\pid_d.out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25765_ (.CLK(clknet_leaf_67_clk),
    .D(_00638_),
    .RESET_B(net8453),
    .Q(\pid_d.out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25766_ (.CLK(clknet_leaf_67_clk),
    .D(_00639_),
    .RESET_B(net8646),
    .Q(\pid_d.out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25767_ (.CLK(clknet_leaf_27_clk),
    .D(_00640_),
    .RESET_B(net8646),
    .Q(\pid_d.out[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25768_ (.CLK(clknet_leaf_27_clk),
    .D(_00641_),
    .RESET_B(net8646),
    .Q(\pid_d.out[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25769_ (.CLK(clknet_leaf_26_clk),
    .D(_00642_),
    .RESET_B(net8576),
    .Q(\pid_d.out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25770_ (.CLK(clknet_leaf_27_clk),
    .D(_00643_),
    .RESET_B(net8650),
    .Q(\pid_d.out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25771_ (.CLK(clknet_leaf_27_clk),
    .D(_00644_),
    .RESET_B(net8650),
    .Q(\pid_d.out[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25772_ (.CLK(clknet_leaf_27_clk),
    .D(_00645_),
    .RESET_B(net8650),
    .Q(\pid_d.out[13] ));
 sky130_fd_sc_hd__dfrtp_2 _25773_ (.CLK(clknet_leaf_24_clk),
    .D(_00646_),
    .RESET_B(net8583),
    .Q(\pid_d.out[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25774_ (.CLK(clknet_leaf_26_clk),
    .D(_00647_),
    .RESET_B(net8650),
    .Q(\pid_d.out[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25775_ (.CLK(clknet_leaf_64_clk),
    .D(_00648_),
    .RESET_B(net8662),
    .Q(\matmul0.beta_pass[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25776_ (.CLK(clknet_leaf_57_clk),
    .D(_00649_),
    .RESET_B(net8711),
    .Q(\matmul0.beta_pass[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25777_ (.CLK(clknet_leaf_81_clk),
    .D(_00650_),
    .RESET_B(net8496),
    .Q(\matmul0.beta_pass[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25778_ (.CLK(clknet_leaf_74_clk),
    .D(_00651_),
    .RESET_B(net8473),
    .Q(\matmul0.beta_pass[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25779_ (.CLK(clknet_leaf_81_clk),
    .D(_00652_),
    .RESET_B(net8500),
    .Q(\matmul0.beta_pass[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25780_ (.CLK(clknet_leaf_73_clk),
    .D(_00653_),
    .RESET_B(net8499),
    .Q(\matmul0.beta_pass[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25781_ (.CLK(clknet_leaf_58_clk),
    .D(_00654_),
    .RESET_B(net8713),
    .Q(\matmul0.beta_pass[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25782_ (.CLK(clknet_leaf_82_clk),
    .D(_00655_),
    .RESET_B(net8500),
    .Q(\matmul0.beta_pass[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25783_ (.CLK(clknet_leaf_73_clk),
    .D(_00656_),
    .RESET_B(net8476),
    .Q(\matmul0.beta_pass[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25784_ (.CLK(clknet_leaf_57_clk),
    .D(_00657_),
    .RESET_B(net8709),
    .Q(\matmul0.beta_pass[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25785_ (.CLK(clknet_leaf_57_clk),
    .D(_00658_),
    .RESET_B(net8716),
    .Q(\matmul0.beta_pass[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25786_ (.CLK(clknet_leaf_58_clk),
    .D(_00659_),
    .RESET_B(net8712),
    .Q(\matmul0.beta_pass[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25787_ (.CLK(clknet_leaf_64_clk),
    .D(_00660_),
    .RESET_B(net8663),
    .Q(\matmul0.beta_pass[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25788_ (.CLK(clknet_leaf_63_clk),
    .D(_00661_),
    .RESET_B(net8672),
    .Q(\matmul0.beta_pass[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25789_ (.CLK(clknet_leaf_64_clk),
    .D(_00662_),
    .RESET_B(net8672),
    .Q(\matmul0.beta_pass[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25790_ (.CLK(clknet_leaf_64_clk),
    .D(_00663_),
    .RESET_B(net8668),
    .Q(\matmul0.beta_pass[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25791_ (.CLK(clknet_leaf_60_clk),
    .D(_00664_),
    .RESET_B(net8669),
    .Q(\svm0.in_valid ));
 sky130_fd_sc_hd__dfrtp_2 _25792_ (.CLK(clknet_leaf_32_clk),
    .D(_00665_),
    .RESET_B(net8681),
    .Q(\pid_q.curr_int[0] ));
 sky130_fd_sc_hd__dfrtp_2 _25793_ (.CLK(clknet_leaf_32_clk),
    .D(_00666_),
    .RESET_B(net8681),
    .Q(\pid_q.curr_int[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25794_ (.CLK(clknet_leaf_33_clk),
    .D(_00667_),
    .RESET_B(net8681),
    .Q(\pid_q.curr_int[2] ));
 sky130_fd_sc_hd__dfrtp_4 _25795_ (.CLK(clknet_leaf_33_clk),
    .D(_00668_),
    .RESET_B(net8678),
    .Q(\pid_q.curr_int[3] ));
 sky130_fd_sc_hd__dfrtp_4 _25796_ (.CLK(clknet_leaf_33_clk),
    .D(_00669_),
    .RESET_B(net8679),
    .Q(\pid_q.curr_int[4] ));
 sky130_fd_sc_hd__dfrtp_2 _25797_ (.CLK(clknet_leaf_32_clk),
    .D(_00670_),
    .RESET_B(net8682),
    .Q(\pid_q.curr_int[5] ));
 sky130_fd_sc_hd__dfrtp_2 _25798_ (.CLK(clknet_leaf_32_clk),
    .D(_00671_),
    .RESET_B(net8683),
    .Q(\pid_q.curr_int[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25799_ (.CLK(clknet_leaf_29_clk),
    .D(_00672_),
    .RESET_B(net8678),
    .Q(\pid_q.curr_int[7] ));
 sky130_fd_sc_hd__dfrtp_2 _25800_ (.CLK(clknet_leaf_30_clk),
    .D(_00673_),
    .RESET_B(net8677),
    .Q(\pid_q.curr_int[8] ));
 sky130_fd_sc_hd__dfrtp_2 _25801_ (.CLK(clknet_leaf_30_clk),
    .D(_00674_),
    .RESET_B(net8677),
    .Q(\pid_q.curr_int[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25802_ (.CLK(clknet_leaf_30_clk),
    .D(_00675_),
    .RESET_B(net8676),
    .Q(\pid_q.curr_int[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25803_ (.CLK(clknet_leaf_30_clk),
    .D(_00676_),
    .RESET_B(net8675),
    .Q(\pid_q.curr_int[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25804_ (.CLK(clknet_leaf_30_clk),
    .D(_00677_),
    .RESET_B(net8675),
    .Q(\pid_q.curr_int[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25805_ (.CLK(clknet_leaf_30_clk),
    .D(_00678_),
    .RESET_B(net8673),
    .Q(\pid_q.curr_int[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25806_ (.CLK(clknet_leaf_30_clk),
    .D(_00679_),
    .RESET_B(net8675),
    .Q(\pid_q.curr_int[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25807_ (.CLK(clknet_leaf_30_clk),
    .D(_00680_),
    .RESET_B(net8673),
    .Q(\pid_q.curr_int[15] ));
 sky130_fd_sc_hd__dfrtp_4 _25808_ (.CLK(clknet_leaf_38_clk),
    .D(_00681_),
    .RESET_B(net8755),
    .Q(\pid_q.prev_error[0] ));
 sky130_fd_sc_hd__dfrtp_2 _25809_ (.CLK(clknet_leaf_38_clk),
    .D(_00682_),
    .RESET_B(net8755),
    .Q(\pid_q.prev_error[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25810_ (.CLK(clknet_leaf_36_clk),
    .D(_00683_),
    .RESET_B(net8797),
    .Q(\pid_q.prev_error[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25811_ (.CLK(clknet_leaf_36_clk),
    .D(_00684_),
    .RESET_B(net8797),
    .Q(\pid_q.prev_error[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25812_ (.CLK(clknet_leaf_36_clk),
    .D(_00685_),
    .RESET_B(net8748),
    .Q(\pid_q.prev_error[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25813_ (.CLK(clknet_leaf_36_clk),
    .D(_00686_),
    .RESET_B(net8748),
    .Q(\pid_q.prev_error[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25814_ (.CLK(clknet_leaf_32_clk),
    .D(_00687_),
    .RESET_B(net8680),
    .Q(\pid_q.prev_error[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25815_ (.CLK(clknet_leaf_37_clk),
    .D(_00688_),
    .RESET_B(net8749),
    .Q(\pid_q.prev_error[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25816_ (.CLK(clknet_leaf_37_clk),
    .D(_00689_),
    .RESET_B(net8750),
    .Q(\pid_q.prev_error[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25817_ (.CLK(clknet_leaf_37_clk),
    .D(_00690_),
    .RESET_B(net8746),
    .Q(\pid_q.prev_error[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25818_ (.CLK(clknet_leaf_37_clk),
    .D(_00691_),
    .RESET_B(net8744),
    .Q(\pid_q.prev_error[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25819_ (.CLK(clknet_leaf_32_clk),
    .D(_00692_),
    .RESET_B(net8685),
    .Q(\pid_q.prev_error[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25820_ (.CLK(clknet_leaf_31_clk),
    .D(_00693_),
    .RESET_B(net8686),
    .Q(\pid_q.prev_error[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25821_ (.CLK(clknet_leaf_31_clk),
    .D(_00694_),
    .RESET_B(net8686),
    .Q(\pid_q.prev_error[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25822_ (.CLK(clknet_leaf_30_clk),
    .D(_00695_),
    .RESET_B(net8686),
    .Q(\pid_q.prev_error[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25823_ (.CLK(clknet_leaf_31_clk),
    .D(_00696_),
    .RESET_B(net8684),
    .Q(\pid_q.prev_error[15] ));
 sky130_fd_sc_hd__dfrtp_4 _25824_ (.CLK(clknet_leaf_38_clk),
    .D(_00697_),
    .RESET_B(net8746),
    .Q(\pid_q.curr_error[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25825_ (.CLK(clknet_leaf_37_clk),
    .D(_00698_),
    .RESET_B(net8744),
    .Q(\pid_q.curr_error[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25826_ (.CLK(clknet_leaf_36_clk),
    .D(_00699_),
    .RESET_B(net8750),
    .Q(\pid_q.curr_error[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25827_ (.CLK(clknet_leaf_36_clk),
    .D(_00700_),
    .RESET_B(net8748),
    .Q(\pid_q.curr_error[3] ));
 sky130_fd_sc_hd__dfrtp_2 _25828_ (.CLK(clknet_leaf_36_clk),
    .D(_00701_),
    .RESET_B(net8753),
    .Q(\pid_q.curr_error[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25829_ (.CLK(clknet_leaf_36_clk),
    .D(_00702_),
    .RESET_B(net8752),
    .Q(\pid_q.curr_error[5] ));
 sky130_fd_sc_hd__dfrtp_2 _25830_ (.CLK(clknet_leaf_37_clk),
    .D(_00703_),
    .RESET_B(net8680),
    .Q(\pid_q.curr_error[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25831_ (.CLK(clknet_leaf_36_clk),
    .D(_00704_),
    .RESET_B(net8752),
    .Q(\pid_q.curr_error[7] ));
 sky130_fd_sc_hd__dfrtp_2 _25832_ (.CLK(clknet_leaf_36_clk),
    .D(_00705_),
    .RESET_B(net8753),
    .Q(\pid_q.curr_error[8] ));
 sky130_fd_sc_hd__dfrtp_2 _25833_ (.CLK(clknet_leaf_37_clk),
    .D(_00706_),
    .RESET_B(net8746),
    .Q(\pid_q.curr_error[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25834_ (.CLK(clknet_leaf_37_clk),
    .D(_00707_),
    .RESET_B(net8745),
    .Q(\pid_q.curr_error[10] ));
 sky130_fd_sc_hd__dfrtp_2 _25835_ (.CLK(clknet_leaf_31_clk),
    .D(_00708_),
    .RESET_B(net8696),
    .Q(\pid_q.curr_error[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25836_ (.CLK(clknet_leaf_31_clk),
    .D(_00709_),
    .RESET_B(net8685),
    .Q(\pid_q.curr_error[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25837_ (.CLK(clknet_leaf_31_clk),
    .D(_00710_),
    .RESET_B(net8684),
    .Q(\pid_q.curr_error[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25838_ (.CLK(clknet_leaf_31_clk),
    .D(_00711_),
    .RESET_B(net8684),
    .Q(\pid_q.curr_error[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25839_ (.CLK(clknet_leaf_31_clk),
    .D(_00712_),
    .RESET_B(net8684),
    .Q(\pid_q.curr_error[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25840_ (.CLK(clknet_leaf_38_clk),
    .D(_00713_),
    .RESET_B(net8743),
    .Q(\pid_q.mult0.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25841_ (.CLK(clknet_leaf_20_clk),
    .D(_00714_),
    .RESET_B(net8610),
    .Q(\pid_q.mult0.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25842_ (.CLK(clknet_leaf_20_clk),
    .D(_00715_),
    .RESET_B(net8743),
    .Q(\pid_q.mult0.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25843_ (.CLK(clknet_leaf_20_clk),
    .D(_00716_),
    .RESET_B(net8747),
    .Q(\pid_q.mult0.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25844_ (.CLK(clknet_leaf_38_clk),
    .D(_00717_),
    .RESET_B(net8747),
    .Q(\pid_q.mult0.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25845_ (.CLK(clknet_leaf_38_clk),
    .D(_00718_),
    .RESET_B(net8747),
    .Q(\pid_q.mult0.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25846_ (.CLK(clknet_leaf_20_clk),
    .D(_00719_),
    .RESET_B(net8616),
    .Q(\pid_q.mult0.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25847_ (.CLK(clknet_leaf_20_clk),
    .D(_00720_),
    .RESET_B(net8616),
    .Q(\pid_q.mult0.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25848_ (.CLK(clknet_leaf_20_clk),
    .D(_00721_),
    .RESET_B(net8615),
    .Q(\pid_q.mult0.b[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25849_ (.CLK(clknet_leaf_20_clk),
    .D(_00722_),
    .RESET_B(net8616),
    .Q(\pid_q.mult0.b[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25850_ (.CLK(clknet_leaf_20_clk),
    .D(_00723_),
    .RESET_B(net8745),
    .Q(\pid_q.mult0.b[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25851_ (.CLK(clknet_leaf_20_clk),
    .D(_00724_),
    .RESET_B(net8616),
    .Q(\pid_q.mult0.b[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25852_ (.CLK(clknet_leaf_23_clk),
    .D(_00725_),
    .RESET_B(net8586),
    .Q(\pid_q.mult0.b[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25853_ (.CLK(clknet_leaf_38_clk),
    .D(_00726_),
    .RESET_B(net8745),
    .Q(\pid_q.mult0.b[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25854_ (.CLK(clknet_leaf_23_clk),
    .D(_00727_),
    .RESET_B(net8586),
    .Q(\pid_q.mult0.b[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25855_ (.CLK(clknet_leaf_23_clk),
    .D(_00728_),
    .RESET_B(net8586),
    .Q(\pid_q.mult0.b[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25856_ (.CLK(clknet_leaf_19_clk),
    .D(_00729_),
    .RESET_B(net8624),
    .Q(\pid_q.mult0.a[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25857_ (.CLK(clknet_leaf_19_clk),
    .D(_00730_),
    .RESET_B(net8624),
    .Q(\pid_q.mult0.a[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25858_ (.CLK(clknet_leaf_16_clk),
    .D(_00731_),
    .RESET_B(net8619),
    .Q(\pid_q.mult0.a[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25859_ (.CLK(clknet_leaf_16_clk),
    .D(_00732_),
    .RESET_B(net8619),
    .Q(\pid_q.mult0.a[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25860_ (.CLK(clknet_leaf_16_clk),
    .D(_00733_),
    .RESET_B(net8619),
    .Q(\pid_q.mult0.a[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25861_ (.CLK(clknet_leaf_15_clk),
    .D(_00734_),
    .RESET_B(net8617),
    .Q(\pid_q.mult0.a[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25862_ (.CLK(clknet_leaf_14_clk),
    .D(_00735_),
    .RESET_B(net8617),
    .Q(\pid_q.mult0.a[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25863_ (.CLK(clknet_leaf_15_clk),
    .D(_00736_),
    .RESET_B(net8617),
    .Q(\pid_q.mult0.a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25864_ (.CLK(clknet_leaf_16_clk),
    .D(_00737_),
    .RESET_B(net8619),
    .Q(\pid_q.mult0.a[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25865_ (.CLK(clknet_leaf_16_clk),
    .D(_00738_),
    .RESET_B(net8619),
    .Q(\pid_q.mult0.a[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25866_ (.CLK(clknet_leaf_16_clk),
    .D(_00739_),
    .RESET_B(net8625),
    .Q(\pid_q.mult0.a[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25867_ (.CLK(clknet_leaf_16_clk),
    .D(_00740_),
    .RESET_B(net8625),
    .Q(\pid_q.mult0.a[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25868_ (.CLK(clknet_leaf_17_clk),
    .D(_00741_),
    .RESET_B(net8624),
    .Q(\pid_q.mult0.a[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25869_ (.CLK(clknet_leaf_18_clk),
    .D(_00742_),
    .RESET_B(net8630),
    .Q(\pid_q.mult0.a[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25870_ (.CLK(clknet_leaf_17_clk),
    .D(_00743_),
    .RESET_B(net8631),
    .Q(\pid_q.mult0.a[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25871_ (.CLK(clknet_leaf_18_clk),
    .D(_00744_),
    .RESET_B(net8630),
    .Q(\pid_q.mult0.a[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25872_ (.CLK(clknet_leaf_17_clk),
    .D(_00745_),
    .RESET_B(net8626),
    .Q(\pid_q.ki[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25873_ (.CLK(clknet_leaf_17_clk),
    .D(_00746_),
    .RESET_B(net8626),
    .Q(\pid_q.ki[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25874_ (.CLK(clknet_leaf_14_clk),
    .D(_00747_),
    .RESET_B(net8621),
    .Q(\pid_q.ki[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25875_ (.CLK(clknet_leaf_15_clk),
    .D(_00748_),
    .RESET_B(net8618),
    .Q(\pid_q.ki[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25876_ (.CLK(clknet_leaf_15_clk),
    .D(_00749_),
    .RESET_B(net8618),
    .Q(\pid_q.ki[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25877_ (.CLK(clknet_leaf_14_clk),
    .D(_00750_),
    .RESET_B(net8620),
    .Q(\pid_q.ki[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25878_ (.CLK(clknet_leaf_14_clk),
    .D(_00751_),
    .RESET_B(net8621),
    .Q(\pid_q.ki[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25879_ (.CLK(clknet_leaf_14_clk),
    .D(_00752_),
    .RESET_B(net8621),
    .Q(\pid_q.ki[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25880_ (.CLK(clknet_leaf_15_clk),
    .D(_00753_),
    .RESET_B(net8622),
    .Q(\pid_q.ki[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25881_ (.CLK(clknet_leaf_14_clk),
    .D(_00754_),
    .RESET_B(net8620),
    .Q(\pid_q.ki[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25882_ (.CLK(clknet_leaf_16_clk),
    .D(_00755_),
    .RESET_B(net8625),
    .Q(\pid_q.ki[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25883_ (.CLK(clknet_leaf_16_clk),
    .D(_00756_),
    .RESET_B(net8625),
    .Q(\pid_q.ki[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25884_ (.CLK(clknet_leaf_17_clk),
    .D(_00757_),
    .RESET_B(net8626),
    .Q(\pid_q.ki[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25885_ (.CLK(clknet_leaf_18_clk),
    .D(_00758_),
    .RESET_B(net8630),
    .Q(\pid_q.ki[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25886_ (.CLK(clknet_leaf_17_clk),
    .D(_00759_),
    .RESET_B(net8632),
    .Q(\pid_q.ki[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25887_ (.CLK(clknet_leaf_40_clk),
    .D(_00760_),
    .RESET_B(net8769),
    .Q(\pid_q.ki[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25888_ (.CLK(clknet_leaf_17_clk),
    .D(_00761_),
    .RESET_B(net8628),
    .Q(\pid_q.kp[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25889_ (.CLK(clknet_leaf_17_clk),
    .D(_00762_),
    .RESET_B(net8628),
    .Q(\pid_q.kp[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25890_ (.CLK(clknet_leaf_14_clk),
    .D(_00763_),
    .RESET_B(net8621),
    .Q(\pid_q.kp[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25891_ (.CLK(clknet_leaf_16_clk),
    .D(_00764_),
    .RESET_B(net8622),
    .Q(\pid_q.kp[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25892_ (.CLK(clknet_leaf_15_clk),
    .D(_00765_),
    .RESET_B(net8622),
    .Q(\pid_q.kp[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25893_ (.CLK(clknet_leaf_14_clk),
    .D(_00766_),
    .RESET_B(net8620),
    .Q(\pid_q.kp[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25894_ (.CLK(clknet_leaf_14_clk),
    .D(_00767_),
    .RESET_B(net8621),
    .Q(\pid_q.kp[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25895_ (.CLK(clknet_leaf_14_clk),
    .D(_00768_),
    .RESET_B(net8621),
    .Q(\pid_q.kp[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25896_ (.CLK(clknet_leaf_15_clk),
    .D(_00769_),
    .RESET_B(net8622),
    .Q(\pid_q.kp[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25897_ (.CLK(clknet_leaf_14_clk),
    .D(_00770_),
    .RESET_B(net8620),
    .Q(\pid_q.kp[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25898_ (.CLK(clknet_leaf_16_clk),
    .D(_00771_),
    .RESET_B(net8627),
    .Q(\pid_q.kp[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25899_ (.CLK(clknet_leaf_16_clk),
    .D(_00772_),
    .RESET_B(net8627),
    .Q(\pid_q.kp[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25900_ (.CLK(clknet_leaf_17_clk),
    .D(_00773_),
    .RESET_B(net8628),
    .Q(\pid_q.kp[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25901_ (.CLK(clknet_leaf_17_clk),
    .D(_00774_),
    .RESET_B(net8630),
    .Q(\pid_q.kp[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25902_ (.CLK(clknet_leaf_17_clk),
    .D(_00775_),
    .RESET_B(net8632),
    .Q(\pid_q.kp[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25903_ (.CLK(clknet_leaf_40_clk),
    .D(_00776_),
    .RESET_B(net8769),
    .Q(\pid_q.kp[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25904_ (.CLK(clknet_leaf_65_clk),
    .D(_00777_),
    .RESET_B(net8654),
    .Q(\pid_q.out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _25905_ (.CLK(clknet_leaf_65_clk),
    .D(_00778_),
    .RESET_B(net8703),
    .Q(\pid_q.out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25906_ (.CLK(clknet_leaf_65_clk),
    .D(_00779_),
    .RESET_B(net8703),
    .Q(\pid_q.out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25907_ (.CLK(clknet_leaf_60_clk),
    .D(_00780_),
    .RESET_B(net8691),
    .Q(\pid_q.out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25908_ (.CLK(clknet_leaf_33_clk),
    .D(_00781_),
    .RESET_B(net8691),
    .Q(\pid_q.out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25909_ (.CLK(clknet_leaf_29_clk),
    .D(_00782_),
    .RESET_B(net8656),
    .Q(\pid_q.out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25910_ (.CLK(clknet_leaf_28_clk),
    .D(_00783_),
    .RESET_B(net8656),
    .Q(\pid_q.out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25911_ (.CLK(clknet_leaf_29_clk),
    .D(_00784_),
    .RESET_B(net8654),
    .Q(\pid_q.out[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25912_ (.CLK(clknet_leaf_66_clk),
    .D(_00785_),
    .RESET_B(net8659),
    .Q(\pid_q.out[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25913_ (.CLK(clknet_leaf_66_clk),
    .D(_00786_),
    .RESET_B(net8659),
    .Q(\pid_q.out[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25914_ (.CLK(clknet_leaf_67_clk),
    .D(_00787_),
    .RESET_B(net8648),
    .Q(\pid_q.out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25915_ (.CLK(clknet_leaf_27_clk),
    .D(_00788_),
    .RESET_B(net8648),
    .Q(\pid_q.out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25916_ (.CLK(clknet_leaf_27_clk),
    .D(_00789_),
    .RESET_B(net8651),
    .Q(\pid_q.out[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25917_ (.CLK(clknet_leaf_28_clk),
    .D(_00790_),
    .RESET_B(net8657),
    .Q(\pid_q.out[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25918_ (.CLK(clknet_leaf_28_clk),
    .D(_00791_),
    .RESET_B(net8651),
    .Q(\pid_q.out[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25919_ (.CLK(clknet_leaf_28_clk),
    .D(_00792_),
    .RESET_B(net8656),
    .Q(\pid_q.out[15] ));
 sky130_fd_sc_hd__dfrtp_1 _25920_ (.CLK(clknet_leaf_96_clk),
    .D(_00793_),
    .RESET_B(net8400),
    .Q(\pid_d.prev_int[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25921_ (.CLK(clknet_leaf_97_clk),
    .D(_00794_),
    .RESET_B(net8412),
    .Q(\pid_d.prev_int[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25922_ (.CLK(clknet_leaf_96_clk),
    .D(_00795_),
    .RESET_B(net8412),
    .Q(\pid_d.prev_int[2] ));
 sky130_fd_sc_hd__dfrtp_2 _25923_ (.CLK(clknet_leaf_96_clk),
    .D(_00796_),
    .RESET_B(net8402),
    .Q(\pid_d.prev_int[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25924_ (.CLK(clknet_leaf_1_clk),
    .D(_00797_),
    .RESET_B(net8404),
    .Q(\pid_d.prev_int[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25925_ (.CLK(clknet_leaf_1_clk),
    .D(_00798_),
    .RESET_B(net8404),
    .Q(\pid_d.prev_int[5] ));
 sky130_fd_sc_hd__dfrtp_1 _25926_ (.CLK(clknet_leaf_1_clk),
    .D(net9197),
    .RESET_B(net8413),
    .Q(\pid_d.prev_int[6] ));
 sky130_fd_sc_hd__dfrtp_1 _25927_ (.CLK(clknet_leaf_1_clk),
    .D(_00800_),
    .RESET_B(net8574),
    .Q(\pid_d.prev_int[7] ));
 sky130_fd_sc_hd__dfrtp_1 _25928_ (.CLK(clknet_leaf_2_clk),
    .D(_00801_),
    .RESET_B(net8574),
    .Q(\pid_d.prev_int[8] ));
 sky130_fd_sc_hd__dfrtp_1 _25929_ (.CLK(clknet_leaf_2_clk),
    .D(_00802_),
    .RESET_B(net8574),
    .Q(\pid_d.prev_int[9] ));
 sky130_fd_sc_hd__dfrtp_1 _25930_ (.CLK(clknet_leaf_26_clk),
    .D(net9170),
    .RESET_B(net8573),
    .Q(\pid_d.prev_int[10] ));
 sky130_fd_sc_hd__dfrtp_1 _25931_ (.CLK(clknet_leaf_26_clk),
    .D(_00804_),
    .RESET_B(net8577),
    .Q(\pid_d.prev_int[11] ));
 sky130_fd_sc_hd__dfrtp_1 _25932_ (.CLK(clknet_leaf_25_clk),
    .D(_00805_),
    .RESET_B(net8579),
    .Q(\pid_d.prev_int[12] ));
 sky130_fd_sc_hd__dfrtp_1 _25933_ (.CLK(clknet_leaf_25_clk),
    .D(_00806_),
    .RESET_B(net8591),
    .Q(\pid_d.prev_int[13] ));
 sky130_fd_sc_hd__dfrtp_1 _25934_ (.CLK(clknet_leaf_25_clk),
    .D(_00807_),
    .RESET_B(net8583),
    .Q(\pid_d.prev_int[14] ));
 sky130_fd_sc_hd__dfrtp_1 _25935_ (.CLK(clknet_leaf_24_clk),
    .D(_00808_),
    .RESET_B(net8589),
    .Q(\pid_d.prev_int[15] ));
 sky130_fd_sc_hd__dfstp_1 _25936_ (.CLK(clknet_4_7__leaf_clk),
    .D(_00015_),
    .SET_B(net8581),
    .Q(\pid_d.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _25937_ (.CLK(clknet_leaf_25_clk),
    .D(_00002_),
    .RESET_B(net8581),
    .Q(\pid_d.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _25938_ (.CLK(clknet_4_4__leaf_clk),
    .D(net2997),
    .RESET_B(net8556),
    .Q(\pid_d.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _25939_ (.CLK(clknet_leaf_24_clk),
    .D(_00004_),
    .RESET_B(net8588),
    .Q(\pid_d.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _25940_ (.CLK(clknet_leaf_25_clk),
    .D(_00005_),
    .RESET_B(net8581),
    .Q(\pid_d.state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _25941_ (.CLK(clknet_leaf_120_clk),
    .D(net2379),
    .RESET_B(net8419),
    .Q(\pid_d.state[5] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Right_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Right_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Right_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Right_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Right_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Right_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Right_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Right_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Right_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Right_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Right_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Right_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Right_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Right_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Right_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Right_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Right_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Right_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Right_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Right_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Right_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Right_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Right_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Left_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Left_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Left_365 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Left_366 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Left_367 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Left_368 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Left_369 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Left_370 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Left_371 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Left_372 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Left_373 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Left_374 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Left_375 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Left_376 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Left_377 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Left_378 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Left_379 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Left_380 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Left_381 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Left_382 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Left_383 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Left_384 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Left_385 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Left_386 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Left_387 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Left_388 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Left_389 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Left_390 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Left_391 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Left_392 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Left_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4472 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(angle_in[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(angle_in[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(angle_in[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(angle_in[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(angle_in[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(angle_in[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(angle_in[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(angle_in[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(angle_in[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(angle_in[3]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(angle_in[4]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(angle_in[5]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(angle_in[6]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(angle_in[7]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(angle_in[8]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(angle_in[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(currA_in[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(currA_in[10]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(currA_in[11]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(currA_in[12]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(currA_in[13]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(currA_in[14]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(currA_in[15]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(currA_in[1]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(currA_in[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(currA_in[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(currA_in[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(currA_in[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(currA_in[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(currA_in[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(currA_in[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(currA_in[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(currB_in[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(currB_in[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(currB_in[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(currB_in[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(currB_in[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(currB_in[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(currB_in[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(currB_in[1]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(currB_in[2]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(currB_in[3]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(currB_in[4]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(currB_in[5]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(currB_in[6]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(currB_in[7]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(currB_in[8]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(currB_in[9]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(currT_in[0]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(currT_in[10]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(currT_in[11]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(currT_in[12]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(currT_in[13]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(currT_in[14]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(currT_in[15]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(currT_in[1]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(currT_in[2]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(currT_in[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(currT_in[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(currT_in[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(currT_in[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(currT_in[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(currT_in[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(currT_in[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(periodTop[0]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(periodTop[10]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(periodTop[11]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(periodTop[12]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(periodTop[13]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(periodTop[14]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(periodTop[15]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(periodTop[1]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(periodTop[2]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(periodTop[3]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(periodTop[4]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(periodTop[5]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(periodTop[6]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(periodTop[7]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(periodTop[8]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(periodTop[9]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(pid_d_addr[0]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(pid_d_addr[10]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(pid_d_addr[11]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(pid_d_addr[12]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(pid_d_addr[13]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(pid_d_addr[14]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(pid_d_addr[15]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(pid_d_addr[1]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(pid_d_addr[2]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(pid_d_addr[3]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(pid_d_addr[4]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(pid_d_addr[5]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(pid_d_addr[6]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(pid_d_addr[7]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(pid_d_addr[8]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(pid_d_addr[9]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(pid_d_data[0]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(pid_d_data[10]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(pid_d_data[11]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(pid_d_data[12]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(pid_d_data[13]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(pid_d_data[14]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(pid_d_data[15]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(pid_d_data[1]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(pid_d_data[2]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(pid_d_data[3]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(pid_d_data[4]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(pid_d_data[5]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(pid_d_data[6]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input110 (.A(pid_d_data[7]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(pid_d_data[8]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(pid_d_data[9]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(pid_d_wen),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(pid_q_addr[0]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(pid_q_addr[10]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(pid_q_addr[11]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 input117 (.A(pid_q_addr[12]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(pid_q_addr[13]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(pid_q_addr[14]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(pid_q_addr[15]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(pid_q_addr[1]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(pid_q_addr[2]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(pid_q_addr[3]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(pid_q_addr[4]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(pid_q_addr[5]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(pid_q_addr[6]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(pid_q_addr[7]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(pid_q_addr[8]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(pid_q_addr[9]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(pid_q_data[0]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(pid_q_data[10]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(pid_q_data[11]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(pid_q_data[12]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(pid_q_data[13]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(pid_q_data[14]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(pid_q_data[15]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(pid_q_data[1]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(pid_q_data[2]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(pid_q_data[3]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(pid_q_data[4]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(pid_q_data[5]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 input142 (.A(pid_q_data[6]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(pid_q_data[7]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(pid_q_data[8]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 input145 (.A(pid_q_data[9]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 input146 (.A(pid_q_wen),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 input147 (.A(rstb),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(valid),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_4 output149 (.A(net6682),
    .X(pwmA_out));
 sky130_fd_sc_hd__clkbuf_4 output150 (.A(net150),
    .X(pwmB_out));
 sky130_fd_sc_hd__clkbuf_4 output151 (.A(net6683),
    .X(pwmC_out));
 sky130_fd_sc_hd__clkbuf_4 output152 (.A(net8075),
    .X(ready));
 sky130_fd_sc_hd__buf_1 wire153 (.A(_06495_),
    .X(net153));
 sky130_fd_sc_hd__buf_1 wire154 (.A(_06489_),
    .X(net154));
 sky130_fd_sc_hd__buf_1 wire155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__buf_1 wire156 (.A(_06479_),
    .X(net156));
 sky130_fd_sc_hd__buf_1 wire157 (.A(_06431_),
    .X(net157));
 sky130_fd_sc_hd__buf_1 wire158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 wire159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__buf_1 wire160 (.A(_06462_),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 wire161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 wire162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 wire163 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 wire164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 wire165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 wire166 (.A(_08634_),
    .X(net166));
 sky130_fd_sc_hd__buf_1 wire167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 wire168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 wire169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 wire170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 wire171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 wire172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 wire173 (.A(_08592_),
    .X(net173));
 sky130_fd_sc_hd__buf_1 wire174 (.A(_06399_),
    .X(net174));
 sky130_fd_sc_hd__buf_1 wire175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 wire176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 wire177 (.A(_04640_),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 wire178 (.A(_02618_),
    .X(net178));
 sky130_fd_sc_hd__buf_1 wire179 (.A(_12027_),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 wire180 (.A(_10616_),
    .X(net180));
 sky130_fd_sc_hd__buf_1 wire181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 wire182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 wire183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 wire184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 wire185 (.A(net186),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 wire186 (.A(_08545_),
    .X(net186));
 sky130_fd_sc_hd__buf_1 wire187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__buf_1 wire188 (.A(_06363_),
    .X(net188));
 sky130_fd_sc_hd__buf_1 wire189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__buf_1 wire190 (.A(_06270_),
    .X(net190));
 sky130_fd_sc_hd__buf_1 wire191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__buf_1 wire192 (.A(_06152_),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 wire193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 wire194 (.A(_04814_),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 wire195 (.A(_04505_),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 wire196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 wire197 (.A(_04501_),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 wire198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 wire199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__buf_1 wire200 (.A(_04382_),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 wire201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 wire202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 wire203 (.A(_02842_),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 wire204 (.A(_02516_),
    .X(net204));
 sky130_fd_sc_hd__buf_1 wire205 (.A(_02459_),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 wire206 (.A(_02407_),
    .X(net206));
 sky130_fd_sc_hd__buf_1 wire207 (.A(_10780_),
    .X(net207));
 sky130_fd_sc_hd__buf_1 wire208 (.A(_08496_),
    .X(net208));
 sky130_fd_sc_hd__buf_1 wire209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_1 wire210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_1 wire211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 wire212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 wire213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 wire214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 wire215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_1 wire216 (.A(_08489_),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 wire217 (.A(_06364_),
    .X(net217));
 sky130_fd_sc_hd__buf_1 max_length218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__buf_1 wire219 (.A(_06321_),
    .X(net219));
 sky130_fd_sc_hd__buf_1 wire220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__buf_1 wire221 (.A(net222),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_1 wire222 (.A(_06216_),
    .X(net222));
 sky130_fd_sc_hd__buf_1 wire223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__buf_1 wire224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_1 wire225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 wire226 (.A(_06011_),
    .X(net226));
 sky130_fd_sc_hd__buf_1 wire227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 wire228 (.A(net229),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_1 wire229 (.A(_04632_),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 wire230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__buf_1 wire231 (.A(_04453_),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_1 wire232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 wire233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__buf_1 wire234 (.A(_04445_),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 wire235 (.A(net236),
    .X(net235));
 sky130_fd_sc_hd__buf_1 wire236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_1 wire237 (.A(_04320_),
    .X(net237));
 sky130_fd_sc_hd__buf_1 wire238 (.A(_04170_),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 wire239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 wire240 (.A(net241),
    .X(net240));
 sky130_fd_sc_hd__buf_1 wire241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_1 wire242 (.A(_04028_),
    .X(net242));
 sky130_fd_sc_hd__buf_1 wire243 (.A(_12014_),
    .X(net243));
 sky130_fd_sc_hd__buf_1 wire244 (.A(_11987_),
    .X(net244));
 sky130_fd_sc_hd__buf_1 wire245 (.A(_10766_),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_1 wire246 (.A(_10511_),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_1 wire247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_1 wire248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 wire249 (.A(net250),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 wire250 (.A(net251),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 wire251 (.A(net252),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 wire252 (.A(net253),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_1 wire253 (.A(_08370_),
    .X(net253));
 sky130_fd_sc_hd__buf_1 wire254 (.A(_06361_),
    .X(net254));
 sky130_fd_sc_hd__buf_1 wire255 (.A(_06360_),
    .X(net255));
 sky130_fd_sc_hd__buf_1 wire256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_1 wire257 (.A(_06086_),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_1 wire258 (.A(_04656_),
    .X(net258));
 sky130_fd_sc_hd__buf_1 wire259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 wire260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 wire261 (.A(net262),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 wire262 (.A(_04624_),
    .X(net262));
 sky130_fd_sc_hd__buf_1 wire263 (.A(_04402_),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_1 wire264 (.A(_04388_),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_1 max_length265 (.A(_04388_),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 wire266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_1 wire267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_1 max_length268 (.A(net269),
    .X(net268));
 sky130_fd_sc_hd__buf_1 wire269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_1 wire270 (.A(_04108_),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_1 wire271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__buf_1 wire272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 wire273 (.A(_02390_),
    .X(net273));
 sky130_fd_sc_hd__buf_1 wire274 (.A(_11958_),
    .X(net274));
 sky130_fd_sc_hd__buf_1 wire275 (.A(_10746_),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_1 wire276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_1 wire277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_1 wire278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 wire279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 wire280 (.A(_08432_),
    .X(net280));
 sky130_fd_sc_hd__buf_1 wire281 (.A(_06760_),
    .X(net281));
 sky130_fd_sc_hd__buf_1 wire282 (.A(_06275_),
    .X(net282));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire283 (.A(_06020_),
    .X(net283));
 sky130_fd_sc_hd__buf_1 wire284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__buf_1 wire285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_1 wire286 (.A(_05936_),
    .X(net286));
 sky130_fd_sc_hd__buf_1 wire287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__buf_1 wire288 (.A(net289),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_1 wire289 (.A(_05856_),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_1 wire290 (.A(_04327_),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_1 wire291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__buf_1 wire292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_1 wire293 (.A(_04250_),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_1 wire294 (.A(_02614_),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 wire295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_1 wire296 (.A(net297),
    .X(net296));
 sky130_fd_sc_hd__buf_1 wire297 (.A(_02327_),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_1 wire298 (.A(net299),
    .X(net298));
 sky130_fd_sc_hd__buf_1 wire299 (.A(net300),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_1 wire300 (.A(net301),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_1 wire301 (.A(_02253_),
    .X(net301));
 sky130_fd_sc_hd__buf_1 wire302 (.A(_10728_),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_2 wire303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 wire304 (.A(_08377_),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_1 wire305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 wire306 (.A(net307),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 wire307 (.A(net308),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_1 wire308 (.A(net309),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_1 wire309 (.A(net310),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_1 wire310 (.A(_08305_),
    .X(net310));
 sky130_fd_sc_hd__buf_1 wire311 (.A(net312),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_1 wire312 (.A(net313),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_1 wire313 (.A(net314),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_1 wire314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_1 wire315 (.A(net316),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_1 wire316 (.A(net317),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_1 wire317 (.A(_08236_),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_1 wire318 (.A(_06757_),
    .X(net318));
 sky130_fd_sc_hd__buf_1 wire319 (.A(_06276_),
    .X(net319));
 sky130_fd_sc_hd__buf_1 wire320 (.A(_06019_),
    .X(net320));
 sky130_fd_sc_hd__buf_1 wire321 (.A(_06016_),
    .X(net321));
 sky130_fd_sc_hd__buf_1 wire322 (.A(_05862_),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 max_length323 (.A(net324),
    .X(net323));
 sky130_fd_sc_hd__buf_1 wire324 (.A(net325),
    .X(net324));
 sky130_fd_sc_hd__buf_1 wire325 (.A(net326),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_1 wire326 (.A(_05775_),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_1 wire327 (.A(_04655_),
    .X(net327));
 sky130_fd_sc_hd__buf_1 wire328 (.A(_04384_),
    .X(net328));
 sky130_fd_sc_hd__buf_1 wire329 (.A(net330),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_1 wire330 (.A(_03945_),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 wire331 (.A(net332),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_1 wire332 (.A(net333),
    .X(net332));
 sky130_fd_sc_hd__buf_1 wire333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_1 wire334 (.A(net335),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_1 wire335 (.A(_03851_),
    .X(net335));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire336 (.A(_02277_),
    .X(net336));
 sky130_fd_sc_hd__buf_1 wire337 (.A(_02260_),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_1 wire338 (.A(net339),
    .X(net338));
 sky130_fd_sc_hd__buf_1 wire339 (.A(net340),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_1 wire340 (.A(net341),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_1 wire341 (.A(_02172_),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_1 wire342 (.A(net343),
    .X(net342));
 sky130_fd_sc_hd__buf_1 wire343 (.A(net344),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_1 wire344 (.A(net345),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_1 wire345 (.A(_02099_),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_1 wire346 (.A(net347),
    .X(net346));
 sky130_fd_sc_hd__buf_1 wire347 (.A(net348),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_1 wire348 (.A(net349),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_1 wire349 (.A(_02007_),
    .X(net349));
 sky130_fd_sc_hd__buf_1 max_length350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__buf_1 wire351 (.A(_11735_),
    .X(net351));
 sky130_fd_sc_hd__buf_1 wire352 (.A(_10693_),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_1 wire353 (.A(_08732_),
    .X(net353));
 sky130_fd_sc_hd__buf_1 wire354 (.A(net355),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_1 wire355 (.A(net356),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_1 wire356 (.A(net357),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_1 wire357 (.A(net358),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_1 wire358 (.A(_08161_),
    .X(net358));
 sky130_fd_sc_hd__buf_1 wire359 (.A(net360),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_1 wire360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_1 wire361 (.A(net362),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_1 wire362 (.A(net363),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_1 wire363 (.A(net364),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_1 wire364 (.A(net365),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_1 wire365 (.A(_08086_),
    .X(net365));
 sky130_fd_sc_hd__buf_1 wire366 (.A(_06319_),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_2 wire367 (.A(net368),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 wire368 (.A(net369),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_1 wire369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 wire370 (.A(net371),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_1 wire371 (.A(_05681_),
    .X(net371));
 sky130_fd_sc_hd__buf_1 wire372 (.A(net373),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_1 wire373 (.A(_04617_),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_1 wire374 (.A(net375),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_1 max_length375 (.A(_04257_),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_2 wire376 (.A(net377),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_1 wire377 (.A(net378),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_1 wire378 (.A(net379),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_1 wire379 (.A(_03866_),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_1 wire380 (.A(_02513_),
    .X(net380));
 sky130_fd_sc_hd__buf_1 wire381 (.A(_02272_),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_1 wire382 (.A(_10402_),
    .X(net382));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire383 (.A(net384),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_1 wire384 (.A(_08730_),
    .X(net384));
 sky130_fd_sc_hd__buf_1 wire385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__buf_1 wire386 (.A(net387),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_1 wire387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_1 wire388 (.A(_08090_),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_1 wire389 (.A(net390),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_1 wire390 (.A(net391),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_1 wire391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_1 wire392 (.A(net393),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_1 wire393 (.A(net394),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_1 wire394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_1 wire395 (.A(_08010_),
    .X(net395));
 sky130_fd_sc_hd__buf_1 wire396 (.A(net397),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_1 wire397 (.A(net398),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_1 wire398 (.A(net399),
    .X(net398));
 sky130_fd_sc_hd__buf_1 wire399 (.A(net400),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_1 wire400 (.A(net401),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_1 wire401 (.A(net402),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_1 wire402 (.A(_07922_),
    .X(net402));
 sky130_fd_sc_hd__buf_1 wire403 (.A(_06365_),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_2 wire404 (.A(_06002_),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_1 wire405 (.A(net406),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_1 wire406 (.A(net407),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_1 max_length407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__buf_1 wire408 (.A(net409),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_1 wire409 (.A(_03761_),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_1 wire410 (.A(net411),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_1 max_length411 (.A(_02180_),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_1 wire412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__buf_1 wire413 (.A(net414),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_1 wire414 (.A(_01907_),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_1 wire415 (.A(net416),
    .X(net415));
 sky130_fd_sc_hd__buf_1 wire416 (.A(net417),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_1 wire417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_1 wire418 (.A(net419),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_1 wire419 (.A(_01533_),
    .X(net419));
 sky130_fd_sc_hd__buf_1 wire420 (.A(_11926_),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_2 wire421 (.A(_10518_),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_2 max_length422 (.A(_10407_),
    .X(net422));
 sky130_fd_sc_hd__buf_1 wire423 (.A(_08726_),
    .X(net423));
 sky130_fd_sc_hd__buf_1 wire424 (.A(_08240_),
    .X(net424));
 sky130_fd_sc_hd__buf_1 wire425 (.A(_07924_),
    .X(net425));
 sky130_fd_sc_hd__buf_1 wire426 (.A(net427),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_1 wire427 (.A(net428),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_1 wire428 (.A(net429),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_1 wire429 (.A(net430),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_1 wire430 (.A(net431),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_1 wire431 (.A(net432),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_1 wire432 (.A(_07829_),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_1 wire433 (.A(net434),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_1 wire434 (.A(net435),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_1 wire435 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_1 wire436 (.A(net437),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_1 wire437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_1 wire438 (.A(net439),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_1 wire439 (.A(_07740_),
    .X(net439));
 sky130_fd_sc_hd__buf_1 wire440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_1 wire441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_1 wire442 (.A(net443),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_1 wire443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_1 wire444 (.A(net445),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_1 wire445 (.A(net446),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_1 wire446 (.A(net447),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_1 wire447 (.A(_07640_),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_1 wire448 (.A(_06736_),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_2 wire449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_1 wire450 (.A(_06021_),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_2 wire451 (.A(_05933_),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_1 wire452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_1 wire453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_1 wire454 (.A(_05334_),
    .X(net454));
 sky130_fd_sc_hd__buf_1 wire455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_1 wire456 (.A(_04611_),
    .X(net456));
 sky130_fd_sc_hd__buf_1 wire457 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_1 wire458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_1 wire459 (.A(_04603_),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_1 wire460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_1 max_length461 (.A(_04184_),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_1 wire462 (.A(net463),
    .X(net462));
 sky130_fd_sc_hd__buf_1 wire463 (.A(net464),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_1 wire464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_1 wire465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_1 wire466 (.A(_03660_),
    .X(net466));
 sky130_fd_sc_hd__buf_1 wire467 (.A(net468),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_1 wire468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__clkbuf_1 wire469 (.A(net470),
    .X(net469));
 sky130_fd_sc_hd__clkbuf_1 wire470 (.A(_03566_),
    .X(net470));
 sky130_fd_sc_hd__buf_1 wire471 (.A(_01925_),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_1 wire472 (.A(net473),
    .X(net472));
 sky130_fd_sc_hd__buf_1 wire473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_1 wire474 (.A(_01809_),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_1 wire475 (.A(net476),
    .X(net475));
 sky130_fd_sc_hd__buf_1 wire476 (.A(net477),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_1 wire477 (.A(_01635_),
    .X(net477));
 sky130_fd_sc_hd__buf_1 wire478 (.A(_01532_),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_1 wire479 (.A(net480),
    .X(net479));
 sky130_fd_sc_hd__buf_1 wire480 (.A(net481),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_1 wire481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_1 wire482 (.A(net483),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_1 wire483 (.A(net484),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_1 wire484 (.A(net485),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_1 wire485 (.A(net486),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_1 wire486 (.A(_01242_),
    .X(net486));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire487 (.A(_11742_),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_1 wire488 (.A(_11619_),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_1 wire489 (.A(_10341_),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_2 wire490 (.A(_08378_),
    .X(net490));
 sky130_fd_sc_hd__buf_1 wire491 (.A(_08243_),
    .X(net491));
 sky130_fd_sc_hd__buf_1 wire492 (.A(_08234_),
    .X(net492));
 sky130_fd_sc_hd__buf_1 wire493 (.A(_08160_),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_1 wire494 (.A(net495),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_1 wire495 (.A(net496),
    .X(net495));
 sky130_fd_sc_hd__clkbuf_1 wire496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_1 wire497 (.A(net498),
    .X(net497));
 sky130_fd_sc_hd__clkbuf_1 wire498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_1 wire499 (.A(net500),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_1 wire500 (.A(net501),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_1 wire501 (.A(net502),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_1 wire502 (.A(_07559_),
    .X(net502));
 sky130_fd_sc_hd__buf_1 wire503 (.A(_05998_),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_2 wire504 (.A(net505),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_1 wire505 (.A(net506),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_1 wire506 (.A(net507),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_1 wire507 (.A(_05683_),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_1 wire508 (.A(_04653_),
    .X(net508));
 sky130_fd_sc_hd__buf_1 wire509 (.A(_04497_),
    .X(net509));
 sky130_fd_sc_hd__buf_1 wire510 (.A(_04177_),
    .X(net510));
 sky130_fd_sc_hd__buf_1 wire511 (.A(_03846_),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_1 wire512 (.A(net513),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_1 wire513 (.A(net514),
    .X(net513));
 sky130_fd_sc_hd__buf_1 wire514 (.A(net515),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_1 wire515 (.A(net516),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_1 wire516 (.A(_03474_),
    .X(net516));
 sky130_fd_sc_hd__buf_1 wire517 (.A(net518),
    .X(net517));
 sky130_fd_sc_hd__clkbuf_1 wire518 (.A(net519),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_1 wire519 (.A(_02512_),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_1 wire520 (.A(net521),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_1 wire521 (.A(_02415_),
    .X(net521));
 sky130_fd_sc_hd__buf_1 wire522 (.A(_02106_),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_1 wire523 (.A(net524),
    .X(net523));
 sky130_fd_sc_hd__buf_1 wire524 (.A(net525),
    .X(net524));
 sky130_fd_sc_hd__clkbuf_1 wire525 (.A(_01727_),
    .X(net525));
 sky130_fd_sc_hd__buf_1 wire526 (.A(_10612_),
    .X(net526));
 sky130_fd_sc_hd__buf_1 wire527 (.A(_09106_),
    .X(net527));
 sky130_fd_sc_hd__buf_1 wire528 (.A(_08720_),
    .X(net528));
 sky130_fd_sc_hd__buf_1 wire529 (.A(_06258_),
    .X(net529));
 sky130_fd_sc_hd__buf_1 wire530 (.A(_06088_),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_1 wire531 (.A(_06077_),
    .X(net531));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire532 (.A(_06075_),
    .X(net532));
 sky130_fd_sc_hd__buf_1 wire533 (.A(_05847_),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_2 wire534 (.A(_05762_),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_1 wire535 (.A(_05240_),
    .X(net535));
 sky130_fd_sc_hd__clkbuf_1 wire536 (.A(net537),
    .X(net536));
 sky130_fd_sc_hd__clkbuf_1 wire537 (.A(_04115_),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_1 wire538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_1 wire539 (.A(net540),
    .X(net539));
 sky130_fd_sc_hd__buf_1 wire540 (.A(net541),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_1 wire541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_1 wire542 (.A(_03384_),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_1 wire543 (.A(net544),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_1 wire544 (.A(net545),
    .X(net544));
 sky130_fd_sc_hd__buf_1 wire545 (.A(net546),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_1 wire546 (.A(net547),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_1 wire547 (.A(net548),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_1 wire548 (.A(_03310_),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_2 wire549 (.A(net550),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_1 wire550 (.A(_02385_),
    .X(net550));
 sky130_fd_sc_hd__buf_1 wire551 (.A(_02339_),
    .X(net551));
 sky130_fd_sc_hd__buf_1 wire552 (.A(_02323_),
    .X(net552));
 sky130_fd_sc_hd__clkbuf_1 wire553 (.A(net554),
    .X(net553));
 sky130_fd_sc_hd__clkbuf_1 wire554 (.A(net555),
    .X(net554));
 sky130_fd_sc_hd__buf_1 wire555 (.A(net556),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_1 wire556 (.A(net557),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_1 wire557 (.A(net558),
    .X(net557));
 sky130_fd_sc_hd__clkbuf_1 wire558 (.A(net559),
    .X(net558));
 sky130_fd_sc_hd__clkbuf_1 wire559 (.A(_01426_),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_1 wire560 (.A(net561),
    .X(net560));
 sky130_fd_sc_hd__buf_1 wire561 (.A(net562),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_1 wire562 (.A(net563),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_1 wire563 (.A(net564),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_1 wire564 (.A(net565),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_1 wire565 (.A(net566),
    .X(net565));
 sky130_fd_sc_hd__clkbuf_1 wire566 (.A(_01331_),
    .X(net566));
 sky130_fd_sc_hd__buf_1 wire567 (.A(_11666_),
    .X(net567));
 sky130_fd_sc_hd__buf_1 wire568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire569 (.A(net570),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_1 wire570 (.A(_11485_),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_2 wire571 (.A(_08380_),
    .X(net571));
 sky130_fd_sc_hd__buf_1 wire572 (.A(net573),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_1 wire573 (.A(_08093_),
    .X(net573));
 sky130_fd_sc_hd__buf_1 wire574 (.A(net575),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_1 wire575 (.A(net576),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_1 wire576 (.A(_07556_),
    .X(net576));
 sky130_fd_sc_hd__buf_1 wire577 (.A(_05835_),
    .X(net577));
 sky130_fd_sc_hd__buf_1 wire578 (.A(net579),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_1 wire579 (.A(net580),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_1 wire580 (.A(_05769_),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_2 wire581 (.A(net582),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_1 wire582 (.A(_05666_),
    .X(net582));
 sky130_fd_sc_hd__buf_1 wire583 (.A(net584),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_1 wire584 (.A(net585),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_1 max_length585 (.A(_05317_),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_1 wire586 (.A(_04652_),
    .X(net586));
 sky130_fd_sc_hd__buf_1 wire587 (.A(_04248_),
    .X(net587));
 sky130_fd_sc_hd__buf_1 wire588 (.A(_04246_),
    .X(net588));
 sky130_fd_sc_hd__buf_1 wire589 (.A(_04104_),
    .X(net589));
 sky130_fd_sc_hd__buf_1 wire590 (.A(net591),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_1 wire591 (.A(_04025_),
    .X(net591));
 sky130_fd_sc_hd__buf_1 wire592 (.A(net593),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_1 wire593 (.A(net594),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_1 wire594 (.A(_03940_),
    .X(net594));
 sky130_fd_sc_hd__buf_1 wire595 (.A(net596),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_1 wire596 (.A(_03939_),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_1 wire597 (.A(net598),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_1 wire598 (.A(_02454_),
    .X(net598));
 sky130_fd_sc_hd__buf_1 wire599 (.A(_01903_),
    .X(net599));
 sky130_fd_sc_hd__buf_1 wire600 (.A(net601),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_1 wire601 (.A(net602),
    .X(net601));
 sky130_fd_sc_hd__clkbuf_1 wire602 (.A(_01552_),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_1 wire603 (.A(_12186_),
    .X(net603));
 sky130_fd_sc_hd__buf_2 wire604 (.A(_11548_),
    .X(net604));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire605 (.A(_10413_),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_1 wire606 (.A(net607),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_2 wire607 (.A(net608),
    .X(net607));
 sky130_fd_sc_hd__clkbuf_1 wire608 (.A(net609),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_1 wire609 (.A(net610),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_1 wire610 (.A(_10260_),
    .X(net610));
 sky130_fd_sc_hd__buf_1 wire611 (.A(net613),
    .X(net611));
 sky130_fd_sc_hd__buf_1 wire612 (.A(_09282_),
    .X(net612));
 sky130_fd_sc_hd__buf_1 max_length613 (.A(_09282_),
    .X(net613));
 sky130_fd_sc_hd__buf_1 wire614 (.A(_09276_),
    .X(net614));
 sky130_fd_sc_hd__buf_1 wire615 (.A(net616),
    .X(net615));
 sky130_fd_sc_hd__buf_1 max_length616 (.A(_09276_),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_2 wire617 (.A(_09135_),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_2 wire618 (.A(_09125_),
    .X(net618));
 sky130_fd_sc_hd__buf_1 wire619 (.A(net620),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_1 wire620 (.A(_08714_),
    .X(net620));
 sky130_fd_sc_hd__buf_1 wire621 (.A(_05937_),
    .X(net621));
 sky130_fd_sc_hd__buf_1 wire622 (.A(net623),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_1 wire623 (.A(net624),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_1 wire624 (.A(_05760_),
    .X(net624));
 sky130_fd_sc_hd__buf_1 wire625 (.A(net626),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_1 wire626 (.A(net627),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_1 wire627 (.A(_05685_),
    .X(net627));
 sky130_fd_sc_hd__buf_1 wire628 (.A(_05635_),
    .X(net628));
 sky130_fd_sc_hd__buf_1 wire629 (.A(net630),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_1 wire630 (.A(_04595_),
    .X(net630));
 sky130_fd_sc_hd__buf_1 wire631 (.A(net632),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_1 wire632 (.A(_04443_),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_2 wire633 (.A(_04167_),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_2 wire634 (.A(net635),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_1 wire635 (.A(_04166_),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_1 wire636 (.A(net637),
    .X(net636));
 sky130_fd_sc_hd__clkbuf_1 wire637 (.A(net638),
    .X(net637));
 sky130_fd_sc_hd__clkbuf_1 max_length638 (.A(_04035_),
    .X(net638));
 sky130_fd_sc_hd__buf_1 wire639 (.A(_03488_),
    .X(net639));
 sky130_fd_sc_hd__buf_1 wire640 (.A(net641),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_1 wire641 (.A(net642),
    .X(net641));
 sky130_fd_sc_hd__clkbuf_1 wire642 (.A(net643),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_1 wire643 (.A(net644),
    .X(net643));
 sky130_fd_sc_hd__clkbuf_1 wire644 (.A(net645),
    .X(net644));
 sky130_fd_sc_hd__clkbuf_1 wire645 (.A(_03238_),
    .X(net645));
 sky130_fd_sc_hd__buf_1 wire646 (.A(net647),
    .X(net646));
 sky130_fd_sc_hd__clkbuf_1 wire647 (.A(net648),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_1 wire648 (.A(net649),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_1 wire649 (.A(net650),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_1 wire650 (.A(net651),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_1 wire651 (.A(_03181_),
    .X(net651));
 sky130_fd_sc_hd__clkbuf_1 wire652 (.A(_01549_),
    .X(net652));
 sky130_fd_sc_hd__buf_1 wire653 (.A(net654),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_1 wire654 (.A(net655),
    .X(net654));
 sky130_fd_sc_hd__clkbuf_1 wire655 (.A(net656),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_1 wire656 (.A(_11368_),
    .X(net656));
 sky130_fd_sc_hd__buf_1 wire657 (.A(_10702_),
    .X(net657));
 sky130_fd_sc_hd__buf_1 wire658 (.A(_10692_),
    .X(net658));
 sky130_fd_sc_hd__buf_1 wire659 (.A(net660),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_1 wire660 (.A(net661),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_1 wire661 (.A(net662),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_1 wire662 (.A(_10267_),
    .X(net662));
 sky130_fd_sc_hd__buf_1 wire663 (.A(net664),
    .X(net663));
 sky130_fd_sc_hd__clkbuf_1 wire664 (.A(net665),
    .X(net664));
 sky130_fd_sc_hd__clkbuf_1 wire665 (.A(net666),
    .X(net665));
 sky130_fd_sc_hd__clkbuf_1 wire666 (.A(_10266_),
    .X(net666));
 sky130_fd_sc_hd__buf_1 wire667 (.A(net668),
    .X(net667));
 sky130_fd_sc_hd__buf_1 wire668 (.A(_09273_),
    .X(net668));
 sky130_fd_sc_hd__buf_1 wire669 (.A(_09270_),
    .X(net669));
 sky130_fd_sc_hd__buf_1 wire670 (.A(_09116_),
    .X(net670));
 sky130_fd_sc_hd__clkbuf_1 wire671 (.A(_08536_),
    .X(net671));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire672 (.A(_08210_),
    .X(net672));
 sky130_fd_sc_hd__buf_1 wire673 (.A(_08075_),
    .X(net673));
 sky130_fd_sc_hd__buf_1 wire674 (.A(_07562_),
    .X(net674));
 sky130_fd_sc_hd__buf_1 wire675 (.A(_07555_),
    .X(net675));
 sky130_fd_sc_hd__clkbuf_1 wire676 (.A(_06707_),
    .X(net676));
 sky130_fd_sc_hd__buf_1 wire677 (.A(_06204_),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_1 wire678 (.A(_06079_),
    .X(net678));
 sky130_fd_sc_hd__buf_1 wire679 (.A(net680),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_1 wire680 (.A(_05836_),
    .X(net680));
 sky130_fd_sc_hd__buf_1 wire681 (.A(_05808_),
    .X(net681));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire682 (.A(_05470_),
    .X(net682));
 sky130_fd_sc_hd__clkbuf_2 wire683 (.A(_05337_),
    .X(net683));
 sky130_fd_sc_hd__buf_1 wire684 (.A(_05305_),
    .X(net684));
 sky130_fd_sc_hd__buf_1 wire685 (.A(_04801_),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_1 wire686 (.A(net687),
    .X(net686));
 sky130_fd_sc_hd__clkbuf_1 wire687 (.A(_04651_),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_1 wire688 (.A(net689),
    .X(net688));
 sky130_fd_sc_hd__clkbuf_1 wire689 (.A(_04650_),
    .X(net689));
 sky130_fd_sc_hd__buf_1 wire690 (.A(net691),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_1 wire691 (.A(_04591_),
    .X(net691));
 sky130_fd_sc_hd__buf_1 wire692 (.A(net693),
    .X(net692));
 sky130_fd_sc_hd__clkbuf_1 wire693 (.A(_04050_),
    .X(net693));
 sky130_fd_sc_hd__buf_1 wire694 (.A(net695),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_1 wire695 (.A(_04016_),
    .X(net695));
 sky130_fd_sc_hd__buf_1 wire696 (.A(_03468_),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_1 wire697 (.A(_03174_),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_1 wire698 (.A(_01921_),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_1 wire699 (.A(_01914_),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_1 max_length700 (.A(_01914_),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_1 wire701 (.A(_01630_),
    .X(net701));
 sky130_fd_sc_hd__buf_1 wire702 (.A(_01521_),
    .X(net702));
 sky130_fd_sc_hd__buf_1 wire703 (.A(net704),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_1 wire704 (.A(_01252_),
    .X(net704));
 sky130_fd_sc_hd__clkbuf_1 wire705 (.A(net706),
    .X(net705));
 sky130_fd_sc_hd__clkbuf_1 wire706 (.A(_01251_),
    .X(net706));
 sky130_fd_sc_hd__clkbuf_1 wire707 (.A(_12393_),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_2 wire708 (.A(_11669_),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_1 wire709 (.A(net710),
    .X(net709));
 sky130_fd_sc_hd__clkbuf_1 wire710 (.A(net711),
    .X(net710));
 sky130_fd_sc_hd__clkbuf_1 wire711 (.A(_11367_),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_1 wire712 (.A(_11252_),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_1 wire713 (.A(_11118_),
    .X(net713));
 sky130_fd_sc_hd__buf_2 wire714 (.A(_10409_),
    .X(net714));
 sky130_fd_sc_hd__buf_1 wire715 (.A(_10152_),
    .X(net715));
 sky130_fd_sc_hd__buf_1 wire716 (.A(net717),
    .X(net716));
 sky130_fd_sc_hd__clkbuf_1 wire717 (.A(net718),
    .X(net717));
 sky130_fd_sc_hd__clkbuf_1 wire718 (.A(net719),
    .X(net718));
 sky130_fd_sc_hd__clkbuf_1 wire719 (.A(_10023_),
    .X(net719));
 sky130_fd_sc_hd__buf_1 wire720 (.A(net721),
    .X(net720));
 sky130_fd_sc_hd__clkbuf_1 wire721 (.A(net722),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_1 wire722 (.A(_08708_),
    .X(net722));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire723 (.A(_08435_),
    .X(net723));
 sky130_fd_sc_hd__buf_1 wire724 (.A(_08355_),
    .X(net724));
 sky130_fd_sc_hd__clkbuf_1 wire725 (.A(_07466_),
    .X(net725));
 sky130_fd_sc_hd__buf_1 wire726 (.A(_06702_),
    .X(net726));
 sky130_fd_sc_hd__buf_1 wire727 (.A(_05982_),
    .X(net727));
 sky130_fd_sc_hd__buf_1 wire728 (.A(net729),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_1 wire729 (.A(net730),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_1 wire730 (.A(_05697_),
    .X(net730));
 sky130_fd_sc_hd__buf_1 wire731 (.A(_05605_),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_2 wire732 (.A(_05517_),
    .X(net732));
 sky130_fd_sc_hd__buf_1 wire733 (.A(_05431_),
    .X(net733));
 sky130_fd_sc_hd__buf_1 wire734 (.A(_05397_),
    .X(net734));
 sky130_fd_sc_hd__buf_1 max_cap735 (.A(_05245_),
    .X(net735));
 sky130_fd_sc_hd__buf_1 wire736 (.A(_05123_),
    .X(net736));
 sky130_fd_sc_hd__buf_1 wire737 (.A(_04585_),
    .X(net737));
 sky130_fd_sc_hd__buf_1 wire738 (.A(_04576_),
    .X(net738));
 sky130_fd_sc_hd__buf_1 wire739 (.A(net740),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_1 wire740 (.A(_04018_),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_1 wire741 (.A(net742),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_1 wire742 (.A(_03952_),
    .X(net742));
 sky130_fd_sc_hd__buf_1 wire743 (.A(_03863_),
    .X(net743));
 sky130_fd_sc_hd__buf_1 wire744 (.A(_03561_),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_2 wire745 (.A(net746),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_1 wire746 (.A(net747),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_1 wire747 (.A(net748),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_1 wire748 (.A(_03381_),
    .X(net748));
 sky130_fd_sc_hd__buf_1 wire749 (.A(net750),
    .X(net749));
 sky130_fd_sc_hd__clkbuf_1 wire750 (.A(net751),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_1 wire751 (.A(net752),
    .X(net751));
 sky130_fd_sc_hd__clkbuf_1 wire752 (.A(net753),
    .X(net752));
 sky130_fd_sc_hd__clkbuf_1 wire753 (.A(net754),
    .X(net753));
 sky130_fd_sc_hd__clkbuf_1 wire754 (.A(_03240_),
    .X(net754));
 sky130_fd_sc_hd__buf_1 wire755 (.A(_03180_),
    .X(net755));
 sky130_fd_sc_hd__buf_1 wire756 (.A(_02204_),
    .X(net756));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire757 (.A(_01422_),
    .X(net757));
 sky130_fd_sc_hd__buf_1 wire758 (.A(_01327_),
    .X(net758));
 sky130_fd_sc_hd__buf_1 wire759 (.A(_01250_),
    .X(net759));
 sky130_fd_sc_hd__buf_1 wire760 (.A(_01219_),
    .X(net760));
 sky130_fd_sc_hd__buf_1 wire761 (.A(net762),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_1 wire762 (.A(_01216_),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_1 wire763 (.A(_11117_),
    .X(net763));
 sky130_fd_sc_hd__buf_2 wire764 (.A(_10563_),
    .X(net764));
 sky130_fd_sc_hd__clkbuf_2 wire765 (.A(net766),
    .X(net765));
 sky130_fd_sc_hd__clkbuf_1 wire766 (.A(_10338_),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_1 wire767 (.A(_10256_),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_1 wire768 (.A(_10017_),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_1 wire769 (.A(_09471_),
    .X(net769));
 sky130_fd_sc_hd__buf_1 wire770 (.A(_09378_),
    .X(net770));
 sky130_fd_sc_hd__buf_1 wire771 (.A(_09266_),
    .X(net771));
 sky130_fd_sc_hd__buf_1 wire772 (.A(_09046_),
    .X(net772));
 sky130_fd_sc_hd__buf_1 wire773 (.A(_08426_),
    .X(net773));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire774 (.A(net775),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_1 wire775 (.A(_08169_),
    .X(net775));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire776 (.A(net777),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_1 wire777 (.A(_08111_),
    .X(net777));
 sky130_fd_sc_hd__buf_1 wire778 (.A(_07646_),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_1 wire779 (.A(_07452_),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_2 wire780 (.A(_05985_),
    .X(net780));
 sky130_fd_sc_hd__buf_1 wire781 (.A(_05978_),
    .X(net781));
 sky130_fd_sc_hd__buf_1 wire782 (.A(_05959_),
    .X(net782));
 sky130_fd_sc_hd__buf_1 wire783 (.A(net784),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_1 wire784 (.A(_05844_),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_1 wire785 (.A(net786),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_1 wire786 (.A(net787),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_1 wire787 (.A(net788),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_1 wire788 (.A(_05766_),
    .X(net788));
 sky130_fd_sc_hd__buf_1 wire789 (.A(_05225_),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_2 wire790 (.A(_05205_),
    .X(net790));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire791 (.A(_05141_),
    .X(net791));
 sky130_fd_sc_hd__buf_2 wire792 (.A(_04309_),
    .X(net792));
 sky130_fd_sc_hd__buf_1 wire793 (.A(net794),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_1 wire794 (.A(_04053_),
    .X(net794));
 sky130_fd_sc_hd__buf_1 wire795 (.A(_03781_),
    .X(net795));
 sky130_fd_sc_hd__buf_1 wire796 (.A(net797),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_1 wire797 (.A(net798),
    .X(net797));
 sky130_fd_sc_hd__clkbuf_1 wire798 (.A(net799),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_1 wire799 (.A(_03305_),
    .X(net799));
 sky130_fd_sc_hd__buf_1 wire800 (.A(net801),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_1 wire801 (.A(_02595_),
    .X(net801));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire802 (.A(_02074_),
    .X(net802));
 sky130_fd_sc_hd__clkbuf_1 wire803 (.A(_01823_),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_1 wire804 (.A(_01816_),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_1 max_length805 (.A(_01816_),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_2 wire806 (.A(_01411_),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_1 wire807 (.A(_01215_),
    .X(net807));
 sky130_fd_sc_hd__buf_1 wire808 (.A(_01076_),
    .X(net808));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire809 (.A(net810),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_1 wire810 (.A(_12245_),
    .X(net810));
 sky130_fd_sc_hd__buf_1 wire811 (.A(_12196_),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_1 wire812 (.A(net813),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_1 wire813 (.A(_11238_),
    .X(net813));
 sky130_fd_sc_hd__buf_1 wire814 (.A(_10415_),
    .X(net814));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire815 (.A(net816),
    .X(net815));
 sky130_fd_sc_hd__clkbuf_1 wire816 (.A(_10146_),
    .X(net816));
 sky130_fd_sc_hd__clkbuf_1 wire817 (.A(_10019_),
    .X(net817));
 sky130_fd_sc_hd__clkbuf_1 wire818 (.A(_09996_),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_1 wire819 (.A(_09972_),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_1 wire820 (.A(net821),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_1 wire821 (.A(_09470_),
    .X(net821));
 sky130_fd_sc_hd__buf_1 wire822 (.A(_09100_),
    .X(net822));
 sky130_fd_sc_hd__buf_1 wire823 (.A(net824),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_1 wire824 (.A(net825),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_1 wire825 (.A(_08702_),
    .X(net825));
 sky130_fd_sc_hd__buf_1 wire826 (.A(_07961_),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_2 wire827 (.A(net828),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_1 wire828 (.A(_07860_),
    .X(net828));
 sky130_fd_sc_hd__buf_1 wire829 (.A(_07330_),
    .X(net829));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire830 (.A(_07166_),
    .X(net830));
 sky130_fd_sc_hd__clkbuf_2 max_length831 (.A(net832),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_2 max_length832 (.A(_06652_),
    .X(net832));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire833 (.A(_06410_),
    .X(net833));
 sky130_fd_sc_hd__buf_1 wire834 (.A(_06373_),
    .X(net834));
 sky130_fd_sc_hd__buf_1 wire835 (.A(_06240_),
    .X(net835));
 sky130_fd_sc_hd__buf_1 wire836 (.A(_06184_),
    .X(net836));
 sky130_fd_sc_hd__buf_1 wire837 (.A(net838),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_1 wire838 (.A(_06114_),
    .X(net838));
 sky130_fd_sc_hd__buf_1 wire839 (.A(_06109_),
    .X(net839));
 sky130_fd_sc_hd__buf_1 wire840 (.A(_06062_),
    .X(net840));
 sky130_fd_sc_hd__buf_1 wire841 (.A(_06045_),
    .X(net841));
 sky130_fd_sc_hd__buf_1 wire842 (.A(_05631_),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_2 wire843 (.A(_05626_),
    .X(net843));
 sky130_fd_sc_hd__buf_1 wire844 (.A(_05603_),
    .X(net844));
 sky130_fd_sc_hd__buf_1 wire845 (.A(_05576_),
    .X(net845));
 sky130_fd_sc_hd__buf_1 wire846 (.A(_05549_),
    .X(net846));
 sky130_fd_sc_hd__buf_1 wire847 (.A(_05503_),
    .X(net847));
 sky130_fd_sc_hd__buf_1 wire848 (.A(_05402_),
    .X(net848));
 sky130_fd_sc_hd__buf_1 wire849 (.A(_05395_),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_2 wire850 (.A(_05183_),
    .X(net850));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire851 (.A(_05019_),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_1 wire852 (.A(net853),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_1 wire853 (.A(_04100_),
    .X(net853));
 sky130_fd_sc_hd__buf_1 wire854 (.A(_03858_),
    .X(net854));
 sky130_fd_sc_hd__buf_1 wire855 (.A(_03639_),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_1 wire856 (.A(net857),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_1 max_length857 (.A(net858),
    .X(net857));
 sky130_fd_sc_hd__buf_1 wire858 (.A(_02592_),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_2 wire859 (.A(_02158_),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_2 wire860 (.A(_01416_),
    .X(net860));
 sky130_fd_sc_hd__buf_1 wire861 (.A(_01230_),
    .X(net861));
 sky130_fd_sc_hd__buf_1 wire862 (.A(_01015_),
    .X(net862));
 sky130_fd_sc_hd__buf_1 wire863 (.A(net864),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_1 wire864 (.A(_12218_),
    .X(net864));
 sky130_fd_sc_hd__buf_1 wire865 (.A(_12173_),
    .X(net865));
 sky130_fd_sc_hd__buf_1 wire866 (.A(_12026_),
    .X(net866));
 sky130_fd_sc_hd__buf_1 wire867 (.A(_12012_),
    .X(net867));
 sky130_fd_sc_hd__buf_1 wire868 (.A(_11978_),
    .X(net868));
 sky130_fd_sc_hd__clkbuf_1 wire869 (.A(net870),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_1 wire870 (.A(net871),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_1 wire871 (.A(_11240_),
    .X(net871));
 sky130_fd_sc_hd__buf_1 wire872 (.A(_11022_),
    .X(net872));
 sky130_fd_sc_hd__buf_1 wire873 (.A(_10725_),
    .X(net873));
 sky130_fd_sc_hd__buf_1 wire874 (.A(net875),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_1 wire875 (.A(_10269_),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_1 wire876 (.A(_09519_),
    .X(net876));
 sky130_fd_sc_hd__clkbuf_1 wire877 (.A(_09467_),
    .X(net877));
 sky130_fd_sc_hd__buf_1 wire878 (.A(_08940_),
    .X(net878));
 sky130_fd_sc_hd__buf_1 wire879 (.A(_08568_),
    .X(net879));
 sky130_fd_sc_hd__buf_1 wire880 (.A(_08567_),
    .X(net880));
 sky130_fd_sc_hd__buf_1 wire881 (.A(_08446_),
    .X(net881));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire882 (.A(_08386_),
    .X(net882));
 sky130_fd_sc_hd__clkbuf_1 wire883 (.A(_08060_),
    .X(net883));
 sky130_fd_sc_hd__buf_1 wire884 (.A(net885),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_1 wire885 (.A(net886),
    .X(net885));
 sky130_fd_sc_hd__clkbuf_1 wire886 (.A(_07962_),
    .X(net886));
 sky130_fd_sc_hd__buf_1 wire887 (.A(_07777_),
    .X(net887));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire888 (.A(_07669_),
    .X(net888));
 sky130_fd_sc_hd__buf_1 wire889 (.A(_07592_),
    .X(net889));
 sky130_fd_sc_hd__clkbuf_1 wire890 (.A(net891),
    .X(net890));
 sky130_fd_sc_hd__clkbuf_1 wire891 (.A(_06864_),
    .X(net891));
 sky130_fd_sc_hd__buf_1 wire892 (.A(net893),
    .X(net892));
 sky130_fd_sc_hd__buf_1 wire893 (.A(net894),
    .X(net893));
 sky130_fd_sc_hd__buf_1 wire894 (.A(_06651_),
    .X(net894));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire895 (.A(net896),
    .X(net895));
 sky130_fd_sc_hd__clkbuf_2 wire896 (.A(_06606_),
    .X(net896));
 sky130_fd_sc_hd__buf_1 wire897 (.A(net898),
    .X(net897));
 sky130_fd_sc_hd__buf_1 max_length898 (.A(_06606_),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_2 wire899 (.A(_06572_),
    .X(net899));
 sky130_fd_sc_hd__buf_1 wire900 (.A(net901),
    .X(net900));
 sky130_fd_sc_hd__buf_1 wire901 (.A(_06572_),
    .X(net901));
 sky130_fd_sc_hd__clkbuf_2 wire902 (.A(net903),
    .X(net902));
 sky130_fd_sc_hd__buf_1 wire903 (.A(net904),
    .X(net903));
 sky130_fd_sc_hd__buf_1 wire904 (.A(net905),
    .X(net904));
 sky130_fd_sc_hd__buf_1 max_length905 (.A(_06543_),
    .X(net905));
 sky130_fd_sc_hd__buf_1 wire906 (.A(_06199_),
    .X(net906));
 sky130_fd_sc_hd__buf_1 wire907 (.A(net908),
    .X(net907));
 sky130_fd_sc_hd__clkbuf_1 wire908 (.A(_06123_),
    .X(net908));
 sky130_fd_sc_hd__buf_1 wire909 (.A(net910),
    .X(net909));
 sky130_fd_sc_hd__clkbuf_1 wire910 (.A(_05964_),
    .X(net910));
 sky130_fd_sc_hd__clkbuf_1 wire911 (.A(_05890_),
    .X(net911));
 sky130_fd_sc_hd__buf_1 wire912 (.A(_05737_),
    .X(net912));
 sky130_fd_sc_hd__buf_1 wire913 (.A(net914),
    .X(net913));
 sky130_fd_sc_hd__clkbuf_1 wire914 (.A(_05723_),
    .X(net914));
 sky130_fd_sc_hd__buf_1 wire915 (.A(_05718_),
    .X(net915));
 sky130_fd_sc_hd__buf_1 wire916 (.A(_05714_),
    .X(net916));
 sky130_fd_sc_hd__clkbuf_1 wire917 (.A(_05411_),
    .X(net917));
 sky130_fd_sc_hd__buf_1 wire918 (.A(_05409_),
    .X(net918));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire919 (.A(_05356_),
    .X(net919));
 sky130_fd_sc_hd__buf_1 wire920 (.A(net921),
    .X(net920));
 sky130_fd_sc_hd__clkbuf_1 wire921 (.A(_05299_),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_1 wire922 (.A(net923),
    .X(net922));
 sky130_fd_sc_hd__clkbuf_1 wire923 (.A(_04649_),
    .X(net923));
 sky130_fd_sc_hd__clkbuf_1 wire924 (.A(net925),
    .X(net924));
 sky130_fd_sc_hd__clkbuf_1 wire925 (.A(_04648_),
    .X(net925));
 sky130_fd_sc_hd__clkbuf_1 wire926 (.A(_04646_),
    .X(net926));
 sky130_fd_sc_hd__clkbuf_1 wire927 (.A(_04645_),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_1 wire928 (.A(_04311_),
    .X(net928));
 sky130_fd_sc_hd__buf_1 wire929 (.A(_04242_),
    .X(net929));
 sky130_fd_sc_hd__buf_1 wire930 (.A(net931),
    .X(net930));
 sky130_fd_sc_hd__clkbuf_1 wire931 (.A(_04020_),
    .X(net931));
 sky130_fd_sc_hd__buf_1 wire932 (.A(_03828_),
    .X(net932));
 sky130_fd_sc_hd__buf_1 wire933 (.A(_03543_),
    .X(net933));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire934 (.A(net935),
    .X(net934));
 sky130_fd_sc_hd__clkbuf_1 wire935 (.A(net936),
    .X(net935));
 sky130_fd_sc_hd__clkbuf_1 wire936 (.A(net937),
    .X(net936));
 sky130_fd_sc_hd__clkbuf_1 wire937 (.A(_03319_),
    .X(net937));
 sky130_fd_sc_hd__buf_1 wire938 (.A(_03303_),
    .X(net938));
 sky130_fd_sc_hd__clkbuf_1 wire939 (.A(net940),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_1 wire940 (.A(_02587_),
    .X(net940));
 sky130_fd_sc_hd__buf_1 wire941 (.A(net942),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_1 wire942 (.A(_02581_),
    .X(net942));
 sky130_fd_sc_hd__buf_1 wire943 (.A(_02239_),
    .X(net943));
 sky130_fd_sc_hd__clkbuf_4 wire944 (.A(_02201_),
    .X(net944));
 sky130_fd_sc_hd__buf_1 wire945 (.A(_02078_),
    .X(net945));
 sky130_fd_sc_hd__buf_1 wire946 (.A(_01734_),
    .X(net946));
 sky130_fd_sc_hd__buf_1 wire947 (.A(_01517_),
    .X(net947));
 sky130_fd_sc_hd__clkbuf_2 wire948 (.A(_01503_),
    .X(net948));
 sky130_fd_sc_hd__buf_1 wire949 (.A(net950),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_2 wire950 (.A(_12135_),
    .X(net950));
 sky130_fd_sc_hd__buf_1 wire951 (.A(_12122_),
    .X(net951));
 sky130_fd_sc_hd__buf_1 wire952 (.A(_11977_),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_2 wire953 (.A(net954),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_1 wire954 (.A(net955),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_1 wire955 (.A(_11623_),
    .X(net955));
 sky130_fd_sc_hd__buf_1 wire956 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_1 wire957 (.A(_11598_),
    .X(net957));
 sky130_fd_sc_hd__buf_1 wire958 (.A(net959),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_1 wire959 (.A(_11597_),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_1 wire960 (.A(_11304_),
    .X(net960));
 sky130_fd_sc_hd__buf_1 wire961 (.A(_10382_),
    .X(net961));
 sky130_fd_sc_hd__buf_1 wire962 (.A(_09949_),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_2 wire963 (.A(_09824_),
    .X(net963));
 sky130_fd_sc_hd__clkbuf_1 wire964 (.A(_09570_),
    .X(net964));
 sky130_fd_sc_hd__clkbuf_1 wire965 (.A(_09464_),
    .X(net965));
 sky130_fd_sc_hd__buf_1 wire966 (.A(_08993_),
    .X(net966));
 sky130_fd_sc_hd__buf_1 wire967 (.A(net968),
    .X(net967));
 sky130_fd_sc_hd__clkbuf_1 wire968 (.A(net969),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_1 wire969 (.A(net970),
    .X(net969));
 sky130_fd_sc_hd__buf_1 wire970 (.A(net971),
    .X(net970));
 sky130_fd_sc_hd__clkbuf_1 wire971 (.A(_08993_),
    .X(net971));
 sky130_fd_sc_hd__buf_1 wire972 (.A(net973),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_1 wire973 (.A(net974),
    .X(net973));
 sky130_fd_sc_hd__clkbuf_1 wire974 (.A(_08696_),
    .X(net974));
 sky130_fd_sc_hd__buf_1 wire975 (.A(_08520_),
    .X(net975));
 sky130_fd_sc_hd__buf_2 wire976 (.A(net977),
    .X(net976));
 sky130_fd_sc_hd__clkbuf_1 wire977 (.A(_08444_),
    .X(net977));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire978 (.A(_08335_),
    .X(net978));
 sky130_fd_sc_hd__buf_1 wire979 (.A(net980),
    .X(net979));
 sky130_fd_sc_hd__clkbuf_1 wire980 (.A(_08269_),
    .X(net980));
 sky130_fd_sc_hd__buf_1 wire981 (.A(net982),
    .X(net981));
 sky130_fd_sc_hd__clkbuf_1 wire982 (.A(_08266_),
    .X(net982));
 sky130_fd_sc_hd__buf_1 wire983 (.A(_08204_),
    .X(net983));
 sky130_fd_sc_hd__buf_1 wire984 (.A(net985),
    .X(net984));
 sky130_fd_sc_hd__clkbuf_1 wire985 (.A(net986),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_1 wire986 (.A(_07934_),
    .X(net986));
 sky130_fd_sc_hd__buf_1 wire987 (.A(_07833_),
    .X(net987));
 sky130_fd_sc_hd__buf_1 wire988 (.A(net989),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_1 wire989 (.A(_07727_),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_2 wire990 (.A(_07301_),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_2 wire991 (.A(_07168_),
    .X(net991));
 sky130_fd_sc_hd__buf_1 wire992 (.A(net993),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_1 wire993 (.A(_06910_),
    .X(net993));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire994 (.A(net995),
    .X(net994));
 sky130_fd_sc_hd__buf_1 max_length995 (.A(_06542_),
    .X(net995));
 sky130_fd_sc_hd__buf_1 wire996 (.A(_06070_),
    .X(net996));
 sky130_fd_sc_hd__buf_1 wire997 (.A(_05739_),
    .X(net997));
 sky130_fd_sc_hd__buf_1 wire998 (.A(_05735_),
    .X(net998));
 sky130_fd_sc_hd__buf_1 wire999 (.A(_05447_),
    .X(net999));
 sky130_fd_sc_hd__buf_1 wire1000 (.A(_05446_),
    .X(net1000));
 sky130_fd_sc_hd__buf_1 wire1001 (.A(_05359_),
    .X(net1001));
 sky130_fd_sc_hd__clkbuf_1 wire1002 (.A(_05230_),
    .X(net1002));
 sky130_fd_sc_hd__buf_1 wire1003 (.A(_05220_),
    .X(net1003));
 sky130_fd_sc_hd__clkbuf_2 wire1004 (.A(_05198_),
    .X(net1004));
 sky130_fd_sc_hd__buf_1 wire1005 (.A(_05117_),
    .X(net1005));
 sky130_fd_sc_hd__buf_1 wire1006 (.A(_05116_),
    .X(net1006));
 sky130_fd_sc_hd__buf_1 wire1007 (.A(_05049_),
    .X(net1007));
 sky130_fd_sc_hd__buf_2 wire1008 (.A(_04948_),
    .X(net1008));
 sky130_fd_sc_hd__buf_1 wire1009 (.A(_04569_),
    .X(net1009));
 sky130_fd_sc_hd__buf_1 wire1010 (.A(_04549_),
    .X(net1010));
 sky130_fd_sc_hd__buf_1 wire1011 (.A(_04539_),
    .X(net1011));
 sky130_fd_sc_hd__buf_1 wire1012 (.A(_04236_),
    .X(net1012));
 sky130_fd_sc_hd__clkbuf_2 wire1013 (.A(net1014),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_1 wire1014 (.A(_04089_),
    .X(net1014));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1015 (.A(_04006_),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_1 wire1016 (.A(net1017),
    .X(net1016));
 sky130_fd_sc_hd__buf_1 wire1017 (.A(_03768_),
    .X(net1017));
 sky130_fd_sc_hd__buf_1 wire1018 (.A(_03540_),
    .X(net1018));
 sky130_fd_sc_hd__buf_1 wire1019 (.A(_03511_),
    .X(net1019));
 sky130_fd_sc_hd__buf_1 wire1020 (.A(net1021),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_1 wire1021 (.A(net1022),
    .X(net1021));
 sky130_fd_sc_hd__clkbuf_1 wire1022 (.A(net1023),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_1 wire1023 (.A(_03466_),
    .X(net1023));
 sky130_fd_sc_hd__buf_1 wire1024 (.A(net1025),
    .X(net1024));
 sky130_fd_sc_hd__clkbuf_1 wire1025 (.A(net1026),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_1 wire1026 (.A(net1027),
    .X(net1026));
 sky130_fd_sc_hd__clkbuf_1 wire1027 (.A(_03375_),
    .X(net1027));
 sky130_fd_sc_hd__buf_1 wire1028 (.A(net1029),
    .X(net1028));
 sky130_fd_sc_hd__clkbuf_1 wire1029 (.A(net1030),
    .X(net1029));
 sky130_fd_sc_hd__clkbuf_1 wire1030 (.A(_03321_),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_2 wire1031 (.A(_02986_),
    .X(net1031));
 sky130_fd_sc_hd__buf_1 wire1032 (.A(_02921_),
    .X(net1032));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1033 (.A(net1034),
    .X(net1033));
 sky130_fd_sc_hd__clkbuf_1 wire1034 (.A(net1035),
    .X(net1034));
 sky130_fd_sc_hd__clkbuf_1 wire1035 (.A(_02235_),
    .X(net1035));
 sky130_fd_sc_hd__buf_1 wire1036 (.A(net1037),
    .X(net1036));
 sky130_fd_sc_hd__clkbuf_1 wire1037 (.A(_02149_),
    .X(net1037));
 sky130_fd_sc_hd__buf_1 wire1038 (.A(net1039),
    .X(net1038));
 sky130_fd_sc_hd__clkbuf_1 wire1039 (.A(net1040),
    .X(net1039));
 sky130_fd_sc_hd__clkbuf_1 wire1040 (.A(_02053_),
    .X(net1040));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1041 (.A(net1042),
    .X(net1041));
 sky130_fd_sc_hd__clkbuf_1 wire1042 (.A(net1043),
    .X(net1042));
 sky130_fd_sc_hd__clkbuf_1 wire1043 (.A(_02051_),
    .X(net1043));
 sky130_fd_sc_hd__buf_1 wire1044 (.A(_01983_),
    .X(net1044));
 sky130_fd_sc_hd__buf_2 wire1045 (.A(_01954_),
    .X(net1045));
 sky130_fd_sc_hd__buf_1 wire1046 (.A(_01890_),
    .X(net1046));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1047 (.A(_01829_),
    .X(net1047));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1048 (.A(_01746_),
    .X(net1048));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1049 (.A(_01480_),
    .X(net1049));
 sky130_fd_sc_hd__buf_1 wire1050 (.A(_01302_),
    .X(net1050));
 sky130_fd_sc_hd__buf_1 wire1051 (.A(_01013_),
    .X(net1051));
 sky130_fd_sc_hd__buf_1 wire1052 (.A(_00818_),
    .X(net1052));
 sky130_fd_sc_hd__buf_1 wire1053 (.A(_12292_),
    .X(net1053));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1054 (.A(_12145_),
    .X(net1054));
 sky130_fd_sc_hd__buf_1 wire1055 (.A(_11951_),
    .X(net1055));
 sky130_fd_sc_hd__clkbuf_2 wire1056 (.A(_11570_),
    .X(net1056));
 sky130_fd_sc_hd__buf_1 wire1057 (.A(_11540_),
    .X(net1057));
 sky130_fd_sc_hd__buf_1 wire1058 (.A(net1059),
    .X(net1058));
 sky130_fd_sc_hd__clkbuf_1 wire1059 (.A(_11526_),
    .X(net1059));
 sky130_fd_sc_hd__clkbuf_2 wire1060 (.A(_11316_),
    .X(net1060));
 sky130_fd_sc_hd__buf_1 wire1061 (.A(net1062),
    .X(net1061));
 sky130_fd_sc_hd__clkbuf_1 wire1062 (.A(net1063),
    .X(net1062));
 sky130_fd_sc_hd__clkbuf_1 wire1063 (.A(_11205_),
    .X(net1063));
 sky130_fd_sc_hd__buf_1 wire1064 (.A(_11011_),
    .X(net1064));
 sky130_fd_sc_hd__clkbuf_2 wire1065 (.A(_10578_),
    .X(net1065));
 sky130_fd_sc_hd__buf_1 wire1066 (.A(net1067),
    .X(net1066));
 sky130_fd_sc_hd__clkbuf_1 wire1067 (.A(net1068),
    .X(net1067));
 sky130_fd_sc_hd__clkbuf_1 wire1068 (.A(_10529_),
    .X(net1068));
 sky130_fd_sc_hd__buf_1 wire1069 (.A(_10450_),
    .X(net1069));
 sky130_fd_sc_hd__buf_1 wire1070 (.A(_10420_),
    .X(net1070));
 sky130_fd_sc_hd__clkbuf_2 wire1071 (.A(net1072),
    .X(net1071));
 sky130_fd_sc_hd__clkbuf_1 wire1072 (.A(_10356_),
    .X(net1072));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1073 (.A(_10184_),
    .X(net1073));
 sky130_fd_sc_hd__buf_1 wire1074 (.A(net1075),
    .X(net1074));
 sky130_fd_sc_hd__clkbuf_1 wire1075 (.A(_10086_),
    .X(net1075));
 sky130_fd_sc_hd__buf_1 wire1076 (.A(net1077),
    .X(net1076));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1077 (.A(_08992_),
    .X(net1077));
 sky130_fd_sc_hd__clkbuf_2 wire1078 (.A(net1079),
    .X(net1078));
 sky130_fd_sc_hd__clkbuf_2 wire1079 (.A(net1080),
    .X(net1079));
 sky130_fd_sc_hd__clkbuf_1 wire1080 (.A(_08410_),
    .X(net1080));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1081 (.A(net1082),
    .X(net1081));
 sky130_fd_sc_hd__clkbuf_1 wire1082 (.A(_08345_),
    .X(net1082));
 sky130_fd_sc_hd__buf_1 wire1083 (.A(_08316_),
    .X(net1083));
 sky130_fd_sc_hd__buf_1 wire1084 (.A(net1085),
    .X(net1084));
 sky130_fd_sc_hd__buf_1 wire1085 (.A(_08292_),
    .X(net1085));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1086 (.A(net1087),
    .X(net1086));
 sky130_fd_sc_hd__clkbuf_2 wire1087 (.A(_08290_),
    .X(net1087));
 sky130_fd_sc_hd__buf_1 wire1088 (.A(_08219_),
    .X(net1088));
 sky130_fd_sc_hd__buf_1 wire1089 (.A(net1090),
    .X(net1089));
 sky130_fd_sc_hd__clkbuf_1 wire1090 (.A(_08202_),
    .X(net1090));
 sky130_fd_sc_hd__buf_1 wire1091 (.A(_08182_),
    .X(net1091));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1092 (.A(_08129_),
    .X(net1092));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1093 (.A(_08113_),
    .X(net1093));
 sky130_fd_sc_hd__buf_1 wire1094 (.A(net1095),
    .X(net1094));
 sky130_fd_sc_hd__clkbuf_1 wire1095 (.A(net1096),
    .X(net1095));
 sky130_fd_sc_hd__clkbuf_1 wire1096 (.A(_07981_),
    .X(net1096));
 sky130_fd_sc_hd__buf_1 wire1097 (.A(net1098),
    .X(net1097));
 sky130_fd_sc_hd__clkbuf_1 wire1098 (.A(_07758_),
    .X(net1098));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1099 (.A(net1100),
    .X(net1099));
 sky130_fd_sc_hd__clkbuf_1 wire1100 (.A(net1101),
    .X(net1100));
 sky130_fd_sc_hd__clkbuf_1 wire1101 (.A(net1102),
    .X(net1101));
 sky130_fd_sc_hd__clkbuf_1 wire1102 (.A(net1103),
    .X(net1102));
 sky130_fd_sc_hd__clkbuf_1 wire1103 (.A(_07744_),
    .X(net1103));
 sky130_fd_sc_hd__buf_1 wire1104 (.A(net1105),
    .X(net1104));
 sky130_fd_sc_hd__clkbuf_1 wire1105 (.A(net1106),
    .X(net1105));
 sky130_fd_sc_hd__clkbuf_1 wire1106 (.A(net1107),
    .X(net1106));
 sky130_fd_sc_hd__clkbuf_1 wire1107 (.A(_07703_),
    .X(net1107));
 sky130_fd_sc_hd__buf_1 wire1108 (.A(_07660_),
    .X(net1108));
 sky130_fd_sc_hd__clkbuf_2 wire1109 (.A(net1110),
    .X(net1109));
 sky130_fd_sc_hd__clkbuf_1 wire1110 (.A(net1111),
    .X(net1110));
 sky130_fd_sc_hd__clkbuf_1 wire1111 (.A(net1112),
    .X(net1111));
 sky130_fd_sc_hd__clkbuf_1 wire1112 (.A(_07612_),
    .X(net1112));
 sky130_fd_sc_hd__clkbuf_2 wire1113 (.A(net1114),
    .X(net1113));
 sky130_fd_sc_hd__clkbuf_1 wire1114 (.A(net1115),
    .X(net1114));
 sky130_fd_sc_hd__clkbuf_1 wire1115 (.A(_07523_),
    .X(net1115));
 sky130_fd_sc_hd__buf_1 wire1116 (.A(_07428_),
    .X(net1116));
 sky130_fd_sc_hd__buf_1 wire1117 (.A(_07163_),
    .X(net1117));
 sky130_fd_sc_hd__clkbuf_1 wire1118 (.A(_06857_),
    .X(net1118));
 sky130_fd_sc_hd__clkbuf_2 max_length1119 (.A(net1120),
    .X(net1119));
 sky130_fd_sc_hd__buf_1 wire1120 (.A(_06405_),
    .X(net1120));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1121 (.A(net1123),
    .X(net1121));
 sky130_fd_sc_hd__buf_1 wire1122 (.A(net1123),
    .X(net1122));
 sky130_fd_sc_hd__clkbuf_2 wire1123 (.A(_06326_),
    .X(net1123));
 sky130_fd_sc_hd__buf_1 wire1124 (.A(net1125),
    .X(net1124));
 sky130_fd_sc_hd__clkbuf_2 wire1125 (.A(_06218_),
    .X(net1125));
 sky130_fd_sc_hd__clkbuf_2 wire1126 (.A(net1127),
    .X(net1126));
 sky130_fd_sc_hd__clkbuf_2 wire1127 (.A(_05780_),
    .X(net1127));
 sky130_fd_sc_hd__buf_1 wire1128 (.A(_05712_),
    .X(net1128));
 sky130_fd_sc_hd__buf_1 wire1129 (.A(_05706_),
    .X(net1129));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1130 (.A(_05640_),
    .X(net1130));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1131 (.A(_05583_),
    .X(net1131));
 sky130_fd_sc_hd__buf_1 wire1132 (.A(_05557_),
    .X(net1132));
 sky130_fd_sc_hd__buf_1 wire1133 (.A(net1134),
    .X(net1133));
 sky130_fd_sc_hd__clkbuf_1 wire1134 (.A(_05513_),
    .X(net1134));
 sky130_fd_sc_hd__buf_1 wire1135 (.A(_05494_),
    .X(net1135));
 sky130_fd_sc_hd__buf_1 wire1136 (.A(_05439_),
    .X(net1136));
 sky130_fd_sc_hd__buf_1 wire1137 (.A(_05438_),
    .X(net1137));
 sky130_fd_sc_hd__buf_1 wire1138 (.A(net1139),
    .X(net1138));
 sky130_fd_sc_hd__clkbuf_1 wire1139 (.A(_05377_),
    .X(net1139));
 sky130_fd_sc_hd__clkbuf_2 wire1140 (.A(net1141),
    .X(net1140));
 sky130_fd_sc_hd__clkbuf_1 wire1141 (.A(net1142),
    .X(net1141));
 sky130_fd_sc_hd__clkbuf_1 wire1142 (.A(_05193_),
    .X(net1142));
 sky130_fd_sc_hd__buf_1 wire1143 (.A(_05174_),
    .X(net1143));
 sky130_fd_sc_hd__clkbuf_1 wire1144 (.A(net1145),
    .X(net1144));
 sky130_fd_sc_hd__clkbuf_1 wire1145 (.A(net1146),
    .X(net1145));
 sky130_fd_sc_hd__clkbuf_1 wire1146 (.A(_05066_),
    .X(net1146));
 sky130_fd_sc_hd__buf_1 wire1147 (.A(_05045_),
    .X(net1147));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1148 (.A(net1149),
    .X(net1148));
 sky130_fd_sc_hd__buf_1 wire1149 (.A(net1151),
    .X(net1149));
 sky130_fd_sc_hd__buf_1 wire1150 (.A(net1151),
    .X(net1150));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1151 (.A(net1152),
    .X(net1151));
 sky130_fd_sc_hd__clkbuf_1 wire1152 (.A(net1153),
    .X(net1152));
 sky130_fd_sc_hd__clkbuf_1 wire1153 (.A(_05026_),
    .X(net1153));
 sky130_fd_sc_hd__clkbuf_1 max_length1154 (.A(_05026_),
    .X(net1154));
 sky130_fd_sc_hd__buf_1 wire1155 (.A(net1156),
    .X(net1155));
 sky130_fd_sc_hd__clkbuf_1 wire1156 (.A(_05023_),
    .X(net1156));
 sky130_fd_sc_hd__buf_1 wire1157 (.A(_04782_),
    .X(net1157));
 sky130_fd_sc_hd__clkbuf_1 wire1158 (.A(_04548_),
    .X(net1158));
 sky130_fd_sc_hd__buf_1 wire1159 (.A(_04077_),
    .X(net1159));
 sky130_fd_sc_hd__buf_1 wire1160 (.A(_03923_),
    .X(net1160));
 sky130_fd_sc_hd__clkbuf_2 wire1161 (.A(_03829_),
    .X(net1161));
 sky130_fd_sc_hd__buf_1 wire1162 (.A(_03708_),
    .X(net1162));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1163 (.A(_03643_),
    .X(net1163));
 sky130_fd_sc_hd__buf_1 wire1164 (.A(_03615_),
    .X(net1164));
 sky130_fd_sc_hd__buf_1 wire1165 (.A(_03545_),
    .X(net1165));
 sky130_fd_sc_hd__buf_1 wire1166 (.A(_03301_),
    .X(net1166));
 sky130_fd_sc_hd__buf_1 wire1167 (.A(_03295_),
    .X(net1167));
 sky130_fd_sc_hd__buf_1 wire1168 (.A(_02147_),
    .X(net1168));
 sky130_fd_sc_hd__buf_1 wire1169 (.A(_02061_),
    .X(net1169));
 sky130_fd_sc_hd__clkbuf_2 wire1170 (.A(_01971_),
    .X(net1170));
 sky130_fd_sc_hd__buf_1 wire1171 (.A(_01858_),
    .X(net1171));
 sky130_fd_sc_hd__buf_1 wire1172 (.A(_01777_),
    .X(net1172));
 sky130_fd_sc_hd__buf_1 wire1173 (.A(_01687_),
    .X(net1173));
 sky130_fd_sc_hd__buf_1 wire1174 (.A(_01656_),
    .X(net1174));
 sky130_fd_sc_hd__clkbuf_1 wire1175 (.A(net1176),
    .X(net1175));
 sky130_fd_sc_hd__clkbuf_1 max_length1176 (.A(_01642_),
    .X(net1176));
 sky130_fd_sc_hd__buf_1 wire1177 (.A(_01584_),
    .X(net1177));
 sky130_fd_sc_hd__buf_1 wire1178 (.A(_01583_),
    .X(net1178));
 sky130_fd_sc_hd__clkbuf_2 wire1179 (.A(_01505_),
    .X(net1179));
 sky130_fd_sc_hd__buf_1 wire1180 (.A(_01482_),
    .X(net1180));
 sky130_fd_sc_hd__buf_1 wire1181 (.A(_01394_),
    .X(net1181));
 sky130_fd_sc_hd__clkbuf_2 wire1182 (.A(_01372_),
    .X(net1182));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1183 (.A(net1184),
    .X(net1183));
 sky130_fd_sc_hd__clkbuf_1 wire1184 (.A(_01020_),
    .X(net1184));
 sky130_fd_sc_hd__buf_1 wire1185 (.A(_01018_),
    .X(net1185));
 sky130_fd_sc_hd__buf_1 wire1186 (.A(_00929_),
    .X(net1186));
 sky130_fd_sc_hd__buf_1 wire1187 (.A(_00913_),
    .X(net1187));
 sky130_fd_sc_hd__clkbuf_2 wire1188 (.A(net1189),
    .X(net1188));
 sky130_fd_sc_hd__clkbuf_1 wire1189 (.A(net1190),
    .X(net1189));
 sky130_fd_sc_hd__clkbuf_1 wire1190 (.A(_11638_),
    .X(net1190));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1191 (.A(_11475_),
    .X(net1191));
 sky130_fd_sc_hd__buf_1 wire1192 (.A(_11218_),
    .X(net1192));
 sky130_fd_sc_hd__buf_1 wire1193 (.A(_11081_),
    .X(net1193));
 sky130_fd_sc_hd__buf_1 wire1194 (.A(_10721_),
    .X(net1194));
 sky130_fd_sc_hd__buf_1 wire1195 (.A(_10497_),
    .X(net1195));
 sky130_fd_sc_hd__buf_1 wire1196 (.A(_10419_),
    .X(net1196));
 sky130_fd_sc_hd__buf_1 wire1197 (.A(net1198),
    .X(net1197));
 sky130_fd_sc_hd__clkbuf_1 wire1198 (.A(_10362_),
    .X(net1198));
 sky130_fd_sc_hd__clkbuf_1 max_length1199 (.A(net1200),
    .X(net1199));
 sky130_fd_sc_hd__buf_1 wire1200 (.A(net1201),
    .X(net1200));
 sky130_fd_sc_hd__clkbuf_1 wire1201 (.A(net1204),
    .X(net1201));
 sky130_fd_sc_hd__buf_1 wire1202 (.A(net1203),
    .X(net1202));
 sky130_fd_sc_hd__buf_1 wire1203 (.A(_10343_),
    .X(net1203));
 sky130_fd_sc_hd__clkbuf_1 max_length1204 (.A(_10343_),
    .X(net1204));
 sky130_fd_sc_hd__buf_1 wire1205 (.A(net1206),
    .X(net1205));
 sky130_fd_sc_hd__clkbuf_1 wire1206 (.A(_10325_),
    .X(net1206));
 sky130_fd_sc_hd__buf_1 wire1207 (.A(_10291_),
    .X(net1207));
 sky130_fd_sc_hd__buf_1 wire1208 (.A(net1209),
    .X(net1208));
 sky130_fd_sc_hd__clkbuf_1 wire1209 (.A(_10272_),
    .X(net1209));
 sky130_fd_sc_hd__buf_1 wire1210 (.A(_10247_),
    .X(net1210));
 sky130_fd_sc_hd__buf_1 wire1211 (.A(_10181_),
    .X(net1211));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1212 (.A(_10007_),
    .X(net1212));
 sky130_fd_sc_hd__buf_1 wire1213 (.A(_09823_),
    .X(net1213));
 sky130_fd_sc_hd__clkbuf_2 max_length1214 (.A(net1215),
    .X(net1214));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1215 (.A(_09700_),
    .X(net1215));
 sky130_fd_sc_hd__buf_1 wire1216 (.A(net1219),
    .X(net1216));
 sky130_fd_sc_hd__buf_1 max_length1217 (.A(net1218),
    .X(net1217));
 sky130_fd_sc_hd__buf_1 wire1218 (.A(net1219),
    .X(net1218));
 sky130_fd_sc_hd__buf_1 wire1219 (.A(_09580_),
    .X(net1219));
 sky130_fd_sc_hd__clkbuf_1 wire1220 (.A(_09250_),
    .X(net1220));
 sky130_fd_sc_hd__buf_1 wire1221 (.A(net1222),
    .X(net1221));
 sky130_fd_sc_hd__clkbuf_1 wire1222 (.A(net1223),
    .X(net1222));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1223 (.A(net1224),
    .X(net1223));
 sky130_fd_sc_hd__clkbuf_1 wire1224 (.A(net1227),
    .X(net1224));
 sky130_fd_sc_hd__clkbuf_1 wire1225 (.A(net1226),
    .X(net1225));
 sky130_fd_sc_hd__buf_1 wire1226 (.A(_08991_),
    .X(net1226));
 sky130_fd_sc_hd__clkbuf_1 max_length1227 (.A(_08991_),
    .X(net1227));
 sky130_fd_sc_hd__clkbuf_1 wire1228 (.A(net1229),
    .X(net1228));
 sky130_fd_sc_hd__buf_1 wire1229 (.A(net1230),
    .X(net1229));
 sky130_fd_sc_hd__clkbuf_1 wire1230 (.A(net1231),
    .X(net1230));
 sky130_fd_sc_hd__buf_1 wire1231 (.A(net1232),
    .X(net1231));
 sky130_fd_sc_hd__buf_1 wire1232 (.A(net1233),
    .X(net1232));
 sky130_fd_sc_hd__buf_1 wire1233 (.A(net1234),
    .X(net1233));
 sky130_fd_sc_hd__buf_1 wire1234 (.A(net1235),
    .X(net1234));
 sky130_fd_sc_hd__clkbuf_1 wire1235 (.A(net1236),
    .X(net1235));
 sky130_fd_sc_hd__clkbuf_1 wire1236 (.A(_08917_),
    .X(net1236));
 sky130_fd_sc_hd__buf_1 wire1237 (.A(net1238),
    .X(net1237));
 sky130_fd_sc_hd__clkbuf_1 wire1238 (.A(net1239),
    .X(net1238));
 sky130_fd_sc_hd__buf_1 wire1239 (.A(_08917_),
    .X(net1239));
 sky130_fd_sc_hd__buf_1 wire1240 (.A(net1241),
    .X(net1240));
 sky130_fd_sc_hd__clkbuf_1 wire1241 (.A(_08690_),
    .X(net1241));
 sky130_fd_sc_hd__buf_1 wire1242 (.A(_08615_),
    .X(net1242));
 sky130_fd_sc_hd__buf_1 wire1243 (.A(_08578_),
    .X(net1243));
 sky130_fd_sc_hd__clkbuf_2 wire1244 (.A(_08515_),
    .X(net1244));
 sky130_fd_sc_hd__clkbuf_1 wire1245 (.A(_08509_),
    .X(net1245));
 sky130_fd_sc_hd__buf_1 wire1246 (.A(_08463_),
    .X(net1246));
 sky130_fd_sc_hd__buf_1 wire1247 (.A(_08419_),
    .X(net1247));
 sky130_fd_sc_hd__buf_1 wire1248 (.A(_08391_),
    .X(net1248));
 sky130_fd_sc_hd__buf_1 wire1249 (.A(_08331_),
    .X(net1249));
 sky130_fd_sc_hd__buf_2 wire1250 (.A(_08262_),
    .X(net1250));
 sky130_fd_sc_hd__buf_1 wire1251 (.A(_08252_),
    .X(net1251));
 sky130_fd_sc_hd__buf_1 max_length1252 (.A(net1253),
    .X(net1252));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1253 (.A(_08184_),
    .X(net1253));
 sky130_fd_sc_hd__buf_1 wire1254 (.A(net1255),
    .X(net1254));
 sky130_fd_sc_hd__clkbuf_1 wire1255 (.A(_08183_),
    .X(net1255));
 sky130_fd_sc_hd__buf_1 wire1256 (.A(_08145_),
    .X(net1256));
 sky130_fd_sc_hd__buf_1 wire1257 (.A(_08071_),
    .X(net1257));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1258 (.A(net1259),
    .X(net1258));
 sky130_fd_sc_hd__clkbuf_1 wire1259 (.A(net1260),
    .X(net1259));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1260 (.A(_08058_),
    .X(net1260));
 sky130_fd_sc_hd__buf_1 wire1261 (.A(_08035_),
    .X(net1261));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1262 (.A(_07993_),
    .X(net1262));
 sky130_fd_sc_hd__buf_1 wire1263 (.A(_07903_),
    .X(net1263));
 sky130_fd_sc_hd__buf_1 wire1264 (.A(_07845_),
    .X(net1264));
 sky130_fd_sc_hd__buf_1 wire1265 (.A(_07807_),
    .X(net1265));
 sky130_fd_sc_hd__buf_1 wire1266 (.A(net1267),
    .X(net1266));
 sky130_fd_sc_hd__clkbuf_1 wire1267 (.A(_07706_),
    .X(net1267));
 sky130_fd_sc_hd__buf_1 wire1268 (.A(_07665_),
    .X(net1268));
 sky130_fd_sc_hd__buf_1 wire1269 (.A(_07662_),
    .X(net1269));
 sky130_fd_sc_hd__clkbuf_2 wire1270 (.A(net1271),
    .X(net1270));
 sky130_fd_sc_hd__clkbuf_1 wire1271 (.A(_07610_),
    .X(net1271));
 sky130_fd_sc_hd__buf_1 wire1272 (.A(_07587_),
    .X(net1272));
 sky130_fd_sc_hd__buf_1 wire1273 (.A(_07498_),
    .X(net1273));
 sky130_fd_sc_hd__clkbuf_2 wire1274 (.A(_07356_),
    .X(net1274));
 sky130_fd_sc_hd__clkbuf_2 wire1275 (.A(_07324_),
    .X(net1275));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1276 (.A(_07294_),
    .X(net1276));
 sky130_fd_sc_hd__buf_1 wire1277 (.A(_07201_),
    .X(net1277));
 sky130_fd_sc_hd__clkbuf_2 wire1278 (.A(net1279),
    .X(net1278));
 sky130_fd_sc_hd__clkbuf_1 wire1279 (.A(_07185_),
    .X(net1279));
 sky130_fd_sc_hd__clkbuf_2 wire1280 (.A(net1281),
    .X(net1280));
 sky130_fd_sc_hd__clkbuf_1 wire1281 (.A(net1282),
    .X(net1281));
 sky130_fd_sc_hd__clkbuf_1 wire1282 (.A(_07161_),
    .X(net1282));
 sky130_fd_sc_hd__buf_1 wire1283 (.A(net1284),
    .X(net1283));
 sky130_fd_sc_hd__clkbuf_1 wire1284 (.A(_07122_),
    .X(net1284));
 sky130_fd_sc_hd__buf_1 wire1285 (.A(_07105_),
    .X(net1285));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1286 (.A(_07070_),
    .X(net1286));
 sky130_fd_sc_hd__buf_1 wire1287 (.A(_07054_),
    .X(net1287));
 sky130_fd_sc_hd__clkbuf_1 wire1288 (.A(net1289),
    .X(net1288));
 sky130_fd_sc_hd__clkbuf_1 wire1289 (.A(_06854_),
    .X(net1289));
 sky130_fd_sc_hd__clkbuf_1 wire1290 (.A(net1291),
    .X(net1290));
 sky130_fd_sc_hd__clkbuf_1 wire1291 (.A(_06852_),
    .X(net1291));
 sky130_fd_sc_hd__clkbuf_2 wire1292 (.A(_06655_),
    .X(net1292));
 sky130_fd_sc_hd__buf_1 wire1293 (.A(net1294),
    .X(net1293));
 sky130_fd_sc_hd__buf_1 wire1294 (.A(_06608_),
    .X(net1294));
 sky130_fd_sc_hd__buf_1 wire1295 (.A(_06608_),
    .X(net1295));
 sky130_fd_sc_hd__buf_1 wire1296 (.A(net1297),
    .X(net1296));
 sky130_fd_sc_hd__clkbuf_2 max_length1297 (.A(net1298),
    .X(net1297));
 sky130_fd_sc_hd__buf_1 max_length1298 (.A(_06574_),
    .X(net1298));
 sky130_fd_sc_hd__clkbuf_2 wire1299 (.A(net1300),
    .X(net1299));
 sky130_fd_sc_hd__clkbuf_1 max_length1300 (.A(net1301),
    .X(net1300));
 sky130_fd_sc_hd__buf_1 max_length1301 (.A(net1302),
    .X(net1301));
 sky130_fd_sc_hd__buf_1 wire1302 (.A(_06522_),
    .X(net1302));
 sky130_fd_sc_hd__clkbuf_1 max_length1303 (.A(_06522_),
    .X(net1303));
 sky130_fd_sc_hd__clkbuf_2 wire1304 (.A(_06374_),
    .X(net1304));
 sky130_fd_sc_hd__buf_1 wire1305 (.A(_06245_),
    .X(net1305));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1306 (.A(net1307),
    .X(net1306));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1307 (.A(_05873_),
    .X(net1307));
 sky130_fd_sc_hd__buf_1 wire1308 (.A(net1309),
    .X(net1308));
 sky130_fd_sc_hd__clkbuf_1 wire1309 (.A(_05779_),
    .X(net1309));
 sky130_fd_sc_hd__buf_1 wire1310 (.A(_05753_),
    .X(net1310));
 sky130_fd_sc_hd__buf_1 wire1311 (.A(net1312),
    .X(net1311));
 sky130_fd_sc_hd__buf_1 wire1312 (.A(_05730_),
    .X(net1312));
 sky130_fd_sc_hd__buf_1 max_length1313 (.A(_05730_),
    .X(net1313));
 sky130_fd_sc_hd__buf_1 wire1314 (.A(net1315),
    .X(net1314));
 sky130_fd_sc_hd__buf_1 wire1315 (.A(net1316),
    .X(net1315));
 sky130_fd_sc_hd__buf_1 wire1316 (.A(_05687_),
    .X(net1316));
 sky130_fd_sc_hd__buf_1 wire1317 (.A(net1318),
    .X(net1317));
 sky130_fd_sc_hd__buf_1 wire1318 (.A(net1319),
    .X(net1318));
 sky130_fd_sc_hd__buf_1 wire1319 (.A(_05687_),
    .X(net1319));
 sky130_fd_sc_hd__buf_1 wire1320 (.A(_05611_),
    .X(net1320));
 sky130_fd_sc_hd__clkbuf_1 wire1321 (.A(net1322),
    .X(net1321));
 sky130_fd_sc_hd__buf_1 wire1322 (.A(net1323),
    .X(net1322));
 sky130_fd_sc_hd__buf_1 wire1323 (.A(net1324),
    .X(net1323));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1324 (.A(net1325),
    .X(net1324));
 sky130_fd_sc_hd__clkbuf_1 wire1325 (.A(net1326),
    .X(net1325));
 sky130_fd_sc_hd__buf_1 wire1326 (.A(net1327),
    .X(net1326));
 sky130_fd_sc_hd__buf_1 wire1327 (.A(net1328),
    .X(net1327));
 sky130_fd_sc_hd__buf_1 wire1328 (.A(net1329),
    .X(net1328));
 sky130_fd_sc_hd__clkbuf_1 wire1329 (.A(_05556_),
    .X(net1329));
 sky130_fd_sc_hd__buf_1 wire1330 (.A(_05526_),
    .X(net1330));
 sky130_fd_sc_hd__buf_1 wire1331 (.A(net1332),
    .X(net1331));
 sky130_fd_sc_hd__clkbuf_2 wire1332 (.A(_05294_),
    .X(net1332));
 sky130_fd_sc_hd__buf_1 wire1333 (.A(net1334),
    .X(net1333));
 sky130_fd_sc_hd__clkbuf_1 wire1334 (.A(net1335),
    .X(net1334));
 sky130_fd_sc_hd__clkbuf_1 wire1335 (.A(_05133_),
    .X(net1335));
 sky130_fd_sc_hd__clkbuf_2 wire1336 (.A(_05098_),
    .X(net1336));
 sky130_fd_sc_hd__clkbuf_1 max_length1337 (.A(net1338),
    .X(net1337));
 sky130_fd_sc_hd__clkbuf_2 wire1338 (.A(net1339),
    .X(net1338));
 sky130_fd_sc_hd__buf_1 wire1339 (.A(net1340),
    .X(net1339));
 sky130_fd_sc_hd__buf_1 wire1340 (.A(net1341),
    .X(net1340));
 sky130_fd_sc_hd__clkbuf_1 max_length1341 (.A(net1342),
    .X(net1341));
 sky130_fd_sc_hd__buf_1 wire1342 (.A(_05012_),
    .X(net1342));
 sky130_fd_sc_hd__clkbuf_2 wire1343 (.A(net1344),
    .X(net1343));
 sky130_fd_sc_hd__clkbuf_1 wire1344 (.A(net1345),
    .X(net1344));
 sky130_fd_sc_hd__clkbuf_1 wire1345 (.A(_04967_),
    .X(net1345));
 sky130_fd_sc_hd__buf_1 wire1346 (.A(_04921_),
    .X(net1346));
 sky130_fd_sc_hd__clkbuf_1 wire1347 (.A(net1348),
    .X(net1347));
 sky130_fd_sc_hd__clkbuf_1 wire1348 (.A(net1349),
    .X(net1348));
 sky130_fd_sc_hd__clkbuf_1 wire1349 (.A(net1351),
    .X(net1349));
 sky130_fd_sc_hd__clkbuf_2 max_length1350 (.A(net1351),
    .X(net1350));
 sky130_fd_sc_hd__buf_1 wire1351 (.A(_04921_),
    .X(net1351));
 sky130_fd_sc_hd__buf_1 wire1352 (.A(net1353),
    .X(net1352));
 sky130_fd_sc_hd__buf_1 wire1353 (.A(net1354),
    .X(net1353));
 sky130_fd_sc_hd__buf_1 wire1354 (.A(net1355),
    .X(net1354));
 sky130_fd_sc_hd__buf_1 max_length1355 (.A(net1356),
    .X(net1355));
 sky130_fd_sc_hd__buf_1 wire1356 (.A(_04902_),
    .X(net1356));
 sky130_fd_sc_hd__buf_1 wire1357 (.A(net1358),
    .X(net1357));
 sky130_fd_sc_hd__clkbuf_2 wire1358 (.A(net1359),
    .X(net1358));
 sky130_fd_sc_hd__buf_1 wire1359 (.A(_04735_),
    .X(net1359));
 sky130_fd_sc_hd__buf_1 wire1360 (.A(net1361),
    .X(net1360));
 sky130_fd_sc_hd__clkbuf_2 wire1361 (.A(net1362),
    .X(net1361));
 sky130_fd_sc_hd__buf_1 wire1362 (.A(_04702_),
    .X(net1362));
 sky130_fd_sc_hd__clkbuf_1 wire1363 (.A(net1364),
    .X(net1363));
 sky130_fd_sc_hd__clkbuf_1 wire1364 (.A(_04647_),
    .X(net1364));
 sky130_fd_sc_hd__buf_1 wire1365 (.A(net1366),
    .X(net1365));
 sky130_fd_sc_hd__buf_1 wire1366 (.A(_04543_),
    .X(net1366));
 sky130_fd_sc_hd__buf_1 wire1367 (.A(_04543_),
    .X(net1367));
 sky130_fd_sc_hd__buf_1 wire1368 (.A(net1369),
    .X(net1368));
 sky130_fd_sc_hd__buf_1 max_length1369 (.A(net1370),
    .X(net1369));
 sky130_fd_sc_hd__buf_1 wire1370 (.A(_04530_),
    .X(net1370));
 sky130_fd_sc_hd__buf_1 wire1371 (.A(_04530_),
    .X(net1371));
 sky130_fd_sc_hd__buf_1 wire1372 (.A(net1373),
    .X(net1372));
 sky130_fd_sc_hd__buf_1 wire1373 (.A(_04510_),
    .X(net1373));
 sky130_fd_sc_hd__buf_1 wire1374 (.A(_04510_),
    .X(net1374));
 sky130_fd_sc_hd__clkbuf_1 max_length1375 (.A(net1376),
    .X(net1375));
 sky130_fd_sc_hd__buf_1 wire1376 (.A(_04508_),
    .X(net1376));
 sky130_fd_sc_hd__buf_1 max_length1377 (.A(net1378),
    .X(net1377));
 sky130_fd_sc_hd__buf_1 wire1378 (.A(_04508_),
    .X(net1378));
 sky130_fd_sc_hd__buf_1 wire1379 (.A(_04072_),
    .X(net1379));
 sky130_fd_sc_hd__buf_1 wire1380 (.A(_04071_),
    .X(net1380));
 sky130_fd_sc_hd__clkbuf_1 wire1381 (.A(net1382),
    .X(net1381));
 sky130_fd_sc_hd__clkbuf_1 wire1382 (.A(net1383),
    .X(net1382));
 sky130_fd_sc_hd__buf_1 wire1383 (.A(_03668_),
    .X(net1383));
 sky130_fd_sc_hd__buf_1 wire1384 (.A(_03408_),
    .X(net1384));
 sky130_fd_sc_hd__buf_1 wire1385 (.A(net1386),
    .X(net1385));
 sky130_fd_sc_hd__clkbuf_1 wire1386 (.A(net1387),
    .X(net1386));
 sky130_fd_sc_hd__clkbuf_1 wire1387 (.A(_03280_),
    .X(net1387));
 sky130_fd_sc_hd__buf_1 wire1388 (.A(_02571_),
    .X(net1388));
 sky130_fd_sc_hd__buf_1 wire1389 (.A(_02121_),
    .X(net1389));
 sky130_fd_sc_hd__buf_1 wire1390 (.A(_01300_),
    .X(net1390));
 sky130_fd_sc_hd__buf_1 wire1391 (.A(_01277_),
    .X(net1391));
 sky130_fd_sc_hd__buf_1 wire1392 (.A(_00890_),
    .X(net1392));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1393 (.A(_00858_),
    .X(net1393));
 sky130_fd_sc_hd__buf_1 wire1394 (.A(_12428_),
    .X(net1394));
 sky130_fd_sc_hd__buf_1 wire1395 (.A(_12396_),
    .X(net1395));
 sky130_fd_sc_hd__clkbuf_2 wire1396 (.A(net1397),
    .X(net1396));
 sky130_fd_sc_hd__clkbuf_1 wire1397 (.A(_12378_),
    .X(net1397));
 sky130_fd_sc_hd__buf_1 wire1398 (.A(net1400),
    .X(net1398));
 sky130_fd_sc_hd__buf_1 wire1399 (.A(net1400),
    .X(net1399));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1400 (.A(net1401),
    .X(net1400));
 sky130_fd_sc_hd__clkbuf_1 wire1401 (.A(net1402),
    .X(net1401));
 sky130_fd_sc_hd__clkbuf_1 wire1402 (.A(net1403),
    .X(net1402));
 sky130_fd_sc_hd__buf_1 max_length1403 (.A(_12142_),
    .X(net1403));
 sky130_fd_sc_hd__clkbuf_2 wire1404 (.A(net1405),
    .X(net1404));
 sky130_fd_sc_hd__clkbuf_1 wire1405 (.A(_11857_),
    .X(net1405));
 sky130_fd_sc_hd__clkbuf_2 wire1406 (.A(net1407),
    .X(net1406));
 sky130_fd_sc_hd__clkbuf_1 wire1407 (.A(_11796_),
    .X(net1407));
 sky130_fd_sc_hd__buf_1 wire1408 (.A(_11770_),
    .X(net1408));
 sky130_fd_sc_hd__clkbuf_2 wire1409 (.A(_11760_),
    .X(net1409));
 sky130_fd_sc_hd__buf_1 wire1410 (.A(net1411),
    .X(net1410));
 sky130_fd_sc_hd__clkbuf_1 wire1411 (.A(_11753_),
    .X(net1411));
 sky130_fd_sc_hd__buf_1 wire1412 (.A(net1413),
    .X(net1412));
 sky130_fd_sc_hd__clkbuf_1 wire1413 (.A(net1414),
    .X(net1413));
 sky130_fd_sc_hd__clkbuf_1 wire1414 (.A(_11685_),
    .X(net1414));
 sky130_fd_sc_hd__buf_1 wire1415 (.A(_11510_),
    .X(net1415));
 sky130_fd_sc_hd__buf_1 wire1416 (.A(_11407_),
    .X(net1416));
 sky130_fd_sc_hd__buf_1 wire1417 (.A(_11399_),
    .X(net1417));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1418 (.A(_11390_),
    .X(net1418));
 sky130_fd_sc_hd__buf_1 wire1419 (.A(_11340_),
    .X(net1419));
 sky130_fd_sc_hd__clkbuf_1 wire1420 (.A(_11305_),
    .X(net1420));
 sky130_fd_sc_hd__buf_1 wire1421 (.A(_11173_),
    .X(net1421));
 sky130_fd_sc_hd__buf_1 wire1422 (.A(net1423),
    .X(net1422));
 sky130_fd_sc_hd__clkbuf_1 wire1423 (.A(net1424),
    .X(net1423));
 sky130_fd_sc_hd__clkbuf_1 wire1424 (.A(net1425),
    .X(net1424));
 sky130_fd_sc_hd__clkbuf_1 wire1425 (.A(_11067_),
    .X(net1425));
 sky130_fd_sc_hd__buf_1 wire1426 (.A(_11007_),
    .X(net1426));
 sky130_fd_sc_hd__clkbuf_1 wire1427 (.A(_10759_),
    .X(net1427));
 sky130_fd_sc_hd__buf_1 wire1428 (.A(_10674_),
    .X(net1428));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1429 (.A(_10586_),
    .X(net1429));
 sky130_fd_sc_hd__buf_1 wire1430 (.A(_10537_),
    .X(net1430));
 sky130_fd_sc_hd__buf_1 wire1431 (.A(net1432),
    .X(net1431));
 sky130_fd_sc_hd__clkbuf_1 wire1432 (.A(_10477_),
    .X(net1432));
 sky130_fd_sc_hd__buf_1 wire1433 (.A(net1434),
    .X(net1433));
 sky130_fd_sc_hd__clkbuf_1 wire1434 (.A(_10471_),
    .X(net1434));
 sky130_fd_sc_hd__clkbuf_1 wire1435 (.A(_10418_),
    .X(net1435));
 sky130_fd_sc_hd__buf_1 wire1436 (.A(_10392_),
    .X(net1436));
 sky130_fd_sc_hd__buf_1 wire1437 (.A(net1438),
    .X(net1437));
 sky130_fd_sc_hd__buf_1 wire1438 (.A(net1439),
    .X(net1438));
 sky130_fd_sc_hd__buf_1 wire1439 (.A(_10344_),
    .X(net1439));
 sky130_fd_sc_hd__buf_1 wire1440 (.A(_10306_),
    .X(net1440));
 sky130_fd_sc_hd__buf_1 wire1441 (.A(net1442),
    .X(net1441));
 sky130_fd_sc_hd__clkbuf_1 wire1442 (.A(_10274_),
    .X(net1442));
 sky130_fd_sc_hd__buf_1 wire1443 (.A(_10261_),
    .X(net1443));
 sky130_fd_sc_hd__buf_1 wire1444 (.A(net1445),
    .X(net1444));
 sky130_fd_sc_hd__buf_1 wire1445 (.A(net1446),
    .X(net1445));
 sky130_fd_sc_hd__buf_1 max_length1446 (.A(_10261_),
    .X(net1446));
 sky130_fd_sc_hd__clkbuf_2 wire1447 (.A(_09828_),
    .X(net1447));
 sky130_fd_sc_hd__buf_1 wire1448 (.A(_09628_),
    .X(net1448));
 sky130_fd_sc_hd__buf_1 wire1449 (.A(_09598_),
    .X(net1449));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1450 (.A(_09598_),
    .X(net1450));
 sky130_fd_sc_hd__buf_1 max_length1451 (.A(net1452),
    .X(net1451));
 sky130_fd_sc_hd__buf_1 wire1452 (.A(net1453),
    .X(net1452));
 sky130_fd_sc_hd__buf_1 wire1453 (.A(net1454),
    .X(net1453));
 sky130_fd_sc_hd__buf_1 wire1454 (.A(_09584_),
    .X(net1454));
 sky130_fd_sc_hd__buf_1 wire1455 (.A(_09579_),
    .X(net1455));
 sky130_fd_sc_hd__buf_1 wire1456 (.A(net1457),
    .X(net1456));
 sky130_fd_sc_hd__buf_1 wire1457 (.A(_09579_),
    .X(net1457));
 sky130_fd_sc_hd__clkbuf_1 wire1458 (.A(net1459),
    .X(net1458));
 sky130_fd_sc_hd__clkbuf_1 wire1459 (.A(_09509_),
    .X(net1459));
 sky130_fd_sc_hd__clkbuf_1 wire1460 (.A(_09455_),
    .X(net1460));
 sky130_fd_sc_hd__buf_1 wire1461 (.A(_09304_),
    .X(net1461));
 sky130_fd_sc_hd__clkbuf_1 wire1462 (.A(net1463),
    .X(net1462));
 sky130_fd_sc_hd__clkbuf_1 wire1463 (.A(net1464),
    .X(net1463));
 sky130_fd_sc_hd__clkbuf_1 wire1464 (.A(net1465),
    .X(net1464));
 sky130_fd_sc_hd__buf_1 max_length1465 (.A(_09204_),
    .X(net1465));
 sky130_fd_sc_hd__clkbuf_1 wire1466 (.A(net1467),
    .X(net1466));
 sky130_fd_sc_hd__clkbuf_1 wire1467 (.A(net1468),
    .X(net1467));
 sky130_fd_sc_hd__clkbuf_1 wire1468 (.A(net1469),
    .X(net1468));
 sky130_fd_sc_hd__clkbuf_1 max_length1469 (.A(_09068_),
    .X(net1469));
 sky130_fd_sc_hd__buf_1 max_length1470 (.A(net1471),
    .X(net1470));
 sky130_fd_sc_hd__buf_1 wire1471 (.A(net1472),
    .X(net1471));
 sky130_fd_sc_hd__clkbuf_1 wire1472 (.A(net1473),
    .X(net1472));
 sky130_fd_sc_hd__buf_1 wire1473 (.A(net1474),
    .X(net1473));
 sky130_fd_sc_hd__clkbuf_1 wire1474 (.A(net1475),
    .X(net1474));
 sky130_fd_sc_hd__buf_1 wire1475 (.A(_09068_),
    .X(net1475));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1476 (.A(net1477),
    .X(net1476));
 sky130_fd_sc_hd__clkbuf_1 wire1477 (.A(_09057_),
    .X(net1477));
 sky130_fd_sc_hd__buf_1 wire1478 (.A(_09036_),
    .X(net1478));
 sky130_fd_sc_hd__buf_1 max_length1479 (.A(net1480),
    .X(net1479));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1480 (.A(net1481),
    .X(net1480));
 sky130_fd_sc_hd__buf_1 wire1481 (.A(net1482),
    .X(net1481));
 sky130_fd_sc_hd__buf_1 wire1482 (.A(_08990_),
    .X(net1482));
 sky130_fd_sc_hd__buf_1 max_length1483 (.A(_08975_),
    .X(net1483));
 sky130_fd_sc_hd__clkbuf_2 wire1484 (.A(net1485),
    .X(net1484));
 sky130_fd_sc_hd__buf_1 wire1485 (.A(net1486),
    .X(net1485));
 sky130_fd_sc_hd__buf_1 wire1486 (.A(_08952_),
    .X(net1486));
 sky130_fd_sc_hd__clkbuf_1 wire1487 (.A(net1488),
    .X(net1487));
 sky130_fd_sc_hd__clkbuf_1 wire1488 (.A(net1489),
    .X(net1488));
 sky130_fd_sc_hd__clkbuf_1 wire1489 (.A(net1498),
    .X(net1489));
 sky130_fd_sc_hd__clkbuf_1 wire1490 (.A(net1491),
    .X(net1490));
 sky130_fd_sc_hd__buf_1 wire1491 (.A(net1493),
    .X(net1491));
 sky130_fd_sc_hd__clkbuf_1 wire1492 (.A(net1494),
    .X(net1492));
 sky130_fd_sc_hd__clkbuf_1 max_length1493 (.A(net1494),
    .X(net1493));
 sky130_fd_sc_hd__buf_1 wire1494 (.A(net1495),
    .X(net1494));
 sky130_fd_sc_hd__buf_1 wire1495 (.A(net1496),
    .X(net1495));
 sky130_fd_sc_hd__buf_1 wire1496 (.A(net1497),
    .X(net1496));
 sky130_fd_sc_hd__clkbuf_1 wire1497 (.A(_08916_),
    .X(net1497));
 sky130_fd_sc_hd__clkbuf_1 max_length1498 (.A(_08916_),
    .X(net1498));
 sky130_fd_sc_hd__clkbuf_1 wire1499 (.A(net1500),
    .X(net1499));
 sky130_fd_sc_hd__buf_1 wire1500 (.A(net1501),
    .X(net1500));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1501 (.A(_08905_),
    .X(net1501));
 sky130_fd_sc_hd__clkbuf_1 wire1502 (.A(net1503),
    .X(net1502));
 sky130_fd_sc_hd__clkbuf_1 wire1503 (.A(net1504),
    .X(net1503));
 sky130_fd_sc_hd__buf_1 wire1504 (.A(net1505),
    .X(net1504));
 sky130_fd_sc_hd__buf_1 wire1505 (.A(net1506),
    .X(net1505));
 sky130_fd_sc_hd__buf_1 wire1506 (.A(_08905_),
    .X(net1506));
 sky130_fd_sc_hd__buf_1 wire1507 (.A(_08417_),
    .X(net1507));
 sky130_fd_sc_hd__buf_1 wire1508 (.A(_08254_),
    .X(net1508));
 sky130_fd_sc_hd__buf_1 wire1509 (.A(net1510),
    .X(net1509));
 sky130_fd_sc_hd__clkbuf_1 max_length1510 (.A(_08251_),
    .X(net1510));
 sky130_fd_sc_hd__buf_1 wire1511 (.A(_08220_),
    .X(net1511));
 sky130_fd_sc_hd__buf_1 wire1512 (.A(_08175_),
    .X(net1512));
 sky130_fd_sc_hd__buf_1 wire1513 (.A(net1514),
    .X(net1513));
 sky130_fd_sc_hd__clkbuf_1 max_length1514 (.A(net1515),
    .X(net1514));
 sky130_fd_sc_hd__clkbuf_2 wire1515 (.A(_08106_),
    .X(net1515));
 sky130_fd_sc_hd__buf_1 wire1516 (.A(_08101_),
    .X(net1516));
 sky130_fd_sc_hd__buf_1 wire1517 (.A(_08070_),
    .X(net1517));
 sky130_fd_sc_hd__buf_1 wire1518 (.A(net1519),
    .X(net1518));
 sky130_fd_sc_hd__clkbuf_1 wire1519 (.A(_08045_),
    .X(net1519));
 sky130_fd_sc_hd__buf_1 wire1520 (.A(_08043_),
    .X(net1520));
 sky130_fd_sc_hd__buf_1 wire1521 (.A(_07992_),
    .X(net1521));
 sky130_fd_sc_hd__buf_1 wire1522 (.A(_07975_),
    .X(net1522));
 sky130_fd_sc_hd__buf_1 wire1523 (.A(net1524),
    .X(net1523));
 sky130_fd_sc_hd__clkbuf_1 wire1524 (.A(_07956_),
    .X(net1524));
 sky130_fd_sc_hd__buf_1 wire1525 (.A(net1526),
    .X(net1525));
 sky130_fd_sc_hd__buf_1 wire1526 (.A(_07950_),
    .X(net1526));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1527 (.A(net1528),
    .X(net1527));
 sky130_fd_sc_hd__clkbuf_1 max_length1528 (.A(_07902_),
    .X(net1528));
 sky130_fd_sc_hd__buf_1 wire1529 (.A(_07809_),
    .X(net1529));
 sky130_fd_sc_hd__clkbuf_2 wire1530 (.A(net1531),
    .X(net1530));
 sky130_fd_sc_hd__clkbuf_1 wire1531 (.A(net1532),
    .X(net1531));
 sky130_fd_sc_hd__clkbuf_1 wire1532 (.A(net1533),
    .X(net1532));
 sky130_fd_sc_hd__clkbuf_1 wire1533 (.A(net1534),
    .X(net1533));
 sky130_fd_sc_hd__clkbuf_1 wire1534 (.A(_07771_),
    .X(net1534));
 sky130_fd_sc_hd__buf_1 wire1535 (.A(_07766_),
    .X(net1535));
 sky130_fd_sc_hd__buf_1 wire1536 (.A(_07751_),
    .X(net1536));
 sky130_fd_sc_hd__buf_1 wire1537 (.A(_07678_),
    .X(net1537));
 sky130_fd_sc_hd__buf_1 wire1538 (.A(_07531_),
    .X(net1538));
 sky130_fd_sc_hd__clkbuf_2 wire1539 (.A(net1540),
    .X(net1539));
 sky130_fd_sc_hd__clkbuf_1 wire1540 (.A(net1541),
    .X(net1540));
 sky130_fd_sc_hd__clkbuf_1 wire1541 (.A(_07380_),
    .X(net1541));
 sky130_fd_sc_hd__buf_1 wire1542 (.A(_07359_),
    .X(net1542));
 sky130_fd_sc_hd__buf_1 wire1543 (.A(_07349_),
    .X(net1543));
 sky130_fd_sc_hd__buf_1 wire1544 (.A(_07277_),
    .X(net1544));
 sky130_fd_sc_hd__buf_1 wire1545 (.A(net1546),
    .X(net1545));
 sky130_fd_sc_hd__clkbuf_1 wire1546 (.A(_07244_),
    .X(net1546));
 sky130_fd_sc_hd__clkbuf_1 wire1547 (.A(_06849_),
    .X(net1547));
 sky130_fd_sc_hd__buf_1 wire1548 (.A(net1550),
    .X(net1548));
 sky130_fd_sc_hd__clkbuf_1 max_length1549 (.A(net1550),
    .X(net1549));
 sky130_fd_sc_hd__buf_1 wire1550 (.A(_06521_),
    .X(net1550));
 sky130_fd_sc_hd__buf_1 wire1551 (.A(net1552),
    .X(net1551));
 sky130_fd_sc_hd__buf_1 wire1552 (.A(net1553),
    .X(net1552));
 sky130_fd_sc_hd__buf_1 wire1553 (.A(_06509_),
    .X(net1553));
 sky130_fd_sc_hd__buf_1 wire1554 (.A(net1555),
    .X(net1554));
 sky130_fd_sc_hd__clkbuf_1 wire1555 (.A(net1556),
    .X(net1555));
 sky130_fd_sc_hd__buf_1 wire1556 (.A(net1557),
    .X(net1556));
 sky130_fd_sc_hd__clkbuf_1 wire1557 (.A(net1558),
    .X(net1557));
 sky130_fd_sc_hd__buf_1 wire1558 (.A(net1559),
    .X(net1558));
 sky130_fd_sc_hd__buf_1 wire1559 (.A(_06509_),
    .X(net1559));
 sky130_fd_sc_hd__clkbuf_2 wire1560 (.A(_06292_),
    .X(net1560));
 sky130_fd_sc_hd__buf_1 wire1561 (.A(_06175_),
    .X(net1561));
 sky130_fd_sc_hd__clkbuf_1 wire1562 (.A(_05973_),
    .X(net1562));
 sky130_fd_sc_hd__clkbuf_2 wire1563 (.A(_05909_),
    .X(net1563));
 sky130_fd_sc_hd__clkbuf_1 wire1564 (.A(net1565),
    .X(net1564));
 sky130_fd_sc_hd__clkbuf_1 wire1565 (.A(net1566),
    .X(net1565));
 sky130_fd_sc_hd__buf_1 wire1566 (.A(net1567),
    .X(net1566));
 sky130_fd_sc_hd__buf_1 wire1567 (.A(_05764_),
    .X(net1567));
 sky130_fd_sc_hd__buf_1 wire1568 (.A(net1569),
    .X(net1568));
 sky130_fd_sc_hd__clkbuf_1 wire1569 (.A(net1570),
    .X(net1569));
 sky130_fd_sc_hd__buf_1 wire1570 (.A(_05764_),
    .X(net1570));
 sky130_fd_sc_hd__buf_1 wire1571 (.A(_05686_),
    .X(net1571));
 sky130_fd_sc_hd__buf_1 wire1572 (.A(_05578_),
    .X(net1572));
 sky130_fd_sc_hd__clkbuf_1 wire1573 (.A(net1574),
    .X(net1573));
 sky130_fd_sc_hd__buf_1 wire1574 (.A(_05577_),
    .X(net1574));
 sky130_fd_sc_hd__clkbuf_1 wire1575 (.A(net1576),
    .X(net1575));
 sky130_fd_sc_hd__clkbuf_1 wire1576 (.A(_05555_),
    .X(net1576));
 sky130_fd_sc_hd__buf_1 wire1577 (.A(net1578),
    .X(net1577));
 sky130_fd_sc_hd__buf_1 wire1578 (.A(net1579),
    .X(net1578));
 sky130_fd_sc_hd__buf_1 wire1579 (.A(net1580),
    .X(net1579));
 sky130_fd_sc_hd__buf_1 max_length1580 (.A(net1581),
    .X(net1580));
 sky130_fd_sc_hd__clkbuf_1 wire1581 (.A(net1582),
    .X(net1581));
 sky130_fd_sc_hd__buf_1 wire1582 (.A(_05555_),
    .X(net1582));
 sky130_fd_sc_hd__clkbuf_2 wire1583 (.A(net1584),
    .X(net1583));
 sky130_fd_sc_hd__buf_1 wire1584 (.A(_05504_),
    .X(net1584));
 sky130_fd_sc_hd__buf_1 wire1585 (.A(_05387_),
    .X(net1585));
 sky130_fd_sc_hd__buf_1 wire1586 (.A(net1587),
    .X(net1586));
 sky130_fd_sc_hd__buf_1 wire1587 (.A(net1588),
    .X(net1587));
 sky130_fd_sc_hd__buf_1 wire1588 (.A(net1589),
    .X(net1588));
 sky130_fd_sc_hd__buf_1 wire1589 (.A(net1591),
    .X(net1589));
 sky130_fd_sc_hd__buf_1 wire1590 (.A(net1591),
    .X(net1590));
 sky130_fd_sc_hd__buf_1 wire1591 (.A(_05293_),
    .X(net1591));
 sky130_fd_sc_hd__buf_1 max_length1592 (.A(_05293_),
    .X(net1592));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1593 (.A(_05215_),
    .X(net1593));
 sky130_fd_sc_hd__buf_1 wire1594 (.A(net1595),
    .X(net1594));
 sky130_fd_sc_hd__clkbuf_1 wire1595 (.A(_05135_),
    .X(net1595));
 sky130_fd_sc_hd__buf_1 wire1596 (.A(_05132_),
    .X(net1596));
 sky130_fd_sc_hd__buf_1 wire1597 (.A(_05132_),
    .X(net1597));
 sky130_fd_sc_hd__clkbuf_2 wire1598 (.A(net1599),
    .X(net1598));
 sky130_fd_sc_hd__clkbuf_1 wire1599 (.A(net1600),
    .X(net1599));
 sky130_fd_sc_hd__clkbuf_1 wire1600 (.A(net1601),
    .X(net1600));
 sky130_fd_sc_hd__buf_1 wire1601 (.A(net1602),
    .X(net1601));
 sky130_fd_sc_hd__buf_1 wire1602 (.A(net1603),
    .X(net1602));
 sky130_fd_sc_hd__buf_1 max_length1603 (.A(_05057_),
    .X(net1603));
 sky130_fd_sc_hd__buf_1 wire1604 (.A(_05037_),
    .X(net1604));
 sky130_fd_sc_hd__buf_1 wire1605 (.A(net1606),
    .X(net1605));
 sky130_fd_sc_hd__buf_1 wire1606 (.A(net1607),
    .X(net1606));
 sky130_fd_sc_hd__clkbuf_1 wire1607 (.A(net1608),
    .X(net1607));
 sky130_fd_sc_hd__buf_1 wire1608 (.A(net1609),
    .X(net1608));
 sky130_fd_sc_hd__clkbuf_1 wire1609 (.A(_05015_),
    .X(net1609));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length1610 (.A(_05015_),
    .X(net1610));
 sky130_fd_sc_hd__clkbuf_2 wire1611 (.A(net1612),
    .X(net1611));
 sky130_fd_sc_hd__clkbuf_1 wire1612 (.A(net1613),
    .X(net1612));
 sky130_fd_sc_hd__clkbuf_1 wire1613 (.A(net1614),
    .X(net1613));
 sky130_fd_sc_hd__clkbuf_1 wire1614 (.A(_04977_),
    .X(net1614));
 sky130_fd_sc_hd__buf_1 wire1615 (.A(_04920_),
    .X(net1615));
 sky130_fd_sc_hd__buf_1 wire1616 (.A(net1617),
    .X(net1616));
 sky130_fd_sc_hd__buf_1 max_length1617 (.A(_04920_),
    .X(net1617));
 sky130_fd_sc_hd__clkbuf_1 max_length1618 (.A(_04901_),
    .X(net1618));
 sky130_fd_sc_hd__buf_1 wire1619 (.A(net1620),
    .X(net1619));
 sky130_fd_sc_hd__buf_1 max_length1620 (.A(_04901_),
    .X(net1620));
 sky130_fd_sc_hd__buf_1 wire1621 (.A(net1626),
    .X(net1621));
 sky130_fd_sc_hd__buf_1 wire1622 (.A(net1623),
    .X(net1622));
 sky130_fd_sc_hd__clkbuf_1 wire1623 (.A(net1624),
    .X(net1623));
 sky130_fd_sc_hd__buf_1 wire1624 (.A(net1625),
    .X(net1624));
 sky130_fd_sc_hd__buf_1 wire1625 (.A(_04860_),
    .X(net1625));
 sky130_fd_sc_hd__buf_1 max_length1626 (.A(_04860_),
    .X(net1626));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1627 (.A(_04785_),
    .X(net1627));
 sky130_fd_sc_hd__buf_1 wire1628 (.A(_04785_),
    .X(net1628));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1629 (.A(_04780_),
    .X(net1629));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1630 (.A(_04780_),
    .X(net1630));
 sky130_fd_sc_hd__buf_1 wire1631 (.A(net1632),
    .X(net1631));
 sky130_fd_sc_hd__buf_1 wire1632 (.A(_04752_),
    .X(net1632));
 sky130_fd_sc_hd__buf_1 wire1633 (.A(_04752_),
    .X(net1633));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length1634 (.A(net1635),
    .X(net1634));
 sky130_fd_sc_hd__buf_1 wire1635 (.A(_04734_),
    .X(net1635));
 sky130_fd_sc_hd__clkbuf_2 wire1636 (.A(net1637),
    .X(net1636));
 sky130_fd_sc_hd__buf_1 wire1637 (.A(_04701_),
    .X(net1637));
 sky130_fd_sc_hd__buf_1 wire1638 (.A(net1639),
    .X(net1638));
 sky130_fd_sc_hd__clkbuf_1 wire1639 (.A(_04589_),
    .X(net1639));
 sky130_fd_sc_hd__buf_1 wire1640 (.A(net1641),
    .X(net1640));
 sky130_fd_sc_hd__clkbuf_1 wire1641 (.A(_04554_),
    .X(net1641));
 sky130_fd_sc_hd__buf_1 wire1642 (.A(_04542_),
    .X(net1642));
 sky130_fd_sc_hd__buf_1 wire1643 (.A(_04529_),
    .X(net1643));
 sky130_fd_sc_hd__buf_1 max_length1644 (.A(_04529_),
    .X(net1644));
 sky130_fd_sc_hd__buf_1 max_length1645 (.A(net1646),
    .X(net1645));
 sky130_fd_sc_hd__buf_1 wire1646 (.A(_04509_),
    .X(net1646));
 sky130_fd_sc_hd__buf_1 wire1647 (.A(_04507_),
    .X(net1647));
 sky130_fd_sc_hd__buf_1 wire1648 (.A(_04507_),
    .X(net1648));
 sky130_fd_sc_hd__clkbuf_2 wire1649 (.A(net1650),
    .X(net1649));
 sky130_fd_sc_hd__buf_2 wire1650 (.A(_04283_),
    .X(net1650));
 sky130_fd_sc_hd__clkbuf_4 wire1651 (.A(_04281_),
    .X(net1651));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1652 (.A(_04219_),
    .X(net1652));
 sky130_fd_sc_hd__buf_1 wire1653 (.A(_04149_),
    .X(net1653));
 sky130_fd_sc_hd__buf_1 wire1654 (.A(_04141_),
    .X(net1654));
 sky130_fd_sc_hd__buf_1 wire1655 (.A(_04139_),
    .X(net1655));
 sky130_fd_sc_hd__buf_1 wire1656 (.A(_04093_),
    .X(net1656));
 sky130_fd_sc_hd__buf_1 wire1657 (.A(_04085_),
    .X(net1657));
 sky130_fd_sc_hd__buf_1 wire1658 (.A(_04011_),
    .X(net1658));
 sky130_fd_sc_hd__buf_1 max_cap1659 (.A(_03706_),
    .X(net1659));
 sky130_fd_sc_hd__buf_1 wire1660 (.A(_03693_),
    .X(net1660));
 sky130_fd_sc_hd__clkbuf_1 wire1661 (.A(_03631_),
    .X(net1661));
 sky130_fd_sc_hd__buf_1 wire1662 (.A(_03599_),
    .X(net1662));
 sky130_fd_sc_hd__clkbuf_1 wire1663 (.A(net1664),
    .X(net1663));
 sky130_fd_sc_hd__clkbuf_1 wire1664 (.A(net1665),
    .X(net1664));
 sky130_fd_sc_hd__clkbuf_1 max_length1665 (.A(_03575_),
    .X(net1665));
 sky130_fd_sc_hd__buf_1 wire1666 (.A(_03505_),
    .X(net1666));
 sky130_fd_sc_hd__clkbuf_2 wire1667 (.A(net1668),
    .X(net1667));
 sky130_fd_sc_hd__clkbuf_1 wire1668 (.A(net1669),
    .X(net1668));
 sky130_fd_sc_hd__clkbuf_1 wire1669 (.A(_03366_),
    .X(net1669));
 sky130_fd_sc_hd__clkbuf_2 wire1670 (.A(net1671),
    .X(net1670));
 sky130_fd_sc_hd__clkbuf_1 wire1671 (.A(net1672),
    .X(net1671));
 sky130_fd_sc_hd__clkbuf_1 wire1672 (.A(net1673),
    .X(net1672));
 sky130_fd_sc_hd__clkbuf_1 wire1673 (.A(_03364_),
    .X(net1673));
 sky130_fd_sc_hd__buf_1 wire1674 (.A(_03214_),
    .X(net1674));
 sky130_fd_sc_hd__clkbuf_2 wire1675 (.A(_03185_),
    .X(net1675));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1676 (.A(_03004_),
    .X(net1676));
 sky130_fd_sc_hd__buf_1 wire1677 (.A(_02983_),
    .X(net1677));
 sky130_fd_sc_hd__buf_1 wire1678 (.A(_02931_),
    .X(net1678));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1679 (.A(net1680),
    .X(net1679));
 sky130_fd_sc_hd__clkbuf_2 wire1680 (.A(net1681),
    .X(net1680));
 sky130_fd_sc_hd__clkbuf_2 wire1681 (.A(net1682),
    .X(net1681));
 sky130_fd_sc_hd__clkbuf_1 wire1682 (.A(net1683),
    .X(net1682));
 sky130_fd_sc_hd__clkbuf_1 wire1683 (.A(net1684),
    .X(net1683));
 sky130_fd_sc_hd__clkbuf_1 wire1684 (.A(net1685),
    .X(net1684));
 sky130_fd_sc_hd__clkbuf_1 wire1685 (.A(net1686),
    .X(net1685));
 sky130_fd_sc_hd__clkbuf_1 wire1686 (.A(net1687),
    .X(net1686));
 sky130_fd_sc_hd__buf_1 wire1687 (.A(_02695_),
    .X(net1687));
 sky130_fd_sc_hd__clkbuf_2 wire1688 (.A(net1689),
    .X(net1688));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1689 (.A(net1690),
    .X(net1689));
 sky130_fd_sc_hd__buf_1 wire1690 (.A(net1691),
    .X(net1690));
 sky130_fd_sc_hd__clkbuf_1 wire1691 (.A(net1692),
    .X(net1691));
 sky130_fd_sc_hd__clkbuf_1 wire1692 (.A(net1693),
    .X(net1692));
 sky130_fd_sc_hd__clkbuf_1 wire1693 (.A(net1694),
    .X(net1693));
 sky130_fd_sc_hd__clkbuf_1 wire1694 (.A(net1695),
    .X(net1694));
 sky130_fd_sc_hd__clkbuf_1 wire1695 (.A(net1696),
    .X(net1695));
 sky130_fd_sc_hd__buf_1 wire1696 (.A(_02662_),
    .X(net1696));
 sky130_fd_sc_hd__clkbuf_1 wire1697 (.A(net1698),
    .X(net1697));
 sky130_fd_sc_hd__buf_1 wire1698 (.A(_02568_),
    .X(net1698));
 sky130_fd_sc_hd__buf_1 wire1699 (.A(net1700),
    .X(net1699));
 sky130_fd_sc_hd__buf_1 wire1700 (.A(net1701),
    .X(net1700));
 sky130_fd_sc_hd__buf_1 wire1701 (.A(_02522_),
    .X(net1701));
 sky130_fd_sc_hd__buf_1 wire1702 (.A(_02297_),
    .X(net1702));
 sky130_fd_sc_hd__buf_1 wire1703 (.A(_02231_),
    .X(net1703));
 sky130_fd_sc_hd__buf_1 wire1704 (.A(net1705),
    .X(net1704));
 sky130_fd_sc_hd__clkbuf_1 wire1705 (.A(_02223_),
    .X(net1705));
 sky130_fd_sc_hd__clkbuf_2 wire1706 (.A(net1707),
    .X(net1706));
 sky130_fd_sc_hd__clkbuf_1 wire1707 (.A(_02206_),
    .X(net1707));
 sky130_fd_sc_hd__buf_1 wire1708 (.A(net1709),
    .X(net1708));
 sky130_fd_sc_hd__clkbuf_1 wire1709 (.A(_02154_),
    .X(net1709));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1710 (.A(net1711),
    .X(net1710));
 sky130_fd_sc_hd__clkbuf_1 wire1711 (.A(_02063_),
    .X(net1711));
 sky130_fd_sc_hd__buf_1 wire1712 (.A(_02059_),
    .X(net1712));
 sky130_fd_sc_hd__buf_1 wire1713 (.A(_01961_),
    .X(net1713));
 sky130_fd_sc_hd__buf_1 wire1714 (.A(_01939_),
    .X(net1714));
 sky130_fd_sc_hd__buf_1 max_length1715 (.A(net1716),
    .X(net1715));
 sky130_fd_sc_hd__buf_1 wire1716 (.A(_01887_),
    .X(net1716));
 sky130_fd_sc_hd__buf_1 wire1717 (.A(_01887_),
    .X(net1717));
 sky130_fd_sc_hd__buf_1 wire1718 (.A(_01874_),
    .X(net1718));
 sky130_fd_sc_hd__buf_1 wire1719 (.A(_01843_),
    .X(net1719));
 sky130_fd_sc_hd__buf_1 wire1720 (.A(_01700_),
    .X(net1720));
 sky130_fd_sc_hd__buf_1 wire1721 (.A(_01597_),
    .X(net1721));
 sky130_fd_sc_hd__buf_1 wire1722 (.A(_01568_),
    .X(net1722));
 sky130_fd_sc_hd__clkbuf_1 wire1723 (.A(_01539_),
    .X(net1723));
 sky130_fd_sc_hd__clkbuf_1 max_length1724 (.A(_01539_),
    .X(net1724));
 sky130_fd_sc_hd__buf_1 wire1725 (.A(_01497_),
    .X(net1725));
 sky130_fd_sc_hd__buf_1 wire1726 (.A(_01465_),
    .X(net1726));
 sky130_fd_sc_hd__buf_1 wire1727 (.A(_01461_),
    .X(net1727));
 sky130_fd_sc_hd__buf_1 wire1728 (.A(_01388_),
    .X(net1728));
 sky130_fd_sc_hd__buf_1 wire1729 (.A(_01358_),
    .X(net1729));
 sky130_fd_sc_hd__buf_1 wire1730 (.A(_01272_),
    .X(net1730));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1731 (.A(_01048_),
    .X(net1731));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1732 (.A(net1733),
    .X(net1732));
 sky130_fd_sc_hd__clkbuf_1 wire1733 (.A(_01006_),
    .X(net1733));
 sky130_fd_sc_hd__clkbuf_2 wire1734 (.A(_00958_),
    .X(net1734));
 sky130_fd_sc_hd__buf_1 wire1735 (.A(_00839_),
    .X(net1735));
 sky130_fd_sc_hd__buf_1 wire1736 (.A(_00836_),
    .X(net1736));
 sky130_fd_sc_hd__clkbuf_2 wire1737 (.A(_00832_),
    .X(net1737));
 sky130_fd_sc_hd__buf_1 wire1738 (.A(_12418_),
    .X(net1738));
 sky130_fd_sc_hd__buf_1 wire1739 (.A(_12408_),
    .X(net1739));
 sky130_fd_sc_hd__clkbuf_2 wire1740 (.A(net1741),
    .X(net1740));
 sky130_fd_sc_hd__clkbuf_1 wire1741 (.A(_12365_),
    .X(net1741));
 sky130_fd_sc_hd__buf_1 wire1742 (.A(net1743),
    .X(net1742));
 sky130_fd_sc_hd__clkbuf_1 wire1743 (.A(net1744),
    .X(net1743));
 sky130_fd_sc_hd__clkbuf_1 wire1744 (.A(_12354_),
    .X(net1744));
 sky130_fd_sc_hd__clkbuf_2 wire1745 (.A(net1746),
    .X(net1745));
 sky130_fd_sc_hd__clkbuf_1 wire1746 (.A(_12341_),
    .X(net1746));
 sky130_fd_sc_hd__buf_1 wire1747 (.A(net1748),
    .X(net1747));
 sky130_fd_sc_hd__clkbuf_1 wire1748 (.A(_11644_),
    .X(net1748));
 sky130_fd_sc_hd__buf_1 wire1749 (.A(net1750),
    .X(net1749));
 sky130_fd_sc_hd__clkbuf_1 wire1750 (.A(_11464_),
    .X(net1750));
 sky130_fd_sc_hd__buf_1 wire1751 (.A(_11322_),
    .X(net1751));
 sky130_fd_sc_hd__clkbuf_1 wire1752 (.A(_11172_),
    .X(net1752));
 sky130_fd_sc_hd__buf_1 wire1753 (.A(net1754),
    .X(net1753));
 sky130_fd_sc_hd__clkbuf_1 wire1754 (.A(net1755),
    .X(net1754));
 sky130_fd_sc_hd__clkbuf_1 wire1755 (.A(_11087_),
    .X(net1755));
 sky130_fd_sc_hd__buf_1 wire1756 (.A(_10932_),
    .X(net1756));
 sky130_fd_sc_hd__buf_1 wire1757 (.A(_10921_),
    .X(net1757));
 sky130_fd_sc_hd__buf_1 wire1758 (.A(_10902_),
    .X(net1758));
 sky130_fd_sc_hd__clkbuf_1 wire1759 (.A(_10848_),
    .X(net1759));
 sky130_fd_sc_hd__buf_1 wire1760 (.A(net1761),
    .X(net1760));
 sky130_fd_sc_hd__clkbuf_1 wire1761 (.A(_10540_),
    .X(net1761));
 sky130_fd_sc_hd__buf_1 wire1762 (.A(net1763),
    .X(net1762));
 sky130_fd_sc_hd__clkbuf_1 wire1763 (.A(net1764),
    .X(net1763));
 sky130_fd_sc_hd__clkbuf_1 wire1764 (.A(_10428_),
    .X(net1764));
 sky130_fd_sc_hd__clkbuf_1 wire1765 (.A(_10366_),
    .X(net1765));
 sky130_fd_sc_hd__buf_1 wire1766 (.A(_10299_),
    .X(net1766));
 sky130_fd_sc_hd__buf_1 max_length1767 (.A(net1768),
    .X(net1767));
 sky130_fd_sc_hd__buf_1 wire1768 (.A(net1769),
    .X(net1768));
 sky130_fd_sc_hd__clkbuf_1 wire1769 (.A(_10264_),
    .X(net1769));
 sky130_fd_sc_hd__buf_1 wire1770 (.A(net1771),
    .X(net1770));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1771 (.A(net1772),
    .X(net1771));
 sky130_fd_sc_hd__clkbuf_1 max_length1772 (.A(_10264_),
    .X(net1772));
 sky130_fd_sc_hd__buf_1 wire1773 (.A(_10238_),
    .X(net1773));
 sky130_fd_sc_hd__buf_1 wire1774 (.A(_10230_),
    .X(net1774));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1775 (.A(_10153_),
    .X(net1775));
 sky130_fd_sc_hd__buf_1 wire1776 (.A(_10120_),
    .X(net1776));
 sky130_fd_sc_hd__buf_1 wire1777 (.A(_10092_),
    .X(net1777));
 sky130_fd_sc_hd__clkbuf_1 wire1778 (.A(_09981_),
    .X(net1778));
 sky130_fd_sc_hd__buf_1 wire1779 (.A(_09725_),
    .X(net1779));
 sky130_fd_sc_hd__buf_1 wire1780 (.A(_09714_),
    .X(net1780));
 sky130_fd_sc_hd__buf_1 wire1781 (.A(_09658_),
    .X(net1781));
 sky130_fd_sc_hd__clkbuf_1 wire1782 (.A(net1783),
    .X(net1782));
 sky130_fd_sc_hd__clkbuf_1 wire1783 (.A(_09597_),
    .X(net1783));
 sky130_fd_sc_hd__buf_1 wire1784 (.A(net1785),
    .X(net1784));
 sky130_fd_sc_hd__buf_1 wire1785 (.A(net1786),
    .X(net1785));
 sky130_fd_sc_hd__buf_1 wire1786 (.A(net1787),
    .X(net1786));
 sky130_fd_sc_hd__clkbuf_1 max_length1787 (.A(_09597_),
    .X(net1787));
 sky130_fd_sc_hd__buf_1 wire1788 (.A(_09583_),
    .X(net1788));
 sky130_fd_sc_hd__buf_1 wire1789 (.A(net1790),
    .X(net1789));
 sky130_fd_sc_hd__buf_1 wire1790 (.A(_09583_),
    .X(net1790));
 sky130_fd_sc_hd__buf_1 wire1791 (.A(_09538_),
    .X(net1791));
 sky130_fd_sc_hd__clkbuf_1 wire1792 (.A(net1793),
    .X(net1792));
 sky130_fd_sc_hd__clkbuf_1 wire1793 (.A(_09482_),
    .X(net1793));
 sky130_fd_sc_hd__clkbuf_1 wire1794 (.A(_09438_),
    .X(net1794));
 sky130_fd_sc_hd__buf_1 wire1795 (.A(_09210_),
    .X(net1795));
 sky130_fd_sc_hd__buf_1 wire1796 (.A(_09203_),
    .X(net1796));
 sky130_fd_sc_hd__clkbuf_2 wire1797 (.A(net1798),
    .X(net1797));
 sky130_fd_sc_hd__clkbuf_2 wire1798 (.A(_09194_),
    .X(net1798));
 sky130_fd_sc_hd__buf_1 wire1799 (.A(net1800),
    .X(net1799));
 sky130_fd_sc_hd__clkbuf_2 wire1800 (.A(_09190_),
    .X(net1800));
 sky130_fd_sc_hd__clkbuf_2 wire1801 (.A(_09099_),
    .X(net1801));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1802 (.A(net1803),
    .X(net1802));
 sky130_fd_sc_hd__clkbuf_1 wire1803 (.A(_09010_),
    .X(net1803));
 sky130_fd_sc_hd__clkbuf_2 wire1804 (.A(net1805),
    .X(net1804));
 sky130_fd_sc_hd__buf_1 wire1805 (.A(_08974_),
    .X(net1805));
 sky130_fd_sc_hd__buf_1 wire1806 (.A(_08957_),
    .X(net1806));
 sky130_fd_sc_hd__buf_1 wire1807 (.A(net1809),
    .X(net1807));
 sky130_fd_sc_hd__buf_1 wire1808 (.A(net1809),
    .X(net1808));
 sky130_fd_sc_hd__buf_1 wire1809 (.A(_08918_),
    .X(net1809));
 sky130_fd_sc_hd__clkbuf_1 wire1810 (.A(net1811),
    .X(net1810));
 sky130_fd_sc_hd__clkbuf_1 wire1811 (.A(net1812),
    .X(net1811));
 sky130_fd_sc_hd__clkbuf_1 wire1812 (.A(net1813),
    .X(net1812));
 sky130_fd_sc_hd__buf_1 wire1813 (.A(net1814),
    .X(net1813));
 sky130_fd_sc_hd__clkbuf_1 wire1814 (.A(net1815),
    .X(net1814));
 sky130_fd_sc_hd__buf_1 wire1815 (.A(_08915_),
    .X(net1815));
 sky130_fd_sc_hd__clkbuf_1 wire1816 (.A(net1817),
    .X(net1816));
 sky130_fd_sc_hd__buf_1 wire1817 (.A(_08911_),
    .X(net1817));
 sky130_fd_sc_hd__clkbuf_1 max_length1818 (.A(net1819),
    .X(net1818));
 sky130_fd_sc_hd__buf_1 wire1819 (.A(net1820),
    .X(net1819));
 sky130_fd_sc_hd__buf_1 wire1820 (.A(net1821),
    .X(net1820));
 sky130_fd_sc_hd__buf_1 wire1821 (.A(_08911_),
    .X(net1821));
 sky130_fd_sc_hd__buf_1 wire1822 (.A(net1823),
    .X(net1822));
 sky130_fd_sc_hd__clkbuf_1 wire1823 (.A(net1824),
    .X(net1823));
 sky130_fd_sc_hd__buf_1 wire1824 (.A(net1826),
    .X(net1824));
 sky130_fd_sc_hd__buf_1 wire1825 (.A(net1826),
    .X(net1825));
 sky130_fd_sc_hd__buf_1 wire1826 (.A(net1827),
    .X(net1826));
 sky130_fd_sc_hd__buf_1 wire1827 (.A(_08904_),
    .X(net1827));
 sky130_fd_sc_hd__buf_1 wire1828 (.A(_08838_),
    .X(net1828));
 sky130_fd_sc_hd__buf_1 wire1829 (.A(net1831),
    .X(net1829));
 sky130_fd_sc_hd__clkbuf_1 wire1830 (.A(net1831),
    .X(net1830));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1831 (.A(net1833),
    .X(net1831));
 sky130_fd_sc_hd__clkbuf_1 wire1832 (.A(net1833),
    .X(net1832));
 sky130_fd_sc_hd__buf_1 wire1833 (.A(net1834),
    .X(net1833));
 sky130_fd_sc_hd__clkbuf_1 wire1834 (.A(net1835),
    .X(net1834));
 sky130_fd_sc_hd__buf_1 wire1835 (.A(net1836),
    .X(net1835));
 sky130_fd_sc_hd__clkbuf_1 wire1836 (.A(net1837),
    .X(net1836));
 sky130_fd_sc_hd__buf_1 wire1837 (.A(_08819_),
    .X(net1837));
 sky130_fd_sc_hd__clkbuf_1 wire1838 (.A(net1839),
    .X(net1838));
 sky130_fd_sc_hd__clkbuf_1 wire1839 (.A(_08684_),
    .X(net1839));
 sky130_fd_sc_hd__buf_1 wire1840 (.A(_08396_),
    .X(net1840));
 sky130_fd_sc_hd__clkbuf_1 wire1841 (.A(_08253_),
    .X(net1841));
 sky130_fd_sc_hd__buf_1 wire1842 (.A(net1843),
    .X(net1842));
 sky130_fd_sc_hd__clkbuf_1 wire1843 (.A(net1844),
    .X(net1843));
 sky130_fd_sc_hd__clkbuf_1 wire1844 (.A(_07945_),
    .X(net1844));
 sky130_fd_sc_hd__buf_1 wire1845 (.A(_07942_),
    .X(net1845));
 sky130_fd_sc_hd__buf_1 wire1846 (.A(_07901_),
    .X(net1846));
 sky130_fd_sc_hd__clkbuf_1 wire1847 (.A(net1848),
    .X(net1847));
 sky130_fd_sc_hd__buf_1 max_length1848 (.A(net1849),
    .X(net1848));
 sky130_fd_sc_hd__buf_1 wire1849 (.A(_07901_),
    .X(net1849));
 sky130_fd_sc_hd__buf_1 wire1850 (.A(_07811_),
    .X(net1850));
 sky130_fd_sc_hd__buf_1 wire1851 (.A(_07676_),
    .X(net1851));
 sky130_fd_sc_hd__buf_1 wire1852 (.A(_07653_),
    .X(net1852));
 sky130_fd_sc_hd__buf_1 wire1853 (.A(_07621_),
    .X(net1853));
 sky130_fd_sc_hd__buf_1 wire1854 (.A(net1855),
    .X(net1854));
 sky130_fd_sc_hd__clkbuf_1 wire1855 (.A(net1856),
    .X(net1855));
 sky130_fd_sc_hd__clkbuf_1 wire1856 (.A(_07619_),
    .X(net1856));
 sky130_fd_sc_hd__buf_1 wire1857 (.A(net1858),
    .X(net1857));
 sky130_fd_sc_hd__clkbuf_1 wire1858 (.A(_07600_),
    .X(net1858));
 sky130_fd_sc_hd__buf_1 wire1859 (.A(_07578_),
    .X(net1859));
 sky130_fd_sc_hd__buf_1 wire1860 (.A(_07537_),
    .X(net1860));
 sky130_fd_sc_hd__buf_1 wire1861 (.A(net1862),
    .X(net1861));
 sky130_fd_sc_hd__clkbuf_1 wire1862 (.A(net1863),
    .X(net1862));
 sky130_fd_sc_hd__clkbuf_1 wire1863 (.A(_07533_),
    .X(net1863));
 sky130_fd_sc_hd__buf_1 wire1864 (.A(_07491_),
    .X(net1864));
 sky130_fd_sc_hd__buf_1 wire1865 (.A(_07482_),
    .X(net1865));
 sky130_fd_sc_hd__buf_1 wire1866 (.A(net1867),
    .X(net1866));
 sky130_fd_sc_hd__clkbuf_1 wire1867 (.A(_07396_),
    .X(net1867));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1868 (.A(_07392_),
    .X(net1868));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1869 (.A(net1870),
    .X(net1869));
 sky130_fd_sc_hd__clkbuf_1 wire1870 (.A(net1871),
    .X(net1870));
 sky130_fd_sc_hd__clkbuf_1 wire1871 (.A(_07385_),
    .X(net1871));
 sky130_fd_sc_hd__clkbuf_2 wire1872 (.A(net1873),
    .X(net1872));
 sky130_fd_sc_hd__clkbuf_1 wire1873 (.A(net1874),
    .X(net1873));
 sky130_fd_sc_hd__clkbuf_1 wire1874 (.A(_07376_),
    .X(net1874));
 sky130_fd_sc_hd__clkbuf_2 wire1875 (.A(net1876),
    .X(net1875));
 sky130_fd_sc_hd__clkbuf_1 wire1876 (.A(_07363_),
    .X(net1876));
 sky130_fd_sc_hd__buf_1 wire1877 (.A(_07350_),
    .X(net1877));
 sky130_fd_sc_hd__clkbuf_2 wire1878 (.A(_07308_),
    .X(net1878));
 sky130_fd_sc_hd__buf_1 wire1879 (.A(_07290_),
    .X(net1879));
 sky130_fd_sc_hd__clkbuf_2 wire1880 (.A(_07286_),
    .X(net1880));
 sky130_fd_sc_hd__buf_1 wire1881 (.A(_07283_),
    .X(net1881));
 sky130_fd_sc_hd__buf_1 wire1882 (.A(_07271_),
    .X(net1882));
 sky130_fd_sc_hd__buf_1 wire1883 (.A(_07249_),
    .X(net1883));
 sky130_fd_sc_hd__buf_1 wire1884 (.A(net1885),
    .X(net1884));
 sky130_fd_sc_hd__clkbuf_1 wire1885 (.A(_07225_),
    .X(net1885));
 sky130_fd_sc_hd__buf_1 wire1886 (.A(net1887),
    .X(net1886));
 sky130_fd_sc_hd__clkbuf_1 wire1887 (.A(net1888),
    .X(net1887));
 sky130_fd_sc_hd__clkbuf_1 wire1888 (.A(_07220_),
    .X(net1888));
 sky130_fd_sc_hd__buf_1 wire1889 (.A(net1890),
    .X(net1889));
 sky130_fd_sc_hd__clkbuf_1 wire1890 (.A(net1891),
    .X(net1890));
 sky130_fd_sc_hd__clkbuf_1 wire1891 (.A(_07209_),
    .X(net1891));
 sky130_fd_sc_hd__buf_1 wire1892 (.A(_07197_),
    .X(net1892));
 sky130_fd_sc_hd__clkbuf_2 wire1893 (.A(_07188_),
    .X(net1893));
 sky130_fd_sc_hd__clkbuf_2 wire1894 (.A(_07171_),
    .X(net1894));
 sky130_fd_sc_hd__buf_1 wire1895 (.A(_07103_),
    .X(net1895));
 sky130_fd_sc_hd__buf_1 wire1896 (.A(net1897),
    .X(net1896));
 sky130_fd_sc_hd__clkbuf_1 wire1897 (.A(_07068_),
    .X(net1897));
 sky130_fd_sc_hd__clkbuf_2 wire1898 (.A(net1899),
    .X(net1898));
 sky130_fd_sc_hd__clkbuf_1 wire1899 (.A(net1900),
    .X(net1899));
 sky130_fd_sc_hd__clkbuf_1 wire1900 (.A(_07058_),
    .X(net1900));
 sky130_fd_sc_hd__buf_1 wire1901 (.A(_07033_),
    .X(net1901));
 sky130_fd_sc_hd__buf_1 wire1902 (.A(net1903),
    .X(net1902));
 sky130_fd_sc_hd__clkbuf_1 wire1903 (.A(net1904),
    .X(net1903));
 sky130_fd_sc_hd__clkbuf_1 wire1904 (.A(net1905),
    .X(net1904));
 sky130_fd_sc_hd__clkbuf_1 wire1905 (.A(_06991_),
    .X(net1905));
 sky130_fd_sc_hd__clkbuf_1 wire1906 (.A(net1907),
    .X(net1906));
 sky130_fd_sc_hd__clkbuf_1 wire1907 (.A(_06885_),
    .X(net1907));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1908 (.A(_06850_),
    .X(net1908));
 sky130_fd_sc_hd__clkbuf_1 wire1909 (.A(_06846_),
    .X(net1909));
 sky130_fd_sc_hd__clkbuf_1 wire1910 (.A(_06844_),
    .X(net1910));
 sky130_fd_sc_hd__clkbuf_1 wire1911 (.A(net1912),
    .X(net1911));
 sky130_fd_sc_hd__clkbuf_1 wire1912 (.A(net1913),
    .X(net1912));
 sky130_fd_sc_hd__clkbuf_1 wire1913 (.A(net1914),
    .X(net1913));
 sky130_fd_sc_hd__clkbuf_1 wire1914 (.A(_06508_),
    .X(net1914));
 sky130_fd_sc_hd__buf_1 wire1915 (.A(net1916),
    .X(net1915));
 sky130_fd_sc_hd__buf_1 wire1916 (.A(net1917),
    .X(net1916));
 sky130_fd_sc_hd__buf_1 wire1917 (.A(net1918),
    .X(net1917));
 sky130_fd_sc_hd__buf_1 wire1918 (.A(net1919),
    .X(net1918));
 sky130_fd_sc_hd__clkbuf_1 wire1919 (.A(net1920),
    .X(net1919));
 sky130_fd_sc_hd__clkbuf_1 wire1920 (.A(net1921),
    .X(net1920));
 sky130_fd_sc_hd__buf_1 wire1921 (.A(net1922),
    .X(net1921));
 sky130_fd_sc_hd__buf_1 wire1922 (.A(_06508_),
    .X(net1922));
 sky130_fd_sc_hd__buf_1 wire1923 (.A(_05946_),
    .X(net1923));
 sky130_fd_sc_hd__clkbuf_1 wire1924 (.A(net1925),
    .X(net1924));
 sky130_fd_sc_hd__buf_1 wire1925 (.A(_05857_),
    .X(net1925));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1926 (.A(net1927),
    .X(net1926));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1927 (.A(_05857_),
    .X(net1927));
 sky130_fd_sc_hd__buf_1 wire1928 (.A(net1929),
    .X(net1928));
 sky130_fd_sc_hd__buf_1 wire1929 (.A(net1930),
    .X(net1929));
 sky130_fd_sc_hd__buf_1 wire1930 (.A(net1931),
    .X(net1930));
 sky130_fd_sc_hd__buf_1 wire1931 (.A(net1932),
    .X(net1931));
 sky130_fd_sc_hd__clkbuf_1 wire1932 (.A(net1933),
    .X(net1932));
 sky130_fd_sc_hd__buf_1 wire1933 (.A(net1934),
    .X(net1933));
 sky130_fd_sc_hd__clkbuf_1 wire1934 (.A(net1937),
    .X(net1934));
 sky130_fd_sc_hd__clkbuf_1 wire1935 (.A(net1936),
    .X(net1935));
 sky130_fd_sc_hd__clkbuf_1 wire1936 (.A(net1937),
    .X(net1936));
 sky130_fd_sc_hd__buf_1 wire1937 (.A(_05642_),
    .X(net1937));
 sky130_fd_sc_hd__buf_1 wire1938 (.A(net1939),
    .X(net1938));
 sky130_fd_sc_hd__buf_1 wire1939 (.A(net1941),
    .X(net1939));
 sky130_fd_sc_hd__buf_1 wire1940 (.A(net1941),
    .X(net1940));
 sky130_fd_sc_hd__buf_1 wire1941 (.A(_05617_),
    .X(net1941));
 sky130_fd_sc_hd__buf_1 wire1942 (.A(net1943),
    .X(net1942));
 sky130_fd_sc_hd__buf_1 wire1943 (.A(net1944),
    .X(net1943));
 sky130_fd_sc_hd__clkbuf_1 wire1944 (.A(_05608_),
    .X(net1944));
 sky130_fd_sc_hd__buf_1 wire1945 (.A(_05579_),
    .X(net1945));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1946 (.A(_05487_),
    .X(net1946));
 sky130_fd_sc_hd__buf_1 wire1947 (.A(net1948),
    .X(net1947));
 sky130_fd_sc_hd__buf_1 wire1948 (.A(_05287_),
    .X(net1948));
 sky130_fd_sc_hd__buf_1 wire1949 (.A(_05191_),
    .X(net1949));
 sky130_fd_sc_hd__buf_1 wire1950 (.A(net1951),
    .X(net1950));
 sky130_fd_sc_hd__clkbuf_1 max_length1951 (.A(_05134_),
    .X(net1951));
 sky130_fd_sc_hd__buf_1 wire1952 (.A(net1953),
    .X(net1952));
 sky130_fd_sc_hd__buf_1 wire1953 (.A(net1954),
    .X(net1953));
 sky130_fd_sc_hd__buf_1 wire1954 (.A(net1955),
    .X(net1954));
 sky130_fd_sc_hd__buf_1 wire1955 (.A(_05131_),
    .X(net1955));
 sky130_fd_sc_hd__clkbuf_1 wire1956 (.A(_05110_),
    .X(net1956));
 sky130_fd_sc_hd__clkbuf_2 wire1957 (.A(_05064_),
    .X(net1957));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1958 (.A(net1959),
    .X(net1958));
 sky130_fd_sc_hd__buf_1 wire1959 (.A(_05056_),
    .X(net1959));
 sky130_fd_sc_hd__buf_1 wire1960 (.A(_04976_),
    .X(net1960));
 sky130_fd_sc_hd__buf_1 max_length1961 (.A(_04976_),
    .X(net1961));
 sky130_fd_sc_hd__buf_1 wire1962 (.A(net1965),
    .X(net1962));
 sky130_fd_sc_hd__buf_1 wire1963 (.A(net1964),
    .X(net1963));
 sky130_fd_sc_hd__clkbuf_1 max_length1964 (.A(net1965),
    .X(net1964));
 sky130_fd_sc_hd__clkbuf_2 wire1965 (.A(net1966),
    .X(net1965));
 sky130_fd_sc_hd__clkbuf_1 wire1966 (.A(_04965_),
    .X(net1966));
 sky130_fd_sc_hd__buf_1 wire1967 (.A(_04932_),
    .X(net1967));
 sky130_fd_sc_hd__buf_1 wire1968 (.A(_04932_),
    .X(net1968));
 sky130_fd_sc_hd__buf_1 wire1969 (.A(net1970),
    .X(net1969));
 sky130_fd_sc_hd__clkbuf_1 wire1970 (.A(_04926_),
    .X(net1970));
 sky130_fd_sc_hd__buf_1 wire1971 (.A(_04926_),
    .X(net1971));
 sky130_fd_sc_hd__buf_1 wire1972 (.A(net1973),
    .X(net1972));
 sky130_fd_sc_hd__buf_1 wire1973 (.A(_04924_),
    .X(net1973));
 sky130_fd_sc_hd__buf_1 wire1974 (.A(_04924_),
    .X(net1974));
 sky130_fd_sc_hd__buf_1 wire1975 (.A(net1976),
    .X(net1975));
 sky130_fd_sc_hd__buf_1 wire1976 (.A(net1977),
    .X(net1976));
 sky130_fd_sc_hd__clkbuf_1 wire1977 (.A(net1978),
    .X(net1977));
 sky130_fd_sc_hd__buf_1 wire1978 (.A(net1979),
    .X(net1978));
 sky130_fd_sc_hd__buf_1 wire1979 (.A(net1980),
    .X(net1979));
 sky130_fd_sc_hd__clkbuf_1 max_length1980 (.A(_04913_),
    .X(net1980));
 sky130_fd_sc_hd__clkbuf_1 wire1981 (.A(net1985),
    .X(net1981));
 sky130_fd_sc_hd__buf_1 wire1982 (.A(net1983),
    .X(net1982));
 sky130_fd_sc_hd__buf_1 wire1983 (.A(net1984),
    .X(net1983));
 sky130_fd_sc_hd__clkbuf_1 wire1984 (.A(net1986),
    .X(net1984));
 sky130_fd_sc_hd__clkbuf_1 max_length1985 (.A(net1986),
    .X(net1985));
 sky130_fd_sc_hd__buf_1 wire1986 (.A(_04905_),
    .X(net1986));
 sky130_fd_sc_hd__buf_1 wire1987 (.A(net1989),
    .X(net1987));
 sky130_fd_sc_hd__buf_1 wire1988 (.A(net1989),
    .X(net1988));
 sky130_fd_sc_hd__buf_1 wire1989 (.A(net1990),
    .X(net1989));
 sky130_fd_sc_hd__buf_1 wire1990 (.A(_04859_),
    .X(net1990));
 sky130_fd_sc_hd__clkbuf_1 max_length1991 (.A(_04859_),
    .X(net1991));
 sky130_fd_sc_hd__buf_1 wire1992 (.A(net1993),
    .X(net1992));
 sky130_fd_sc_hd__clkbuf_2 wire1993 (.A(_04853_),
    .X(net1993));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire1994 (.A(_04787_),
    .X(net1994));
 sky130_fd_sc_hd__buf_1 wire1995 (.A(_04787_),
    .X(net1995));
 sky130_fd_sc_hd__buf_2 wire1996 (.A(net1997),
    .X(net1996));
 sky130_fd_sc_hd__clkbuf_2 max_length1997 (.A(net1998),
    .X(net1997));
 sky130_fd_sc_hd__buf_1 wire1998 (.A(_04668_),
    .X(net1998));
 sky130_fd_sc_hd__clkbuf_1 wire1999 (.A(_04665_),
    .X(net1999));
 sky130_fd_sc_hd__clkbuf_2 wire2000 (.A(net2001),
    .X(net2000));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2001 (.A(_04643_),
    .X(net2001));
 sky130_fd_sc_hd__clkbuf_1 wire2002 (.A(net2003),
    .X(net2002));
 sky130_fd_sc_hd__clkbuf_2 wire2003 (.A(net2004),
    .X(net2003));
 sky130_fd_sc_hd__clkbuf_1 wire2004 (.A(net2005),
    .X(net2004));
 sky130_fd_sc_hd__clkbuf_1 wire2005 (.A(net2006),
    .X(net2005));
 sky130_fd_sc_hd__clkbuf_1 wire2006 (.A(net2008),
    .X(net2006));
 sky130_fd_sc_hd__buf_1 wire2007 (.A(net2008),
    .X(net2007));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2008 (.A(_04641_),
    .X(net2008));
 sky130_fd_sc_hd__buf_1 wire2009 (.A(net2010),
    .X(net2009));
 sky130_fd_sc_hd__clkbuf_1 wire2010 (.A(_04583_),
    .X(net2010));
 sky130_fd_sc_hd__buf_1 wire2011 (.A(net2012),
    .X(net2011));
 sky130_fd_sc_hd__clkbuf_1 wire2012 (.A(net2013),
    .X(net2012));
 sky130_fd_sc_hd__clkbuf_1 wire2013 (.A(net2014),
    .X(net2013));
 sky130_fd_sc_hd__clkbuf_1 wire2014 (.A(net2015),
    .X(net2014));
 sky130_fd_sc_hd__buf_1 wire2015 (.A(_04535_),
    .X(net2015));
 sky130_fd_sc_hd__buf_1 wire2016 (.A(net2017),
    .X(net2016));
 sky130_fd_sc_hd__buf_1 wire2017 (.A(_04360_),
    .X(net2017));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2018 (.A(_04280_),
    .X(net2018));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2019 (.A(_04217_),
    .X(net2019));
 sky130_fd_sc_hd__buf_1 wire2020 (.A(net2021),
    .X(net2020));
 sky130_fd_sc_hd__buf_1 wire2021 (.A(_04076_),
    .X(net2021));
 sky130_fd_sc_hd__buf_1 wire2022 (.A(net2023),
    .X(net2022));
 sky130_fd_sc_hd__buf_1 wire2023 (.A(_04010_),
    .X(net2023));
 sky130_fd_sc_hd__buf_2 wire2024 (.A(net2025),
    .X(net2024));
 sky130_fd_sc_hd__buf_1 wire2025 (.A(_03963_),
    .X(net2025));
 sky130_fd_sc_hd__buf_1 wire2026 (.A(_02930_),
    .X(net2026));
 sky130_fd_sc_hd__buf_1 wire2027 (.A(_02870_),
    .X(net2027));
 sky130_fd_sc_hd__buf_1 wire2028 (.A(net2029),
    .X(net2028));
 sky130_fd_sc_hd__buf_1 wire2029 (.A(_02870_),
    .X(net2029));
 sky130_fd_sc_hd__clkbuf_1 wire2030 (.A(net2031),
    .X(net2030));
 sky130_fd_sc_hd__clkbuf_1 wire2031 (.A(net2032),
    .X(net2031));
 sky130_fd_sc_hd__clkbuf_1 wire2032 (.A(_02715_),
    .X(net2032));
 sky130_fd_sc_hd__buf_1 wire2033 (.A(net2034),
    .X(net2033));
 sky130_fd_sc_hd__buf_1 wire2034 (.A(_02715_),
    .X(net2034));
 sky130_fd_sc_hd__buf_1 wire2035 (.A(net2036),
    .X(net2035));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2036 (.A(_02694_),
    .X(net2036));
 sky130_fd_sc_hd__buf_1 wire2037 (.A(net2039),
    .X(net2037));
 sky130_fd_sc_hd__buf_1 max_length2038 (.A(net2039),
    .X(net2038));
 sky130_fd_sc_hd__buf_1 wire2039 (.A(_02661_),
    .X(net2039));
 sky130_fd_sc_hd__buf_1 wire2040 (.A(net2041),
    .X(net2040));
 sky130_fd_sc_hd__clkbuf_1 wire2041 (.A(_02559_),
    .X(net2041));
 sky130_fd_sc_hd__buf_1 wire2042 (.A(_02548_),
    .X(net2042));
 sky130_fd_sc_hd__buf_1 max_length2043 (.A(net2044),
    .X(net2043));
 sky130_fd_sc_hd__buf_1 wire2044 (.A(net2045),
    .X(net2044));
 sky130_fd_sc_hd__buf_1 max_length2045 (.A(_02544_),
    .X(net2045));
 sky130_fd_sc_hd__buf_1 max_length2046 (.A(net2047),
    .X(net2046));
 sky130_fd_sc_hd__buf_1 wire2047 (.A(net2048),
    .X(net2047));
 sky130_fd_sc_hd__buf_1 wire2048 (.A(_02524_),
    .X(net2048));
 sky130_fd_sc_hd__buf_1 wire2049 (.A(_02521_),
    .X(net2049));
 sky130_fd_sc_hd__clkbuf_1 max_length2050 (.A(_02521_),
    .X(net2050));
 sky130_fd_sc_hd__buf_1 wire2051 (.A(_02307_),
    .X(net2051));
 sky130_fd_sc_hd__clkbuf_2 wire2052 (.A(net2053),
    .X(net2052));
 sky130_fd_sc_hd__clkbuf_1 wire2053 (.A(net2054),
    .X(net2053));
 sky130_fd_sc_hd__clkbuf_1 wire2054 (.A(_02209_),
    .X(net2054));
 sky130_fd_sc_hd__buf_1 wire2055 (.A(net2056),
    .X(net2055));
 sky130_fd_sc_hd__buf_1 wire2056 (.A(net2057),
    .X(net2056));
 sky130_fd_sc_hd__clkbuf_2 wire2057 (.A(net2058),
    .X(net2057));
 sky130_fd_sc_hd__clkbuf_2 wire2058 (.A(net2059),
    .X(net2058));
 sky130_fd_sc_hd__buf_1 wire2059 (.A(_01894_),
    .X(net2059));
 sky130_fd_sc_hd__clkbuf_2 wire2060 (.A(net2061),
    .X(net2060));
 sky130_fd_sc_hd__clkbuf_1 wire2061 (.A(_01798_),
    .X(net2061));
 sky130_fd_sc_hd__buf_2 wire2062 (.A(net2063),
    .X(net2062));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2063 (.A(_01798_),
    .X(net2063));
 sky130_fd_sc_hd__buf_1 wire2064 (.A(net2066),
    .X(net2064));
 sky130_fd_sc_hd__buf_1 wire2065 (.A(net2066),
    .X(net2065));
 sky130_fd_sc_hd__clkbuf_2 max_length2066 (.A(_01796_),
    .X(net2066));
 sky130_fd_sc_hd__buf_2 wire2067 (.A(_01779_),
    .X(net2067));
 sky130_fd_sc_hd__buf_1 max_length2068 (.A(_01779_),
    .X(net2068));
 sky130_fd_sc_hd__buf_1 wire2069 (.A(_01711_),
    .X(net2069));
 sky130_fd_sc_hd__clkbuf_1 wire2070 (.A(net2071),
    .X(net2070));
 sky130_fd_sc_hd__clkbuf_1 wire2071 (.A(net2072),
    .X(net2071));
 sky130_fd_sc_hd__clkbuf_1 max_length2072 (.A(_01434_),
    .X(net2072));
 sky130_fd_sc_hd__buf_1 wire2073 (.A(_01155_),
    .X(net2073));
 sky130_fd_sc_hd__clkbuf_2 wire2074 (.A(_01046_),
    .X(net2074));
 sky130_fd_sc_hd__buf_1 wire2075 (.A(_01042_),
    .X(net2075));
 sky130_fd_sc_hd__buf_1 wire2076 (.A(_00974_),
    .X(net2076));
 sky130_fd_sc_hd__clkbuf_2 wire2077 (.A(net2078),
    .X(net2077));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2078 (.A(_12503_),
    .X(net2078));
 sky130_fd_sc_hd__clkbuf_2 wire2079 (.A(net2080),
    .X(net2079));
 sky130_fd_sc_hd__clkbuf_1 wire2080 (.A(net2081),
    .X(net2080));
 sky130_fd_sc_hd__clkbuf_1 wire2081 (.A(_12318_),
    .X(net2081));
 sky130_fd_sc_hd__clkbuf_2 wire2082 (.A(net2083),
    .X(net2082));
 sky130_fd_sc_hd__clkbuf_1 wire2083 (.A(_12300_),
    .X(net2083));
 sky130_fd_sc_hd__clkbuf_2 wire2084 (.A(net2085),
    .X(net2084));
 sky130_fd_sc_hd__clkbuf_1 wire2085 (.A(_12294_),
    .X(net2085));
 sky130_fd_sc_hd__buf_1 wire2086 (.A(_12279_),
    .X(net2086));
 sky130_fd_sc_hd__buf_1 wire2087 (.A(net2088),
    .X(net2087));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2088 (.A(_12271_),
    .X(net2088));
 sky130_fd_sc_hd__buf_1 wire2089 (.A(net2090),
    .X(net2089));
 sky130_fd_sc_hd__clkbuf_1 wire2090 (.A(_12204_),
    .X(net2090));
 sky130_fd_sc_hd__buf_1 wire2091 (.A(_12086_),
    .X(net2091));
 sky130_fd_sc_hd__buf_1 wire2092 (.A(_11805_),
    .X(net2092));
 sky130_fd_sc_hd__clkbuf_2 wire2093 (.A(net2094),
    .X(net2093));
 sky130_fd_sc_hd__clkbuf_1 wire2094 (.A(_11802_),
    .X(net2094));
 sky130_fd_sc_hd__buf_1 wire2095 (.A(net2096),
    .X(net2095));
 sky130_fd_sc_hd__buf_1 wire2096 (.A(_11694_),
    .X(net2096));
 sky130_fd_sc_hd__buf_1 wire2097 (.A(net2098),
    .X(net2097));
 sky130_fd_sc_hd__clkbuf_1 wire2098 (.A(_11692_),
    .X(net2098));
 sky130_fd_sc_hd__buf_1 wire2099 (.A(_11591_),
    .X(net2099));
 sky130_fd_sc_hd__clkbuf_2 wire2100 (.A(_11586_),
    .X(net2100));
 sky130_fd_sc_hd__buf_1 wire2101 (.A(net2102),
    .X(net2101));
 sky130_fd_sc_hd__clkbuf_1 wire2102 (.A(_11468_),
    .X(net2102));
 sky130_fd_sc_hd__buf_1 wire2103 (.A(_11402_),
    .X(net2103));
 sky130_fd_sc_hd__clkbuf_2 wire2104 (.A(net2105),
    .X(net2104));
 sky130_fd_sc_hd__clkbuf_1 wire2105 (.A(_11378_),
    .X(net2105));
 sky130_fd_sc_hd__clkbuf_2 wire2106 (.A(_11378_),
    .X(net2106));
 sky130_fd_sc_hd__buf_1 wire2107 (.A(_11157_),
    .X(net2107));
 sky130_fd_sc_hd__buf_1 wire2108 (.A(_11145_),
    .X(net2108));
 sky130_fd_sc_hd__buf_1 wire2109 (.A(_10956_),
    .X(net2109));
 sky130_fd_sc_hd__buf_1 wire2110 (.A(_10953_),
    .X(net2110));
 sky130_fd_sc_hd__buf_1 wire2111 (.A(_10952_),
    .X(net2111));
 sky130_fd_sc_hd__buf_1 wire2112 (.A(_10951_),
    .X(net2112));
 sky130_fd_sc_hd__clkbuf_1 wire2113 (.A(net2114),
    .X(net2113));
 sky130_fd_sc_hd__clkbuf_1 wire2114 (.A(net2115),
    .X(net2114));
 sky130_fd_sc_hd__clkbuf_1 wire2115 (.A(net2116),
    .X(net2115));
 sky130_fd_sc_hd__clkbuf_1 wire2116 (.A(_10887_),
    .X(net2116));
 sky130_fd_sc_hd__buf_1 wire2117 (.A(net2118),
    .X(net2117));
 sky130_fd_sc_hd__clkbuf_1 wire2118 (.A(net2119),
    .X(net2118));
 sky130_fd_sc_hd__clkbuf_1 wire2119 (.A(net2120),
    .X(net2119));
 sky130_fd_sc_hd__clkbuf_1 wire2120 (.A(_10874_),
    .X(net2120));
 sky130_fd_sc_hd__buf_1 wire2121 (.A(net2124),
    .X(net2121));
 sky130_fd_sc_hd__buf_1 max_length2122 (.A(net2123),
    .X(net2122));
 sky130_fd_sc_hd__buf_1 wire2123 (.A(net2124),
    .X(net2123));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2124 (.A(_10771_),
    .X(net2124));
 sky130_fd_sc_hd__buf_1 wire2125 (.A(_10588_),
    .X(net2125));
 sky130_fd_sc_hd__clkbuf_1 wire2126 (.A(_10546_),
    .X(net2126));
 sky130_fd_sc_hd__clkbuf_2 wire2127 (.A(_10481_),
    .X(net2127));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2128 (.A(_10433_),
    .X(net2128));
 sky130_fd_sc_hd__clkbuf_2 wire2129 (.A(_10368_),
    .X(net2129));
 sky130_fd_sc_hd__buf_1 wire2130 (.A(_10363_),
    .X(net2130));
 sky130_fd_sc_hd__clkbuf_2 wire2131 (.A(_10277_),
    .X(net2131));
 sky130_fd_sc_hd__clkbuf_1 wire2132 (.A(net2133),
    .X(net2132));
 sky130_fd_sc_hd__buf_1 wire2133 (.A(net2134),
    .X(net2133));
 sky130_fd_sc_hd__buf_1 wire2134 (.A(net2135),
    .X(net2134));
 sky130_fd_sc_hd__buf_1 wire2135 (.A(net2136),
    .X(net2135));
 sky130_fd_sc_hd__clkbuf_1 wire2136 (.A(net2137),
    .X(net2136));
 sky130_fd_sc_hd__clkbuf_1 wire2137 (.A(_10263_),
    .X(net2137));
 sky130_fd_sc_hd__buf_1 wire2138 (.A(_10112_),
    .X(net2138));
 sky130_fd_sc_hd__buf_1 wire2139 (.A(net2140),
    .X(net2139));
 sky130_fd_sc_hd__clkbuf_1 wire2140 (.A(_09815_),
    .X(net2140));
 sky130_fd_sc_hd__buf_1 wire2141 (.A(_09719_),
    .X(net2141));
 sky130_fd_sc_hd__clkbuf_1 wire2142 (.A(_09706_),
    .X(net2142));
 sky130_fd_sc_hd__clkbuf_2 wire2143 (.A(net2144),
    .X(net2143));
 sky130_fd_sc_hd__clkbuf_1 wire2144 (.A(_09698_),
    .X(net2144));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2145 (.A(_09692_),
    .X(net2145));
 sky130_fd_sc_hd__buf_1 max_length2146 (.A(_09577_),
    .X(net2146));
 sky130_fd_sc_hd__clkbuf_2 wire2147 (.A(net2148),
    .X(net2147));
 sky130_fd_sc_hd__buf_1 wire2148 (.A(net2149),
    .X(net2148));
 sky130_fd_sc_hd__clkbuf_1 wire2149 (.A(net2150),
    .X(net2149));
 sky130_fd_sc_hd__clkbuf_1 wire2150 (.A(_09577_),
    .X(net2150));
 sky130_fd_sc_hd__clkbuf_1 wire2151 (.A(net2152),
    .X(net2151));
 sky130_fd_sc_hd__clkbuf_1 wire2152 (.A(_09503_),
    .X(net2152));
 sky130_fd_sc_hd__buf_1 wire2153 (.A(_09476_),
    .X(net2153));
 sky130_fd_sc_hd__clkbuf_1 max_length2154 (.A(net2155),
    .X(net2154));
 sky130_fd_sc_hd__buf_1 wire2155 (.A(_09429_),
    .X(net2155));
 sky130_fd_sc_hd__buf_1 wire2156 (.A(net2158),
    .X(net2156));
 sky130_fd_sc_hd__buf_1 max_length2157 (.A(net2158),
    .X(net2157));
 sky130_fd_sc_hd__buf_1 wire2158 (.A(_09193_),
    .X(net2158));
 sky130_fd_sc_hd__buf_1 max_length2159 (.A(net2160),
    .X(net2159));
 sky130_fd_sc_hd__clkbuf_2 wire2160 (.A(_09191_),
    .X(net2160));
 sky130_fd_sc_hd__buf_1 wire2161 (.A(net2163),
    .X(net2161));
 sky130_fd_sc_hd__buf_1 wire2162 (.A(net2163),
    .X(net2162));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2163 (.A(_09189_),
    .X(net2163));
 sky130_fd_sc_hd__buf_1 wire2164 (.A(net2165),
    .X(net2164));
 sky130_fd_sc_hd__clkbuf_2 wire2165 (.A(_09185_),
    .X(net2165));
 sky130_fd_sc_hd__buf_1 wire2166 (.A(net2167),
    .X(net2166));
 sky130_fd_sc_hd__clkbuf_1 wire2167 (.A(net2168),
    .X(net2167));
 sky130_fd_sc_hd__buf_1 wire2168 (.A(_09096_),
    .X(net2168));
 sky130_fd_sc_hd__clkbuf_1 wire2169 (.A(_09081_),
    .X(net2169));
 sky130_fd_sc_hd__clkbuf_1 wire2170 (.A(_09070_),
    .X(net2170));
 sky130_fd_sc_hd__clkbuf_2 wire2171 (.A(net2172),
    .X(net2171));
 sky130_fd_sc_hd__buf_1 wire2172 (.A(_08989_),
    .X(net2172));
 sky130_fd_sc_hd__buf_1 wire2173 (.A(_08951_),
    .X(net2173));
 sky130_fd_sc_hd__buf_1 wire2174 (.A(net2175),
    .X(net2174));
 sky130_fd_sc_hd__clkbuf_1 wire2175 (.A(_08899_),
    .X(net2175));
 sky130_fd_sc_hd__buf_1 wire2176 (.A(_08883_),
    .X(net2176));
 sky130_fd_sc_hd__clkbuf_2 wire2177 (.A(_08851_),
    .X(net2177));
 sky130_fd_sc_hd__buf_1 wire2178 (.A(net2179),
    .X(net2178));
 sky130_fd_sc_hd__buf_1 wire2179 (.A(net2180),
    .X(net2179));
 sky130_fd_sc_hd__buf_1 wire2180 (.A(net2181),
    .X(net2180));
 sky130_fd_sc_hd__buf_1 wire2181 (.A(net2188),
    .X(net2181));
 sky130_fd_sc_hd__clkbuf_1 wire2182 (.A(net2183),
    .X(net2182));
 sky130_fd_sc_hd__buf_1 wire2183 (.A(net2184),
    .X(net2183));
 sky130_fd_sc_hd__clkbuf_1 wire2184 (.A(net2185),
    .X(net2184));
 sky130_fd_sc_hd__clkbuf_1 wire2185 (.A(net2186),
    .X(net2185));
 sky130_fd_sc_hd__buf_1 wire2186 (.A(net2187),
    .X(net2186));
 sky130_fd_sc_hd__buf_1 wire2187 (.A(_08841_),
    .X(net2187));
 sky130_fd_sc_hd__clkbuf_1 max_length2188 (.A(_08841_),
    .X(net2188));
 sky130_fd_sc_hd__buf_1 wire2189 (.A(_08833_),
    .X(net2189));
 sky130_fd_sc_hd__buf_1 wire2190 (.A(net2191),
    .X(net2190));
 sky130_fd_sc_hd__buf_1 wire2191 (.A(net2192),
    .X(net2191));
 sky130_fd_sc_hd__buf_1 wire2192 (.A(net2193),
    .X(net2192));
 sky130_fd_sc_hd__clkbuf_1 wire2193 (.A(net2194),
    .X(net2193));
 sky130_fd_sc_hd__clkbuf_1 wire2194 (.A(_08818_),
    .X(net2194));
 sky130_fd_sc_hd__clkbuf_1 wire2195 (.A(net2196),
    .X(net2195));
 sky130_fd_sc_hd__buf_1 wire2196 (.A(net2197),
    .X(net2196));
 sky130_fd_sc_hd__buf_1 wire2197 (.A(net2198),
    .X(net2197));
 sky130_fd_sc_hd__clkbuf_1 wire2198 (.A(net2199),
    .X(net2198));
 sky130_fd_sc_hd__buf_1 wire2199 (.A(net2200),
    .X(net2199));
 sky130_fd_sc_hd__clkbuf_1 wire2200 (.A(net2201),
    .X(net2200));
 sky130_fd_sc_hd__clkbuf_1 max_length2201 (.A(_08818_),
    .X(net2201));
 sky130_fd_sc_hd__buf_1 wire2202 (.A(net2203),
    .X(net2202));
 sky130_fd_sc_hd__clkbuf_1 wire2203 (.A(_08677_),
    .X(net2203));
 sky130_fd_sc_hd__clkbuf_2 wire2204 (.A(_08258_),
    .X(net2204));
 sky130_fd_sc_hd__buf_1 max_length2205 (.A(net2206),
    .X(net2205));
 sky130_fd_sc_hd__buf_1 wire2206 (.A(net2207),
    .X(net2206));
 sky130_fd_sc_hd__clkbuf_1 wire2207 (.A(_08051_),
    .X(net2207));
 sky130_fd_sc_hd__buf_1 max_length2208 (.A(net2209),
    .X(net2208));
 sky130_fd_sc_hd__buf_1 wire2209 (.A(net2210),
    .X(net2209));
 sky130_fd_sc_hd__buf_1 wire2210 (.A(net2211),
    .X(net2210));
 sky130_fd_sc_hd__buf_1 wire2211 (.A(net2212),
    .X(net2211));
 sky130_fd_sc_hd__buf_1 wire2212 (.A(_07990_),
    .X(net2212));
 sky130_fd_sc_hd__clkbuf_1 wire2213 (.A(net2214),
    .X(net2213));
 sky130_fd_sc_hd__buf_1 wire2214 (.A(_07900_),
    .X(net2214));
 sky130_fd_sc_hd__buf_1 wire2215 (.A(_07898_),
    .X(net2215));
 sky130_fd_sc_hd__clkbuf_1 wire2216 (.A(_07896_),
    .X(net2216));
 sky130_fd_sc_hd__buf_1 wire2217 (.A(net2219),
    .X(net2217));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length2218 (.A(net2219),
    .X(net2218));
 sky130_fd_sc_hd__buf_1 wire2219 (.A(net2220),
    .X(net2219));
 sky130_fd_sc_hd__buf_1 wire2220 (.A(_07896_),
    .X(net2220));
 sky130_fd_sc_hd__clkbuf_1 wire2221 (.A(_07810_),
    .X(net2221));
 sky130_fd_sc_hd__buf_1 wire2222 (.A(net2223),
    .X(net2222));
 sky130_fd_sc_hd__clkbuf_2 max_length2223 (.A(net2224),
    .X(net2223));
 sky130_fd_sc_hd__buf_1 wire2224 (.A(_07810_),
    .X(net2224));
 sky130_fd_sc_hd__buf_1 wire2225 (.A(net2226),
    .X(net2225));
 sky130_fd_sc_hd__clkbuf_1 wire2226 (.A(_07788_),
    .X(net2226));
 sky130_fd_sc_hd__buf_1 wire2227 (.A(_07607_),
    .X(net2227));
 sky130_fd_sc_hd__buf_1 wire2228 (.A(_07570_),
    .X(net2228));
 sky130_fd_sc_hd__clkbuf_2 wire2229 (.A(net2230),
    .X(net2229));
 sky130_fd_sc_hd__clkbuf_1 wire2230 (.A(net2231),
    .X(net2230));
 sky130_fd_sc_hd__clkbuf_1 wire2231 (.A(net2232),
    .X(net2231));
 sky130_fd_sc_hd__clkbuf_1 wire2232 (.A(_07394_),
    .X(net2232));
 sky130_fd_sc_hd__buf_1 wire2233 (.A(_07377_),
    .X(net2233));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2234 (.A(net2235),
    .X(net2234));
 sky130_fd_sc_hd__buf_1 max_length2235 (.A(_07377_),
    .X(net2235));
 sky130_fd_sc_hd__clkbuf_1 wire2236 (.A(net2237),
    .X(net2236));
 sky130_fd_sc_hd__clkbuf_1 max_length2237 (.A(net2238),
    .X(net2237));
 sky130_fd_sc_hd__buf_1 wire2238 (.A(net2241),
    .X(net2238));
 sky130_fd_sc_hd__clkbuf_2 wire2239 (.A(net2240),
    .X(net2239));
 sky130_fd_sc_hd__clkbuf_1 wire2240 (.A(_07275_),
    .X(net2240));
 sky130_fd_sc_hd__clkbuf_1 max_length2241 (.A(_07275_),
    .X(net2241));
 sky130_fd_sc_hd__buf_1 wire2242 (.A(_07231_),
    .X(net2242));
 sky130_fd_sc_hd__clkbuf_1 wire2243 (.A(net2244),
    .X(net2243));
 sky130_fd_sc_hd__clkbuf_1 wire2244 (.A(_07156_),
    .X(net2244));
 sky130_fd_sc_hd__clkbuf_2 wire2245 (.A(net2246),
    .X(net2245));
 sky130_fd_sc_hd__buf_1 wire2246 (.A(net2247),
    .X(net2246));
 sky130_fd_sc_hd__clkbuf_1 wire2247 (.A(net2248),
    .X(net2247));
 sky130_fd_sc_hd__clkbuf_1 max_length2248 (.A(_07156_),
    .X(net2248));
 sky130_fd_sc_hd__buf_1 wire2249 (.A(_07130_),
    .X(net2249));
 sky130_fd_sc_hd__buf_1 wire2250 (.A(net2251),
    .X(net2250));
 sky130_fd_sc_hd__buf_1 wire2251 (.A(_07130_),
    .X(net2251));
 sky130_fd_sc_hd__clkbuf_2 wire2252 (.A(net2253),
    .X(net2252));
 sky130_fd_sc_hd__clkbuf_1 wire2253 (.A(net2254),
    .X(net2253));
 sky130_fd_sc_hd__clkbuf_1 wire2254 (.A(net2255),
    .X(net2254));
 sky130_fd_sc_hd__clkbuf_1 wire2255 (.A(_07006_),
    .X(net2255));
 sky130_fd_sc_hd__clkbuf_2 wire2256 (.A(net2257),
    .X(net2256));
 sky130_fd_sc_hd__clkbuf_1 wire2257 (.A(net2258),
    .X(net2257));
 sky130_fd_sc_hd__clkbuf_1 wire2258 (.A(_06980_),
    .X(net2258));
 sky130_fd_sc_hd__clkbuf_1 wire2259 (.A(_06875_),
    .X(net2259));
 sky130_fd_sc_hd__clkbuf_1 wire2260 (.A(_06841_),
    .X(net2260));
 sky130_fd_sc_hd__clkbuf_1 wire2261 (.A(_06837_),
    .X(net2261));
 sky130_fd_sc_hd__clkbuf_2 wire2262 (.A(_06825_),
    .X(net2262));
 sky130_fd_sc_hd__buf_1 max_length2263 (.A(_06825_),
    .X(net2263));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2264 (.A(_06519_),
    .X(net2264));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2265 (.A(net2266),
    .X(net2265));
 sky130_fd_sc_hd__buf_1 wire2266 (.A(net2267),
    .X(net2266));
 sky130_fd_sc_hd__clkbuf_1 wire2267 (.A(net2268),
    .X(net2267));
 sky130_fd_sc_hd__clkbuf_1 wire2268 (.A(net2269),
    .X(net2268));
 sky130_fd_sc_hd__clkbuf_1 wire2269 (.A(net2270),
    .X(net2269));
 sky130_fd_sc_hd__clkbuf_1 wire2270 (.A(net2271),
    .X(net2270));
 sky130_fd_sc_hd__clkbuf_1 wire2271 (.A(net2272),
    .X(net2271));
 sky130_fd_sc_hd__clkbuf_1 wire2272 (.A(net2273),
    .X(net2272));
 sky130_fd_sc_hd__clkbuf_1 wire2273 (.A(net2274),
    .X(net2273));
 sky130_fd_sc_hd__clkbuf_1 wire2274 (.A(net2275),
    .X(net2274));
 sky130_fd_sc_hd__clkbuf_1 wire2275 (.A(net2276),
    .X(net2275));
 sky130_fd_sc_hd__clkbuf_1 wire2276 (.A(net2277),
    .X(net2276));
 sky130_fd_sc_hd__clkbuf_1 max_length2277 (.A(_06517_),
    .X(net2277));
 sky130_fd_sc_hd__buf_2 wire2278 (.A(_06515_),
    .X(net2278));
 sky130_fd_sc_hd__clkbuf_1 wire2279 (.A(net2280),
    .X(net2279));
 sky130_fd_sc_hd__buf_1 wire2280 (.A(net2281),
    .X(net2280));
 sky130_fd_sc_hd__buf_1 wire2281 (.A(net2282),
    .X(net2281));
 sky130_fd_sc_hd__clkbuf_1 wire2282 (.A(net2283),
    .X(net2282));
 sky130_fd_sc_hd__clkbuf_1 max_length2283 (.A(net2284),
    .X(net2283));
 sky130_fd_sc_hd__buf_1 wire2284 (.A(_06507_),
    .X(net2284));
 sky130_fd_sc_hd__clkbuf_1 wire2285 (.A(net2286),
    .X(net2285));
 sky130_fd_sc_hd__clkbuf_1 wire2286 (.A(_06502_),
    .X(net2286));
 sky130_fd_sc_hd__clkbuf_2 max_length2287 (.A(net2288),
    .X(net2287));
 sky130_fd_sc_hd__buf_1 wire2288 (.A(net2289),
    .X(net2288));
 sky130_fd_sc_hd__buf_1 wire2289 (.A(net2290),
    .X(net2289));
 sky130_fd_sc_hd__clkbuf_1 wire2290 (.A(_06502_),
    .X(net2290));
 sky130_fd_sc_hd__buf_1 wire2291 (.A(net2292),
    .X(net2291));
 sky130_fd_sc_hd__buf_1 wire2292 (.A(net2293),
    .X(net2292));
 sky130_fd_sc_hd__buf_1 wire2293 (.A(_05609_),
    .X(net2293));
 sky130_fd_sc_hd__buf_1 wire2294 (.A(net2295),
    .X(net2294));
 sky130_fd_sc_hd__clkbuf_1 wire2295 (.A(_05532_),
    .X(net2295));
 sky130_fd_sc_hd__buf_1 wire2296 (.A(net2297),
    .X(net2296));
 sky130_fd_sc_hd__buf_1 wire2297 (.A(net2298),
    .X(net2297));
 sky130_fd_sc_hd__buf_1 wire2298 (.A(net2299),
    .X(net2298));
 sky130_fd_sc_hd__clkbuf_1 wire2299 (.A(_05420_),
    .X(net2299));
 sky130_fd_sc_hd__clkbuf_1 wire2300 (.A(net2301),
    .X(net2300));
 sky130_fd_sc_hd__buf_1 wire2301 (.A(net2302),
    .X(net2301));
 sky130_fd_sc_hd__buf_1 wire2302 (.A(_05419_),
    .X(net2302));
 sky130_fd_sc_hd__buf_1 wire2303 (.A(_05348_),
    .X(net2303));
 sky130_fd_sc_hd__buf_1 wire2304 (.A(_05189_),
    .X(net2304));
 sky130_fd_sc_hd__buf_1 wire2305 (.A(net2306),
    .X(net2305));
 sky130_fd_sc_hd__clkbuf_1 wire2306 (.A(_05130_),
    .X(net2306));
 sky130_fd_sc_hd__buf_1 wire2307 (.A(net2308),
    .X(net2307));
 sky130_fd_sc_hd__buf_1 wire2308 (.A(net2309),
    .X(net2308));
 sky130_fd_sc_hd__buf_1 wire2309 (.A(net2310),
    .X(net2309));
 sky130_fd_sc_hd__buf_1 wire2310 (.A(_05129_),
    .X(net2310));
 sky130_fd_sc_hd__buf_1 wire2311 (.A(net2312),
    .X(net2311));
 sky130_fd_sc_hd__buf_1 wire2312 (.A(net2313),
    .X(net2312));
 sky130_fd_sc_hd__clkbuf_1 wire2313 (.A(net2314),
    .X(net2313));
 sky130_fd_sc_hd__clkbuf_1 wire2314 (.A(net2315),
    .X(net2314));
 sky130_fd_sc_hd__buf_1 wire2315 (.A(net2316),
    .X(net2315));
 sky130_fd_sc_hd__buf_1 max_length2316 (.A(_05035_),
    .X(net2316));
 sky130_fd_sc_hd__buf_1 wire2317 (.A(net2318),
    .X(net2317));
 sky130_fd_sc_hd__buf_1 wire2318 (.A(net2319),
    .X(net2318));
 sky130_fd_sc_hd__buf_1 wire2319 (.A(net2320),
    .X(net2319));
 sky130_fd_sc_hd__buf_1 wire2320 (.A(_04975_),
    .X(net2320));
 sky130_fd_sc_hd__buf_1 wire2321 (.A(net2322),
    .X(net2321));
 sky130_fd_sc_hd__buf_1 wire2322 (.A(net2323),
    .X(net2322));
 sky130_fd_sc_hd__buf_1 wire2323 (.A(net2324),
    .X(net2323));
 sky130_fd_sc_hd__buf_1 wire2324 (.A(_04974_),
    .X(net2324));
 sky130_fd_sc_hd__buf_1 wire2325 (.A(net2326),
    .X(net2325));
 sky130_fd_sc_hd__buf_1 wire2326 (.A(net2327),
    .X(net2326));
 sky130_fd_sc_hd__buf_1 wire2327 (.A(net2328),
    .X(net2327));
 sky130_fd_sc_hd__clkbuf_1 wire2328 (.A(net2329),
    .X(net2328));
 sky130_fd_sc_hd__buf_1 wire2329 (.A(_04959_),
    .X(net2329));
 sky130_fd_sc_hd__buf_1 wire2330 (.A(net2331),
    .X(net2330));
 sky130_fd_sc_hd__buf_1 max_length2331 (.A(net2332),
    .X(net2331));
 sky130_fd_sc_hd__buf_1 wire2332 (.A(net2333),
    .X(net2332));
 sky130_fd_sc_hd__clkbuf_1 wire2333 (.A(net2334),
    .X(net2333));
 sky130_fd_sc_hd__buf_1 wire2334 (.A(_04957_),
    .X(net2334));
 sky130_fd_sc_hd__buf_1 wire2335 (.A(net2336),
    .X(net2335));
 sky130_fd_sc_hd__buf_1 wire2336 (.A(net2337),
    .X(net2336));
 sky130_fd_sc_hd__clkbuf_1 wire2337 (.A(_04931_),
    .X(net2337));
 sky130_fd_sc_hd__buf_1 wire2338 (.A(net2339),
    .X(net2338));
 sky130_fd_sc_hd__buf_1 wire2339 (.A(_04930_),
    .X(net2339));
 sky130_fd_sc_hd__clkbuf_1 wire2340 (.A(_04930_),
    .X(net2340));
 sky130_fd_sc_hd__buf_1 wire2341 (.A(net2342),
    .X(net2341));
 sky130_fd_sc_hd__buf_1 wire2342 (.A(net2343),
    .X(net2342));
 sky130_fd_sc_hd__clkbuf_1 wire2343 (.A(_04925_),
    .X(net2343));
 sky130_fd_sc_hd__buf_1 wire2344 (.A(net2345),
    .X(net2344));
 sky130_fd_sc_hd__buf_1 wire2345 (.A(_04923_),
    .X(net2345));
 sky130_fd_sc_hd__buf_1 max_length2346 (.A(net2347),
    .X(net2346));
 sky130_fd_sc_hd__buf_1 wire2347 (.A(net2348),
    .X(net2347));
 sky130_fd_sc_hd__buf_1 wire2348 (.A(net2349),
    .X(net2348));
 sky130_fd_sc_hd__clkbuf_1 wire2349 (.A(_04918_),
    .X(net2349));
 sky130_fd_sc_hd__buf_1 max_length2350 (.A(net2351),
    .X(net2350));
 sky130_fd_sc_hd__buf_1 wire2351 (.A(net2352),
    .X(net2351));
 sky130_fd_sc_hd__clkbuf_1 wire2352 (.A(net2353),
    .X(net2352));
 sky130_fd_sc_hd__buf_1 wire2353 (.A(_04917_),
    .X(net2353));
 sky130_fd_sc_hd__buf_1 wire2354 (.A(net2355),
    .X(net2354));
 sky130_fd_sc_hd__clkbuf_1 wire2355 (.A(_04912_),
    .X(net2355));
 sky130_fd_sc_hd__buf_1 wire2356 (.A(net2357),
    .X(net2356));
 sky130_fd_sc_hd__buf_1 wire2357 (.A(net2358),
    .X(net2357));
 sky130_fd_sc_hd__clkbuf_1 wire2358 (.A(_04910_),
    .X(net2358));
 sky130_fd_sc_hd__clkbuf_1 wire2359 (.A(net2363),
    .X(net2359));
 sky130_fd_sc_hd__buf_1 wire2360 (.A(net2361),
    .X(net2360));
 sky130_fd_sc_hd__buf_1 wire2361 (.A(net2362),
    .X(net2361));
 sky130_fd_sc_hd__clkbuf_1 wire2362 (.A(net2364),
    .X(net2362));
 sky130_fd_sc_hd__clkbuf_1 max_length2363 (.A(net2364),
    .X(net2363));
 sky130_fd_sc_hd__buf_1 wire2364 (.A(_04907_),
    .X(net2364));
 sky130_fd_sc_hd__buf_1 wire2365 (.A(net2366),
    .X(net2365));
 sky130_fd_sc_hd__clkbuf_1 wire2366 (.A(net2367),
    .X(net2366));
 sky130_fd_sc_hd__buf_1 wire2367 (.A(_04899_),
    .X(net2367));
 sky130_fd_sc_hd__buf_1 wire2368 (.A(net2369),
    .X(net2368));
 sky130_fd_sc_hd__clkbuf_1 wire2369 (.A(net2370),
    .X(net2369));
 sky130_fd_sc_hd__buf_1 max_length2370 (.A(_04895_),
    .X(net2370));
 sky130_fd_sc_hd__clkbuf_1 wire2371 (.A(net2372),
    .X(net2371));
 sky130_fd_sc_hd__clkbuf_1 wire2372 (.A(net2373),
    .X(net2372));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2373 (.A(net2376),
    .X(net2373));
 sky130_fd_sc_hd__buf_1 wire2374 (.A(net2375),
    .X(net2374));
 sky130_fd_sc_hd__buf_1 wire2375 (.A(net2376),
    .X(net2375));
 sky130_fd_sc_hd__buf_1 wire2376 (.A(net2377),
    .X(net2376));
 sky130_fd_sc_hd__clkbuf_1 wire2377 (.A(net2378),
    .X(net2377));
 sky130_fd_sc_hd__buf_1 wire2378 (.A(_04891_),
    .X(net2378));
 sky130_fd_sc_hd__buf_1 wire2379 (.A(net2380),
    .X(net2379));
 sky130_fd_sc_hd__buf_1 wire2380 (.A(net2381),
    .X(net2380));
 sky130_fd_sc_hd__buf_1 wire2381 (.A(_00006_),
    .X(net2381));
 sky130_fd_sc_hd__buf_1 wire2382 (.A(_00011_),
    .X(net2382));
 sky130_fd_sc_hd__clkbuf_1 max_length2383 (.A(net2384),
    .X(net2383));
 sky130_fd_sc_hd__buf_1 wire2384 (.A(_00011_),
    .X(net2384));
 sky130_fd_sc_hd__buf_1 wire2385 (.A(_04858_),
    .X(net2385));
 sky130_fd_sc_hd__clkbuf_1 wire2386 (.A(net2387),
    .X(net2386));
 sky130_fd_sc_hd__clkbuf_1 wire2387 (.A(net2388),
    .X(net2387));
 sky130_fd_sc_hd__buf_1 wire2388 (.A(net2389),
    .X(net2388));
 sky130_fd_sc_hd__buf_1 wire2389 (.A(net2390),
    .X(net2389));
 sky130_fd_sc_hd__buf_1 wire2390 (.A(_04858_),
    .X(net2390));
 sky130_fd_sc_hd__buf_1 wire2391 (.A(_04852_),
    .X(net2391));
 sky130_fd_sc_hd__buf_1 wire2392 (.A(net2393),
    .X(net2392));
 sky130_fd_sc_hd__clkbuf_2 wire2393 (.A(_04850_),
    .X(net2393));
 sky130_fd_sc_hd__buf_1 wire2394 (.A(net2395),
    .X(net2394));
 sky130_fd_sc_hd__buf_1 wire2395 (.A(net2396),
    .X(net2395));
 sky130_fd_sc_hd__buf_1 wire2396 (.A(_04753_),
    .X(net2396));
 sky130_fd_sc_hd__clkbuf_2 wire2397 (.A(net2398),
    .X(net2397));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2398 (.A(_04664_),
    .X(net2398));
 sky130_fd_sc_hd__clkbuf_2 wire2399 (.A(net2400),
    .X(net2399));
 sky130_fd_sc_hd__clkbuf_1 wire2400 (.A(net2401),
    .X(net2400));
 sky130_fd_sc_hd__clkbuf_1 wire2401 (.A(net2402),
    .X(net2401));
 sky130_fd_sc_hd__clkbuf_1 wire2402 (.A(net2403),
    .X(net2402));
 sky130_fd_sc_hd__buf_1 wire2403 (.A(_04527_),
    .X(net2403));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2404 (.A(_04224_),
    .X(net2404));
 sky130_fd_sc_hd__buf_1 wire2405 (.A(_04130_),
    .X(net2405));
 sky130_fd_sc_hd__clkbuf_1 wire2406 (.A(net2407),
    .X(net2406));
 sky130_fd_sc_hd__clkbuf_1 max_length2407 (.A(_04009_),
    .X(net2407));
 sky130_fd_sc_hd__buf_1 wire2408 (.A(_03985_),
    .X(net2408));
 sky130_fd_sc_hd__buf_1 wire2409 (.A(net2410),
    .X(net2409));
 sky130_fd_sc_hd__buf_1 wire2410 (.A(_03962_),
    .X(net2410));
 sky130_fd_sc_hd__buf_1 wire2411 (.A(_03786_),
    .X(net2411));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2412 (.A(_03604_),
    .X(net2412));
 sky130_fd_sc_hd__buf_1 wire2413 (.A(_03501_),
    .X(net2413));
 sky130_fd_sc_hd__clkbuf_1 wire2414 (.A(net2415),
    .X(net2414));
 sky130_fd_sc_hd__clkbuf_1 wire2415 (.A(net2416),
    .X(net2415));
 sky130_fd_sc_hd__buf_1 wire2416 (.A(_03480_),
    .X(net2416));
 sky130_fd_sc_hd__clkbuf_1 wire2417 (.A(net2418),
    .X(net2417));
 sky130_fd_sc_hd__clkbuf_1 wire2418 (.A(net2419),
    .X(net2418));
 sky130_fd_sc_hd__buf_1 wire2419 (.A(_03388_),
    .X(net2419));
 sky130_fd_sc_hd__clkbuf_2 wire2420 (.A(net2421),
    .X(net2420));
 sky130_fd_sc_hd__clkbuf_1 wire2421 (.A(net2422),
    .X(net2421));
 sky130_fd_sc_hd__clkbuf_1 wire2422 (.A(net2423),
    .X(net2422));
 sky130_fd_sc_hd__clkbuf_1 wire2423 (.A(_03356_),
    .X(net2423));
 sky130_fd_sc_hd__clkbuf_2 wire2424 (.A(net2425),
    .X(net2424));
 sky130_fd_sc_hd__clkbuf_1 wire2425 (.A(_03343_),
    .X(net2425));
 sky130_fd_sc_hd__buf_1 wire2426 (.A(_03333_),
    .X(net2426));
 sky130_fd_sc_hd__buf_1 wire2427 (.A(_03271_),
    .X(net2427));
 sky130_fd_sc_hd__buf_1 wire2428 (.A(_03225_),
    .X(net2428));
 sky130_fd_sc_hd__buf_1 wire2429 (.A(_03205_),
    .X(net2429));
 sky130_fd_sc_hd__buf_1 wire2430 (.A(_03102_),
    .X(net2430));
 sky130_fd_sc_hd__buf_1 wire2431 (.A(_02995_),
    .X(net2431));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2432 (.A(_02937_),
    .X(net2432));
 sky130_fd_sc_hd__clkbuf_2 wire2433 (.A(_02869_),
    .X(net2433));
 sky130_fd_sc_hd__clkbuf_1 wire2434 (.A(net2435),
    .X(net2434));
 sky130_fd_sc_hd__clkbuf_1 wire2435 (.A(net2436),
    .X(net2435));
 sky130_fd_sc_hd__clkbuf_1 wire2436 (.A(net2437),
    .X(net2436));
 sky130_fd_sc_hd__clkbuf_1 wire2437 (.A(net2438),
    .X(net2437));
 sky130_fd_sc_hd__clkbuf_1 wire2438 (.A(_02660_),
    .X(net2438));
 sky130_fd_sc_hd__buf_1 wire2439 (.A(net2440),
    .X(net2439));
 sky130_fd_sc_hd__buf_1 wire2440 (.A(net2441),
    .X(net2440));
 sky130_fd_sc_hd__clkbuf_1 wire2441 (.A(net2442),
    .X(net2441));
 sky130_fd_sc_hd__clkbuf_1 wire2442 (.A(net2443),
    .X(net2442));
 sky130_fd_sc_hd__clkbuf_1 wire2443 (.A(net2444),
    .X(net2443));
 sky130_fd_sc_hd__clkbuf_1 wire2444 (.A(net2445),
    .X(net2444));
 sky130_fd_sc_hd__buf_1 wire2445 (.A(net2446),
    .X(net2445));
 sky130_fd_sc_hd__buf_1 wire2446 (.A(_02624_),
    .X(net2446));
 sky130_fd_sc_hd__buf_1 max_length2447 (.A(net2448),
    .X(net2447));
 sky130_fd_sc_hd__buf_2 wire2448 (.A(net2449),
    .X(net2448));
 sky130_fd_sc_hd__clkbuf_1 wire2449 (.A(net2450),
    .X(net2449));
 sky130_fd_sc_hd__clkbuf_1 wire2450 (.A(net2454),
    .X(net2450));
 sky130_fd_sc_hd__buf_1 wire2451 (.A(net2452),
    .X(net2451));
 sky130_fd_sc_hd__clkbuf_1 wire2452 (.A(net2453),
    .X(net2452));
 sky130_fd_sc_hd__clkbuf_1 wire2453 (.A(net2454),
    .X(net2453));
 sky130_fd_sc_hd__buf_1 wire2454 (.A(_02620_),
    .X(net2454));
 sky130_fd_sc_hd__clkbuf_1 wire2455 (.A(_02603_),
    .X(net2455));
 sky130_fd_sc_hd__clkbuf_1 wire2456 (.A(_02601_),
    .X(net2456));
 sky130_fd_sc_hd__clkbuf_1 wire2457 (.A(net2458),
    .X(net2457));
 sky130_fd_sc_hd__buf_1 wire2458 (.A(_02556_),
    .X(net2458));
 sky130_fd_sc_hd__buf_1 wire2459 (.A(_02543_),
    .X(net2459));
 sky130_fd_sc_hd__buf_1 wire2460 (.A(net2461),
    .X(net2460));
 sky130_fd_sc_hd__buf_1 max_length2461 (.A(_02523_),
    .X(net2461));
 sky130_fd_sc_hd__clkbuf_1 wire2462 (.A(_02520_),
    .X(net2462));
 sky130_fd_sc_hd__buf_1 max_length2463 (.A(net2465),
    .X(net2463));
 sky130_fd_sc_hd__clkbuf_1 max_length2464 (.A(net2465),
    .X(net2464));
 sky130_fd_sc_hd__buf_1 wire2465 (.A(net2466),
    .X(net2465));
 sky130_fd_sc_hd__buf_1 wire2466 (.A(net2467),
    .X(net2466));
 sky130_fd_sc_hd__buf_1 max_length2467 (.A(net2468),
    .X(net2467));
 sky130_fd_sc_hd__buf_1 wire2468 (.A(net2469),
    .X(net2468));
 sky130_fd_sc_hd__clkbuf_1 wire2469 (.A(_02520_),
    .X(net2469));
 sky130_fd_sc_hd__clkbuf_1 wire2470 (.A(_02362_),
    .X(net2470));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2471 (.A(_02301_),
    .X(net2471));
 sky130_fd_sc_hd__buf_1 wire2472 (.A(_02299_),
    .X(net2472));
 sky130_fd_sc_hd__buf_1 wire2473 (.A(_02225_),
    .X(net2473));
 sky130_fd_sc_hd__buf_1 wire2474 (.A(_01852_),
    .X(net2474));
 sky130_fd_sc_hd__buf_1 wire2475 (.A(_01785_),
    .X(net2475));
 sky130_fd_sc_hd__buf_1 wire2476 (.A(net2477),
    .X(net2476));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2477 (.A(_01710_),
    .X(net2477));
 sky130_fd_sc_hd__clkbuf_1 wire2478 (.A(_01341_),
    .X(net2478));
 sky130_fd_sc_hd__buf_1 wire2479 (.A(_01306_),
    .X(net2479));
 sky130_fd_sc_hd__buf_1 wire2480 (.A(_01052_),
    .X(net2480));
 sky130_fd_sc_hd__buf_1 wire2481 (.A(_00905_),
    .X(net2481));
 sky130_fd_sc_hd__buf_1 wire2482 (.A(_00886_),
    .X(net2482));
 sky130_fd_sc_hd__buf_1 wire2483 (.A(_00846_),
    .X(net2483));
 sky130_fd_sc_hd__buf_1 wire2484 (.A(_00809_),
    .X(net2484));
 sky130_fd_sc_hd__buf_1 wire2485 (.A(_12532_),
    .X(net2485));
 sky130_fd_sc_hd__buf_1 wire2486 (.A(_12525_),
    .X(net2486));
 sky130_fd_sc_hd__buf_1 wire2487 (.A(net2488),
    .X(net2487));
 sky130_fd_sc_hd__buf_1 wire2488 (.A(net2489),
    .X(net2488));
 sky130_fd_sc_hd__buf_1 wire2489 (.A(_12502_),
    .X(net2489));
 sky130_fd_sc_hd__clkbuf_1 wire2490 (.A(_12317_),
    .X(net2490));
 sky130_fd_sc_hd__clkbuf_1 wire2491 (.A(_12299_),
    .X(net2491));
 sky130_fd_sc_hd__buf_1 wire2492 (.A(_12278_),
    .X(net2492));
 sky130_fd_sc_hd__buf_1 wire2493 (.A(_11893_),
    .X(net2493));
 sky130_fd_sc_hd__buf_1 wire2494 (.A(net2495),
    .X(net2494));
 sky130_fd_sc_hd__clkbuf_1 wire2495 (.A(net2496),
    .X(net2495));
 sky130_fd_sc_hd__clkbuf_1 wire2496 (.A(_11865_),
    .X(net2496));
 sky130_fd_sc_hd__clkbuf_1 wire2497 (.A(_11858_),
    .X(net2497));
 sky130_fd_sc_hd__buf_1 wire2498 (.A(net2499),
    .X(net2498));
 sky130_fd_sc_hd__clkbuf_1 wire2499 (.A(_11763_),
    .X(net2499));
 sky130_fd_sc_hd__buf_1 max_length2500 (.A(net2501),
    .X(net2500));
 sky130_fd_sc_hd__buf_1 wire2501 (.A(_11647_),
    .X(net2501));
 sky130_fd_sc_hd__clkbuf_2 wire2502 (.A(net2503),
    .X(net2502));
 sky130_fd_sc_hd__clkbuf_1 wire2503 (.A(_11491_),
    .X(net2503));
 sky130_fd_sc_hd__clkbuf_2 wire2504 (.A(net2505),
    .X(net2504));
 sky130_fd_sc_hd__buf_1 wire2505 (.A(_11446_),
    .X(net2505));
 sky130_fd_sc_hd__clkbuf_2 max_length2506 (.A(_11446_),
    .X(net2506));
 sky130_fd_sc_hd__buf_1 wire2507 (.A(_11270_),
    .X(net2507));
 sky130_fd_sc_hd__clkbuf_1 wire2508 (.A(_11189_),
    .X(net2508));
 sky130_fd_sc_hd__clkbuf_2 wire2509 (.A(net2510),
    .X(net2509));
 sky130_fd_sc_hd__buf_1 wire2510 (.A(_11158_),
    .X(net2510));
 sky130_fd_sc_hd__buf_1 wire2511 (.A(_11149_),
    .X(net2511));
 sky130_fd_sc_hd__buf_1 wire2512 (.A(_11131_),
    .X(net2512));
 sky130_fd_sc_hd__buf_1 wire2513 (.A(net2515),
    .X(net2513));
 sky130_fd_sc_hd__clkbuf_1 wire2514 (.A(net2515),
    .X(net2514));
 sky130_fd_sc_hd__buf_1 wire2515 (.A(_11127_),
    .X(net2515));
 sky130_fd_sc_hd__buf_1 wire2516 (.A(net2517),
    .X(net2516));
 sky130_fd_sc_hd__clkbuf_1 wire2517 (.A(net2518),
    .X(net2517));
 sky130_fd_sc_hd__buf_1 wire2518 (.A(_11127_),
    .X(net2518));
 sky130_fd_sc_hd__buf_1 wire2519 (.A(_11053_),
    .X(net2519));
 sky130_fd_sc_hd__buf_1 wire2520 (.A(_10992_),
    .X(net2520));
 sky130_fd_sc_hd__buf_1 wire2521 (.A(_10980_),
    .X(net2521));
 sky130_fd_sc_hd__buf_1 wire2522 (.A(_10978_),
    .X(net2522));
 sky130_fd_sc_hd__clkbuf_2 wire2523 (.A(net2524),
    .X(net2523));
 sky130_fd_sc_hd__clkbuf_1 wire2524 (.A(net2525),
    .X(net2524));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2525 (.A(_10899_),
    .X(net2525));
 sky130_fd_sc_hd__clkbuf_1 wire2526 (.A(_10894_),
    .X(net2526));
 sky130_fd_sc_hd__buf_1 wire2527 (.A(_10852_),
    .X(net2527));
 sky130_fd_sc_hd__buf_1 wire2528 (.A(_10826_),
    .X(net2528));
 sky130_fd_sc_hd__clkbuf_1 wire2529 (.A(_10816_),
    .X(net2529));
 sky130_fd_sc_hd__clkbuf_2 wire2530 (.A(_10799_),
    .X(net2530));
 sky130_fd_sc_hd__clkbuf_2 wire2531 (.A(net2532),
    .X(net2531));
 sky130_fd_sc_hd__buf_1 wire2532 (.A(net2533),
    .X(net2532));
 sky130_fd_sc_hd__clkbuf_2 wire2533 (.A(net2534),
    .X(net2533));
 sky130_fd_sc_hd__clkbuf_1 wire2534 (.A(net2535),
    .X(net2534));
 sky130_fd_sc_hd__clkbuf_1 wire2535 (.A(net2536),
    .X(net2535));
 sky130_fd_sc_hd__clkbuf_1 wire2536 (.A(_10770_),
    .X(net2536));
 sky130_fd_sc_hd__clkbuf_1 max_length2537 (.A(_10770_),
    .X(net2537));
 sky130_fd_sc_hd__clkbuf_1 wire2538 (.A(_10486_),
    .X(net2538));
 sky130_fd_sc_hd__clkbuf_2 wire2539 (.A(_10435_),
    .X(net2539));
 sky130_fd_sc_hd__buf_1 wire2540 (.A(_10276_),
    .X(net2540));
 sky130_fd_sc_hd__clkbuf_2 wire2541 (.A(net2542),
    .X(net2541));
 sky130_fd_sc_hd__clkbuf_1 wire2542 (.A(_10228_),
    .X(net2542));
 sky130_fd_sc_hd__buf_1 wire2543 (.A(_10177_),
    .X(net2543));
 sky130_fd_sc_hd__buf_1 wire2544 (.A(_10099_),
    .X(net2544));
 sky130_fd_sc_hd__buf_1 wire2545 (.A(_10068_),
    .X(net2545));
 sky130_fd_sc_hd__buf_1 wire2546 (.A(_10067_),
    .X(net2546));
 sky130_fd_sc_hd__buf_1 wire2547 (.A(_10042_),
    .X(net2547));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2548 (.A(_09931_),
    .X(net2548));
 sky130_fd_sc_hd__clkbuf_2 wire2549 (.A(_09869_),
    .X(net2549));
 sky130_fd_sc_hd__clkbuf_2 wire2550 (.A(_09865_),
    .X(net2550));
 sky130_fd_sc_hd__clkbuf_2 wire2551 (.A(_09857_),
    .X(net2551));
 sky130_fd_sc_hd__buf_1 wire2552 (.A(_09794_),
    .X(net2552));
 sky130_fd_sc_hd__buf_1 wire2553 (.A(_09743_),
    .X(net2553));
 sky130_fd_sc_hd__clkbuf_2 max_length2554 (.A(_09720_),
    .X(net2554));
 sky130_fd_sc_hd__clkbuf_2 wire2555 (.A(net2556),
    .X(net2555));
 sky130_fd_sc_hd__buf_1 wire2556 (.A(net2557),
    .X(net2556));
 sky130_fd_sc_hd__clkbuf_2 wire2557 (.A(net2558),
    .X(net2557));
 sky130_fd_sc_hd__buf_1 wire2558 (.A(_09691_),
    .X(net2558));
 sky130_fd_sc_hd__clkbuf_2 wire2559 (.A(net2560),
    .X(net2559));
 sky130_fd_sc_hd__clkbuf_1 wire2560 (.A(_09683_),
    .X(net2560));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2561 (.A(_09677_),
    .X(net2561));
 sky130_fd_sc_hd__buf_1 wire2562 (.A(_09647_),
    .X(net2562));
 sky130_fd_sc_hd__clkbuf_2 wire2563 (.A(_09631_),
    .X(net2563));
 sky130_fd_sc_hd__buf_1 wire2564 (.A(_09601_),
    .X(net2564));
 sky130_fd_sc_hd__clkbuf_1 wire2565 (.A(_09563_),
    .X(net2565));
 sky130_fd_sc_hd__clkbuf_1 wire2566 (.A(_09517_),
    .X(net2566));
 sky130_fd_sc_hd__buf_1 wire2567 (.A(net2570),
    .X(net2567));
 sky130_fd_sc_hd__buf_1 wire2568 (.A(net2569),
    .X(net2568));
 sky130_fd_sc_hd__buf_1 wire2569 (.A(net2570),
    .X(net2569));
 sky130_fd_sc_hd__buf_1 max_length2570 (.A(net2571),
    .X(net2570));
 sky130_fd_sc_hd__buf_1 wire2571 (.A(_09286_),
    .X(net2571));
 sky130_fd_sc_hd__buf_1 wire2572 (.A(net2573),
    .X(net2572));
 sky130_fd_sc_hd__buf_1 max_length2573 (.A(net2574),
    .X(net2573));
 sky130_fd_sc_hd__buf_1 wire2574 (.A(net2575),
    .X(net2574));
 sky130_fd_sc_hd__buf_1 wire2575 (.A(_09278_),
    .X(net2575));
 sky130_fd_sc_hd__buf_1 wire2576 (.A(net2577),
    .X(net2576));
 sky130_fd_sc_hd__buf_1 wire2577 (.A(net2578),
    .X(net2577));
 sky130_fd_sc_hd__buf_1 wire2578 (.A(_09272_),
    .X(net2578));
 sky130_fd_sc_hd__buf_1 wire2579 (.A(_09272_),
    .X(net2579));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2580 (.A(net2581),
    .X(net2580));
 sky130_fd_sc_hd__buf_1 wire2581 (.A(net2582),
    .X(net2581));
 sky130_fd_sc_hd__buf_1 wire2582 (.A(_09170_),
    .X(net2582));
 sky130_fd_sc_hd__buf_1 wire2583 (.A(net2584),
    .X(net2583));
 sky130_fd_sc_hd__clkbuf_1 wire2584 (.A(net2585),
    .X(net2584));
 sky130_fd_sc_hd__clkbuf_1 wire2585 (.A(_09164_),
    .X(net2585));
 sky130_fd_sc_hd__buf_1 max_length2586 (.A(_09164_),
    .X(net2586));
 sky130_fd_sc_hd__buf_1 wire2587 (.A(_09158_),
    .X(net2587));
 sky130_fd_sc_hd__buf_1 wire2588 (.A(net2589),
    .X(net2588));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2589 (.A(_09158_),
    .X(net2589));
 sky130_fd_sc_hd__clkbuf_1 wire2590 (.A(_09069_),
    .X(net2590));
 sky130_fd_sc_hd__clkbuf_1 wire2591 (.A(net2594),
    .X(net2591));
 sky130_fd_sc_hd__buf_1 max_length2592 (.A(net2593),
    .X(net2592));
 sky130_fd_sc_hd__clkbuf_2 max_length2593 (.A(net2594),
    .X(net2593));
 sky130_fd_sc_hd__buf_1 wire2594 (.A(_09069_),
    .X(net2594));
 sky130_fd_sc_hd__buf_1 wire2595 (.A(_09052_),
    .X(net2595));
 sky130_fd_sc_hd__buf_1 wire2596 (.A(net2598),
    .X(net2596));
 sky130_fd_sc_hd__buf_1 wire2597 (.A(net2598),
    .X(net2597));
 sky130_fd_sc_hd__buf_1 wire2598 (.A(_09033_),
    .X(net2598));
 sky130_fd_sc_hd__buf_1 wire2599 (.A(_09004_),
    .X(net2599));
 sky130_fd_sc_hd__buf_1 wire2600 (.A(net2601),
    .X(net2600));
 sky130_fd_sc_hd__buf_1 max_length2601 (.A(net2602),
    .X(net2601));
 sky130_fd_sc_hd__clkbuf_2 max_length2602 (.A(_09004_),
    .X(net2602));
 sky130_fd_sc_hd__clkbuf_1 wire2603 (.A(_08988_),
    .X(net2603));
 sky130_fd_sc_hd__buf_1 wire2604 (.A(_08970_),
    .X(net2604));
 sky130_fd_sc_hd__clkbuf_1 wire2605 (.A(_08950_),
    .X(net2605));
 sky130_fd_sc_hd__buf_1 wire2606 (.A(_08933_),
    .X(net2606));
 sky130_fd_sc_hd__buf_1 wire2607 (.A(net2610),
    .X(net2607));
 sky130_fd_sc_hd__buf_1 wire2608 (.A(net2610),
    .X(net2608));
 sky130_fd_sc_hd__buf_1 wire2609 (.A(_08925_),
    .X(net2609));
 sky130_fd_sc_hd__buf_1 max_length2610 (.A(_08925_),
    .X(net2610));
 sky130_fd_sc_hd__clkbuf_1 wire2611 (.A(_08882_),
    .X(net2611));
 sky130_fd_sc_hd__buf_1 wire2612 (.A(_08849_),
    .X(net2612));
 sky130_fd_sc_hd__buf_1 wire2613 (.A(_08669_),
    .X(net2613));
 sky130_fd_sc_hd__clkbuf_1 wire2614 (.A(net2615),
    .X(net2614));
 sky130_fd_sc_hd__buf_1 wire2615 (.A(_08648_),
    .X(net2615));
 sky130_fd_sc_hd__buf_1 wire2616 (.A(net2617),
    .X(net2616));
 sky130_fd_sc_hd__buf_1 wire2617 (.A(_08636_),
    .X(net2617));
 sky130_fd_sc_hd__buf_1 wire2618 (.A(_08636_),
    .X(net2618));
 sky130_fd_sc_hd__buf_1 wire2619 (.A(net2620),
    .X(net2619));
 sky130_fd_sc_hd__buf_1 max_length2620 (.A(_08636_),
    .X(net2620));
 sky130_fd_sc_hd__clkbuf_2 wire2621 (.A(net2622),
    .X(net2621));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2622 (.A(_08450_),
    .X(net2622));
 sky130_fd_sc_hd__buf_1 wire2623 (.A(_08040_),
    .X(net2623));
 sky130_fd_sc_hd__buf_1 max_length2624 (.A(_08040_),
    .X(net2624));
 sky130_fd_sc_hd__buf_1 wire2625 (.A(net2626),
    .X(net2625));
 sky130_fd_sc_hd__buf_1 max_length2626 (.A(_07936_),
    .X(net2626));
 sky130_fd_sc_hd__buf_1 max_length2627 (.A(_07936_),
    .X(net2627));
 sky130_fd_sc_hd__clkbuf_2 wire2628 (.A(net2629),
    .X(net2628));
 sky130_fd_sc_hd__buf_1 wire2629 (.A(_07933_),
    .X(net2629));
 sky130_fd_sc_hd__buf_1 wire2630 (.A(_07933_),
    .X(net2630));
 sky130_fd_sc_hd__clkbuf_2 wire2631 (.A(net2632),
    .X(net2631));
 sky130_fd_sc_hd__buf_1 wire2632 (.A(net2633),
    .X(net2632));
 sky130_fd_sc_hd__buf_1 wire2633 (.A(_07866_),
    .X(net2633));
 sky130_fd_sc_hd__buf_1 max_length2634 (.A(net2635),
    .X(net2634));
 sky130_fd_sc_hd__buf_1 wire2635 (.A(net2636),
    .X(net2635));
 sky130_fd_sc_hd__buf_1 wire2636 (.A(net2637),
    .X(net2636));
 sky130_fd_sc_hd__buf_1 wire2637 (.A(_07864_),
    .X(net2637));
 sky130_fd_sc_hd__buf_1 wire2638 (.A(net2639),
    .X(net2638));
 sky130_fd_sc_hd__buf_1 wire2639 (.A(_07843_),
    .X(net2639));
 sky130_fd_sc_hd__buf_1 max_length2640 (.A(_07843_),
    .X(net2640));
 sky130_fd_sc_hd__buf_1 wire2641 (.A(net2642),
    .X(net2641));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2642 (.A(net2644),
    .X(net2642));
 sky130_fd_sc_hd__clkbuf_1 max_length2643 (.A(net2644),
    .X(net2643));
 sky130_fd_sc_hd__buf_1 max_length2644 (.A(_07838_),
    .X(net2644));
 sky130_fd_sc_hd__buf_1 wire2645 (.A(net2646),
    .X(net2645));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2646 (.A(net2647),
    .X(net2646));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2647 (.A(_07780_),
    .X(net2647));
 sky130_fd_sc_hd__clkbuf_2 wire2648 (.A(net2649),
    .X(net2648));
 sky130_fd_sc_hd__buf_1 wire2649 (.A(net2650),
    .X(net2649));
 sky130_fd_sc_hd__buf_1 wire2650 (.A(_07763_),
    .X(net2650));
 sky130_fd_sc_hd__clkbuf_2 wire2651 (.A(net2652),
    .X(net2651));
 sky130_fd_sc_hd__buf_1 wire2652 (.A(_07761_),
    .X(net2652));
 sky130_fd_sc_hd__clkbuf_1 wire2653 (.A(_07759_),
    .X(net2653));
 sky130_fd_sc_hd__buf_1 wire2654 (.A(net2655),
    .X(net2654));
 sky130_fd_sc_hd__buf_1 wire2655 (.A(net2657),
    .X(net2655));
 sky130_fd_sc_hd__buf_1 wire2656 (.A(net2657),
    .X(net2656));
 sky130_fd_sc_hd__buf_1 max_length2657 (.A(_07759_),
    .X(net2657));
 sky130_fd_sc_hd__clkbuf_1 wire2658 (.A(_07724_),
    .X(net2658));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2659 (.A(net2660),
    .X(net2659));
 sky130_fd_sc_hd__buf_1 wire2660 (.A(_07724_),
    .X(net2660));
 sky130_fd_sc_hd__buf_1 wire2661 (.A(net2662),
    .X(net2661));
 sky130_fd_sc_hd__clkbuf_2 wire2662 (.A(net2663),
    .X(net2662));
 sky130_fd_sc_hd__clkbuf_1 wire2663 (.A(net2664),
    .X(net2663));
 sky130_fd_sc_hd__buf_1 wire2664 (.A(net2665),
    .X(net2664));
 sky130_fd_sc_hd__buf_1 wire2665 (.A(_07715_),
    .X(net2665));
 sky130_fd_sc_hd__buf_1 wire2666 (.A(net2667),
    .X(net2666));
 sky130_fd_sc_hd__clkbuf_1 wire2667 (.A(net2668),
    .X(net2667));
 sky130_fd_sc_hd__buf_1 wire2668 (.A(net2669),
    .X(net2668));
 sky130_fd_sc_hd__clkbuf_1 wire2669 (.A(_07713_),
    .X(net2669));
 sky130_fd_sc_hd__buf_1 wire2670 (.A(_07694_),
    .X(net2670));
 sky130_fd_sc_hd__buf_1 wire2671 (.A(_07694_),
    .X(net2671));
 sky130_fd_sc_hd__buf_1 wire2672 (.A(net2673),
    .X(net2672));
 sky130_fd_sc_hd__clkbuf_1 wire2673 (.A(net2674),
    .X(net2673));
 sky130_fd_sc_hd__clkbuf_1 wire2674 (.A(net2675),
    .X(net2674));
 sky130_fd_sc_hd__buf_1 wire2675 (.A(_07681_),
    .X(net2675));
 sky130_fd_sc_hd__buf_1 wire2676 (.A(_07670_),
    .X(net2676));
 sky130_fd_sc_hd__buf_1 wire2677 (.A(_07579_),
    .X(net2677));
 sky130_fd_sc_hd__buf_1 wire2678 (.A(_07560_),
    .X(net2678));
 sky130_fd_sc_hd__buf_1 wire2679 (.A(net2680),
    .X(net2679));
 sky130_fd_sc_hd__buf_1 wire2680 (.A(_07560_),
    .X(net2680));
 sky130_fd_sc_hd__buf_1 wire2681 (.A(_07560_),
    .X(net2681));
 sky130_fd_sc_hd__clkbuf_2 wire2682 (.A(net2683),
    .X(net2682));
 sky130_fd_sc_hd__buf_1 wire2683 (.A(net2684),
    .X(net2683));
 sky130_fd_sc_hd__clkbuf_1 wire2684 (.A(net2685),
    .X(net2684));
 sky130_fd_sc_hd__buf_1 wire2685 (.A(net2686),
    .X(net2685));
 sky130_fd_sc_hd__buf_1 wire2686 (.A(_07534_),
    .X(net2686));
 sky130_fd_sc_hd__clkbuf_1 wire2687 (.A(net2688),
    .X(net2687));
 sky130_fd_sc_hd__clkbuf_1 wire2688 (.A(net2689),
    .X(net2688));
 sky130_fd_sc_hd__buf_1 wire2689 (.A(_07508_),
    .X(net2689));
 sky130_fd_sc_hd__clkbuf_1 wire2690 (.A(_07505_),
    .X(net2690));
 sky130_fd_sc_hd__buf_1 wire2691 (.A(net2692),
    .X(net2691));
 sky130_fd_sc_hd__buf_1 max_length2692 (.A(net2693),
    .X(net2692));
 sky130_fd_sc_hd__buf_1 wire2693 (.A(net2694),
    .X(net2693));
 sky130_fd_sc_hd__buf_1 wire2694 (.A(_07505_),
    .X(net2694));
 sky130_fd_sc_hd__buf_1 wire2695 (.A(net2696),
    .X(net2695));
 sky130_fd_sc_hd__buf_1 wire2696 (.A(_07489_),
    .X(net2696));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2697 (.A(net2698),
    .X(net2697));
 sky130_fd_sc_hd__clkbuf_1 max_length2698 (.A(_07489_),
    .X(net2698));
 sky130_fd_sc_hd__buf_1 wire2699 (.A(_07438_),
    .X(net2699));
 sky130_fd_sc_hd__clkbuf_2 wire2700 (.A(net2701),
    .X(net2700));
 sky130_fd_sc_hd__buf_1 wire2701 (.A(net2702),
    .X(net2701));
 sky130_fd_sc_hd__buf_1 wire2702 (.A(_07368_),
    .X(net2702));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2703 (.A(_07354_),
    .X(net2703));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2704 (.A(_07320_),
    .X(net2704));
 sky130_fd_sc_hd__buf_1 wire2705 (.A(net2706),
    .X(net2705));
 sky130_fd_sc_hd__clkbuf_1 wire2706 (.A(_07309_),
    .X(net2706));
 sky130_fd_sc_hd__clkbuf_2 wire2707 (.A(net2708),
    .X(net2707));
 sky130_fd_sc_hd__buf_1 wire2708 (.A(net2709),
    .X(net2708));
 sky130_fd_sc_hd__clkbuf_1 wire2709 (.A(net2710),
    .X(net2709));
 sky130_fd_sc_hd__clkbuf_1 max_length2710 (.A(_07309_),
    .X(net2710));
 sky130_fd_sc_hd__clkbuf_1 wire2711 (.A(net2713),
    .X(net2711));
 sky130_fd_sc_hd__clkbuf_2 max_length2712 (.A(net2714),
    .X(net2712));
 sky130_fd_sc_hd__buf_1 max_length2713 (.A(net2714),
    .X(net2713));
 sky130_fd_sc_hd__buf_1 wire2714 (.A(_07305_),
    .X(net2714));
 sky130_fd_sc_hd__clkbuf_1 wire2715 (.A(_07287_),
    .X(net2715));
 sky130_fd_sc_hd__clkbuf_1 wire2716 (.A(net2718),
    .X(net2716));
 sky130_fd_sc_hd__buf_1 wire2717 (.A(net2718),
    .X(net2717));
 sky130_fd_sc_hd__buf_1 max_length2718 (.A(net2719),
    .X(net2718));
 sky130_fd_sc_hd__buf_1 wire2719 (.A(net2720),
    .X(net2719));
 sky130_fd_sc_hd__buf_1 wire2720 (.A(_07287_),
    .X(net2720));
 sky130_fd_sc_hd__clkbuf_2 wire2721 (.A(net2722),
    .X(net2721));
 sky130_fd_sc_hd__buf_1 wire2722 (.A(net2723),
    .X(net2722));
 sky130_fd_sc_hd__buf_1 wire2723 (.A(net2724),
    .X(net2723));
 sky130_fd_sc_hd__buf_1 wire2724 (.A(net2725),
    .X(net2724));
 sky130_fd_sc_hd__buf_1 wire2725 (.A(_07268_),
    .X(net2725));
 sky130_fd_sc_hd__buf_1 wire2726 (.A(net2729),
    .X(net2726));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2727 (.A(net2728),
    .X(net2727));
 sky130_fd_sc_hd__clkbuf_1 wire2728 (.A(_07241_),
    .X(net2728));
 sky130_fd_sc_hd__buf_1 max_length2729 (.A(_07241_),
    .X(net2729));
 sky130_fd_sc_hd__buf_1 wire2730 (.A(_07240_),
    .X(net2730));
 sky130_fd_sc_hd__clkbuf_1 max_length2731 (.A(net2733),
    .X(net2731));
 sky130_fd_sc_hd__buf_1 max_length2732 (.A(net2733),
    .X(net2732));
 sky130_fd_sc_hd__buf_1 wire2733 (.A(net2734),
    .X(net2733));
 sky130_fd_sc_hd__buf_1 wire2734 (.A(net2735),
    .X(net2734));
 sky130_fd_sc_hd__buf_1 wire2735 (.A(net2736),
    .X(net2735));
 sky130_fd_sc_hd__clkbuf_1 wire2736 (.A(_07240_),
    .X(net2736));
 sky130_fd_sc_hd__clkbuf_1 wire2737 (.A(net2738),
    .X(net2737));
 sky130_fd_sc_hd__clkbuf_1 wire2738 (.A(net2739),
    .X(net2738));
 sky130_fd_sc_hd__clkbuf_1 wire2739 (.A(_07226_),
    .X(net2739));
 sky130_fd_sc_hd__buf_1 wire2740 (.A(net2741),
    .X(net2740));
 sky130_fd_sc_hd__clkbuf_1 wire2741 (.A(net2742),
    .X(net2741));
 sky130_fd_sc_hd__buf_1 wire2742 (.A(_07226_),
    .X(net2742));
 sky130_fd_sc_hd__clkbuf_1 wire2743 (.A(_07207_),
    .X(net2743));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2744 (.A(net2745),
    .X(net2744));
 sky130_fd_sc_hd__clkbuf_1 wire2745 (.A(net2746),
    .X(net2745));
 sky130_fd_sc_hd__buf_1 wire2746 (.A(net2747),
    .X(net2746));
 sky130_fd_sc_hd__buf_1 wire2747 (.A(net2748),
    .X(net2747));
 sky130_fd_sc_hd__buf_1 wire2748 (.A(_07207_),
    .X(net2748));
 sky130_fd_sc_hd__clkbuf_1 wire2749 (.A(_07205_),
    .X(net2749));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2750 (.A(net2751),
    .X(net2750));
 sky130_fd_sc_hd__buf_1 wire2751 (.A(net2752),
    .X(net2751));
 sky130_fd_sc_hd__buf_1 wire2752 (.A(net2753),
    .X(net2752));
 sky130_fd_sc_hd__buf_1 wire2753 (.A(net2754),
    .X(net2753));
 sky130_fd_sc_hd__clkbuf_1 max_length2754 (.A(_07205_),
    .X(net2754));
 sky130_fd_sc_hd__buf_1 wire2755 (.A(net2756),
    .X(net2755));
 sky130_fd_sc_hd__buf_1 wire2756 (.A(net2757),
    .X(net2756));
 sky130_fd_sc_hd__buf_1 wire2757 (.A(_07204_),
    .X(net2757));
 sky130_fd_sc_hd__buf_1 wire2758 (.A(net2759),
    .X(net2758));
 sky130_fd_sc_hd__buf_1 wire2759 (.A(_07204_),
    .X(net2759));
 sky130_fd_sc_hd__buf_1 wire2760 (.A(_07190_),
    .X(net2760));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2761 (.A(net2762),
    .X(net2761));
 sky130_fd_sc_hd__buf_1 wire2762 (.A(net2763),
    .X(net2762));
 sky130_fd_sc_hd__clkbuf_1 max_length2763 (.A(_07190_),
    .X(net2763));
 sky130_fd_sc_hd__buf_1 wire2764 (.A(net2765),
    .X(net2764));
 sky130_fd_sc_hd__buf_1 wire2765 (.A(net2766),
    .X(net2765));
 sky130_fd_sc_hd__buf_1 wire2766 (.A(net2767),
    .X(net2766));
 sky130_fd_sc_hd__clkbuf_1 wire2767 (.A(net2768),
    .X(net2767));
 sky130_fd_sc_hd__clkbuf_2 wire2768 (.A(net2769),
    .X(net2768));
 sky130_fd_sc_hd__clkbuf_1 wire2769 (.A(net2770),
    .X(net2769));
 sky130_fd_sc_hd__clkbuf_1 wire2770 (.A(net2771),
    .X(net2770));
 sky130_fd_sc_hd__clkbuf_1 wire2771 (.A(_07153_),
    .X(net2771));
 sky130_fd_sc_hd__buf_2 wire2772 (.A(net2773),
    .X(net2772));
 sky130_fd_sc_hd__clkbuf_1 wire2773 (.A(net2774),
    .X(net2773));
 sky130_fd_sc_hd__clkbuf_1 wire2774 (.A(net2775),
    .X(net2774));
 sky130_fd_sc_hd__clkbuf_1 wire2775 (.A(_07146_),
    .X(net2775));
 sky130_fd_sc_hd__buf_1 max_length2776 (.A(net2778),
    .X(net2776));
 sky130_fd_sc_hd__clkbuf_1 max_length2777 (.A(net2778),
    .X(net2777));
 sky130_fd_sc_hd__buf_1 wire2778 (.A(_07142_),
    .X(net2778));
 sky130_fd_sc_hd__buf_1 max_length2779 (.A(_07142_),
    .X(net2779));
 sky130_fd_sc_hd__buf_1 max_length2780 (.A(net2781),
    .X(net2780));
 sky130_fd_sc_hd__buf_1 wire2781 (.A(_07140_),
    .X(net2781));
 sky130_fd_sc_hd__buf_1 wire2782 (.A(_07140_),
    .X(net2782));
 sky130_fd_sc_hd__buf_1 wire2783 (.A(net2784),
    .X(net2783));
 sky130_fd_sc_hd__buf_1 wire2784 (.A(net2785),
    .X(net2784));
 sky130_fd_sc_hd__clkbuf_1 wire2785 (.A(net2786),
    .X(net2785));
 sky130_fd_sc_hd__buf_1 wire2786 (.A(net2787),
    .X(net2786));
 sky130_fd_sc_hd__clkbuf_1 wire2787 (.A(net2788),
    .X(net2787));
 sky130_fd_sc_hd__buf_1 wire2788 (.A(_07138_),
    .X(net2788));
 sky130_fd_sc_hd__buf_1 max_length2789 (.A(_07138_),
    .X(net2789));
 sky130_fd_sc_hd__buf_1 wire2790 (.A(_07134_),
    .X(net2790));
 sky130_fd_sc_hd__clkbuf_2 wire2791 (.A(net2792),
    .X(net2791));
 sky130_fd_sc_hd__clkbuf_1 wire2792 (.A(net2793),
    .X(net2792));
 sky130_fd_sc_hd__clkbuf_1 wire2793 (.A(_07134_),
    .X(net2793));
 sky130_fd_sc_hd__buf_1 wire2794 (.A(net2795),
    .X(net2794));
 sky130_fd_sc_hd__buf_1 max_length2795 (.A(net2796),
    .X(net2795));
 sky130_fd_sc_hd__buf_1 wire2796 (.A(net2797),
    .X(net2796));
 sky130_fd_sc_hd__buf_1 wire2797 (.A(net2798),
    .X(net2797));
 sky130_fd_sc_hd__clkbuf_1 max_length2798 (.A(_07129_),
    .X(net2798));
 sky130_fd_sc_hd__buf_1 wire2799 (.A(net2800),
    .X(net2799));
 sky130_fd_sc_hd__buf_1 wire2800 (.A(net2801),
    .X(net2800));
 sky130_fd_sc_hd__buf_1 wire2801 (.A(_07125_),
    .X(net2801));
 sky130_fd_sc_hd__buf_1 max_length2802 (.A(net2803),
    .X(net2802));
 sky130_fd_sc_hd__buf_1 wire2803 (.A(net2804),
    .X(net2803));
 sky130_fd_sc_hd__buf_1 wire2804 (.A(net2805),
    .X(net2804));
 sky130_fd_sc_hd__buf_1 wire2805 (.A(net2806),
    .X(net2805));
 sky130_fd_sc_hd__buf_1 wire2806 (.A(net2807),
    .X(net2806));
 sky130_fd_sc_hd__buf_1 wire2807 (.A(_07108_),
    .X(net2807));
 sky130_fd_sc_hd__clkbuf_1 max_length2808 (.A(_07108_),
    .X(net2808));
 sky130_fd_sc_hd__clkbuf_1 wire2809 (.A(_07100_),
    .X(net2809));
 sky130_fd_sc_hd__clkbuf_1 max_length2810 (.A(net2812),
    .X(net2810));
 sky130_fd_sc_hd__buf_1 wire2811 (.A(net2813),
    .X(net2811));
 sky130_fd_sc_hd__buf_1 max_length2812 (.A(net2813),
    .X(net2812));
 sky130_fd_sc_hd__buf_1 wire2813 (.A(net2814),
    .X(net2813));
 sky130_fd_sc_hd__buf_1 wire2814 (.A(_07100_),
    .X(net2814));
 sky130_fd_sc_hd__clkbuf_2 wire2815 (.A(net2816),
    .X(net2815));
 sky130_fd_sc_hd__buf_1 wire2816 (.A(net2817),
    .X(net2816));
 sky130_fd_sc_hd__clkbuf_1 wire2817 (.A(net2818),
    .X(net2817));
 sky130_fd_sc_hd__clkbuf_1 wire2818 (.A(net2819),
    .X(net2818));
 sky130_fd_sc_hd__buf_1 wire2819 (.A(net2820),
    .X(net2819));
 sky130_fd_sc_hd__buf_1 max_length2820 (.A(_07092_),
    .X(net2820));
 sky130_fd_sc_hd__clkbuf_1 wire2821 (.A(net2822),
    .X(net2821));
 sky130_fd_sc_hd__buf_1 wire2822 (.A(net2823),
    .X(net2822));
 sky130_fd_sc_hd__clkbuf_1 wire2823 (.A(net2826),
    .X(net2823));
 sky130_fd_sc_hd__buf_1 wire2824 (.A(net2825),
    .X(net2824));
 sky130_fd_sc_hd__clkbuf_1 wire2825 (.A(_07087_),
    .X(net2825));
 sky130_fd_sc_hd__buf_1 max_length2826 (.A(_07087_),
    .X(net2826));
 sky130_fd_sc_hd__buf_1 max_length2827 (.A(net2828),
    .X(net2827));
 sky130_fd_sc_hd__buf_1 wire2828 (.A(_07080_),
    .X(net2828));
 sky130_fd_sc_hd__buf_1 wire2829 (.A(net2830),
    .X(net2829));
 sky130_fd_sc_hd__buf_1 wire2830 (.A(_07080_),
    .X(net2830));
 sky130_fd_sc_hd__clkbuf_1 wire2831 (.A(net2832),
    .X(net2831));
 sky130_fd_sc_hd__buf_1 wire2832 (.A(_07077_),
    .X(net2832));
 sky130_fd_sc_hd__buf_1 wire2833 (.A(_07077_),
    .X(net2833));
 sky130_fd_sc_hd__buf_1 wire2834 (.A(net2835),
    .X(net2834));
 sky130_fd_sc_hd__clkbuf_1 wire2835 (.A(_07041_),
    .X(net2835));
 sky130_fd_sc_hd__buf_1 wire2836 (.A(net2837),
    .X(net2836));
 sky130_fd_sc_hd__buf_1 wire2837 (.A(net2838),
    .X(net2837));
 sky130_fd_sc_hd__buf_1 wire2838 (.A(_07041_),
    .X(net2838));
 sky130_fd_sc_hd__buf_1 wire2839 (.A(_07040_),
    .X(net2839));
 sky130_fd_sc_hd__buf_1 wire2840 (.A(net2841),
    .X(net2840));
 sky130_fd_sc_hd__buf_1 wire2841 (.A(net2842),
    .X(net2841));
 sky130_fd_sc_hd__buf_1 wire2842 (.A(net2843),
    .X(net2842));
 sky130_fd_sc_hd__clkbuf_1 wire2843 (.A(net2844),
    .X(net2843));
 sky130_fd_sc_hd__clkbuf_1 wire2844 (.A(net2845),
    .X(net2844));
 sky130_fd_sc_hd__clkbuf_1 max_length2845 (.A(_07016_),
    .X(net2845));
 sky130_fd_sc_hd__clkbuf_2 wire2846 (.A(net2847),
    .X(net2846));
 sky130_fd_sc_hd__clkbuf_1 wire2847 (.A(net2848),
    .X(net2847));
 sky130_fd_sc_hd__buf_1 wire2848 (.A(_07012_),
    .X(net2848));
 sky130_fd_sc_hd__buf_1 max_length2849 (.A(_07012_),
    .X(net2849));
 sky130_fd_sc_hd__buf_1 wire2850 (.A(_06988_),
    .X(net2850));
 sky130_fd_sc_hd__buf_1 wire2851 (.A(net2852),
    .X(net2851));
 sky130_fd_sc_hd__buf_1 max_length2852 (.A(_06988_),
    .X(net2852));
 sky130_fd_sc_hd__buf_1 wire2853 (.A(net2854),
    .X(net2853));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2854 (.A(_06914_),
    .X(net2854));
 sky130_fd_sc_hd__buf_1 wire2855 (.A(_06911_),
    .X(net2855));
 sky130_fd_sc_hd__clkbuf_1 max_length2856 (.A(_06869_),
    .X(net2856));
 sky130_fd_sc_hd__buf_1 wire2857 (.A(net2859),
    .X(net2857));
 sky130_fd_sc_hd__buf_1 wire2858 (.A(net2859),
    .X(net2858));
 sky130_fd_sc_hd__buf_1 wire2859 (.A(_06869_),
    .X(net2859));
 sky130_fd_sc_hd__buf_1 max_length2860 (.A(net2861),
    .X(net2860));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2861 (.A(_06838_),
    .X(net2861));
 sky130_fd_sc_hd__buf_1 wire2862 (.A(_06838_),
    .X(net2862));
 sky130_fd_sc_hd__clkbuf_1 wire2863 (.A(_06834_),
    .X(net2863));
 sky130_fd_sc_hd__clkbuf_1 wire2864 (.A(_06829_),
    .X(net2864));
 sky130_fd_sc_hd__clkbuf_2 wire2865 (.A(_06824_),
    .X(net2865));
 sky130_fd_sc_hd__buf_1 max_length2866 (.A(_06824_),
    .X(net2866));
 sky130_fd_sc_hd__buf_1 wire2867 (.A(net2868),
    .X(net2867));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2868 (.A(net2870),
    .X(net2868));
 sky130_fd_sc_hd__buf_1 wire2869 (.A(_06820_),
    .X(net2869));
 sky130_fd_sc_hd__clkbuf_1 max_length2870 (.A(_06820_),
    .X(net2870));
 sky130_fd_sc_hd__buf_1 wire2871 (.A(_06814_),
    .X(net2871));
 sky130_fd_sc_hd__buf_1 wire2872 (.A(_06814_),
    .X(net2872));
 sky130_fd_sc_hd__clkbuf_1 wire2873 (.A(net2875),
    .X(net2873));
 sky130_fd_sc_hd__buf_1 max_length2874 (.A(net2875),
    .X(net2874));
 sky130_fd_sc_hd__buf_1 max_length2875 (.A(_06805_),
    .X(net2875));
 sky130_fd_sc_hd__buf_1 wire2876 (.A(net2877),
    .X(net2876));
 sky130_fd_sc_hd__buf_1 wire2877 (.A(_06802_),
    .X(net2877));
 sky130_fd_sc_hd__buf_1 max_length2878 (.A(_06802_),
    .X(net2878));
 sky130_fd_sc_hd__buf_1 max_length2879 (.A(net2880),
    .X(net2879));
 sky130_fd_sc_hd__buf_1 wire2880 (.A(_06801_),
    .X(net2880));
 sky130_fd_sc_hd__buf_1 wire2881 (.A(_06719_),
    .X(net2881));
 sky130_fd_sc_hd__buf_1 max_length2882 (.A(net2883),
    .X(net2882));
 sky130_fd_sc_hd__buf_1 wire2883 (.A(net2884),
    .X(net2883));
 sky130_fd_sc_hd__clkbuf_1 wire2884 (.A(net2885),
    .X(net2884));
 sky130_fd_sc_hd__buf_1 wire2885 (.A(_06719_),
    .X(net2885));
 sky130_fd_sc_hd__clkbuf_2 max_length2886 (.A(net2887),
    .X(net2886));
 sky130_fd_sc_hd__clkbuf_2 wire2887 (.A(net2888),
    .X(net2887));
 sky130_fd_sc_hd__buf_1 wire2888 (.A(_06653_),
    .X(net2888));
 sky130_fd_sc_hd__buf_1 wire2889 (.A(net2890),
    .X(net2889));
 sky130_fd_sc_hd__buf_1 wire2890 (.A(_06603_),
    .X(net2890));
 sky130_fd_sc_hd__buf_1 wire2891 (.A(net2892),
    .X(net2891));
 sky130_fd_sc_hd__buf_1 max_length2892 (.A(_06603_),
    .X(net2892));
 sky130_fd_sc_hd__buf_1 wire2893 (.A(_06569_),
    .X(net2893));
 sky130_fd_sc_hd__buf_1 max_length2894 (.A(net2895),
    .X(net2894));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2895 (.A(_06569_),
    .X(net2895));
 sky130_fd_sc_hd__clkbuf_2 wire2896 (.A(net2897),
    .X(net2896));
 sky130_fd_sc_hd__clkbuf_1 max_length2897 (.A(net2899),
    .X(net2897));
 sky130_fd_sc_hd__buf_1 max_length2898 (.A(net2899),
    .X(net2898));
 sky130_fd_sc_hd__buf_1 wire2899 (.A(net2900),
    .X(net2899));
 sky130_fd_sc_hd__buf_1 wire2900 (.A(_06525_),
    .X(net2900));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire2901 (.A(_06518_),
    .X(net2901));
 sky130_fd_sc_hd__clkbuf_2 wire2902 (.A(net2903),
    .X(net2902));
 sky130_fd_sc_hd__buf_1 wire2903 (.A(net2904),
    .X(net2903));
 sky130_fd_sc_hd__clkbuf_1 wire2904 (.A(net2905),
    .X(net2904));
 sky130_fd_sc_hd__clkbuf_1 wire2905 (.A(net2906),
    .X(net2905));
 sky130_fd_sc_hd__clkbuf_1 wire2906 (.A(net2907),
    .X(net2906));
 sky130_fd_sc_hd__clkbuf_1 wire2907 (.A(net2908),
    .X(net2907));
 sky130_fd_sc_hd__clkbuf_1 wire2908 (.A(net2909),
    .X(net2908));
 sky130_fd_sc_hd__clkbuf_1 wire2909 (.A(net2910),
    .X(net2909));
 sky130_fd_sc_hd__clkbuf_1 wire2910 (.A(net2911),
    .X(net2910));
 sky130_fd_sc_hd__clkbuf_1 wire2911 (.A(net2912),
    .X(net2911));
 sky130_fd_sc_hd__clkbuf_1 wire2912 (.A(net2913),
    .X(net2912));
 sky130_fd_sc_hd__clkbuf_1 wire2913 (.A(_06516_),
    .X(net2913));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length2914 (.A(_06516_),
    .X(net2914));
 sky130_fd_sc_hd__buf_1 wire2915 (.A(net2916),
    .X(net2915));
 sky130_fd_sc_hd__clkbuf_1 wire2916 (.A(net2917),
    .X(net2916));
 sky130_fd_sc_hd__clkbuf_1 wire2917 (.A(net2918),
    .X(net2917));
 sky130_fd_sc_hd__clkbuf_1 wire2918 (.A(net2919),
    .X(net2918));
 sky130_fd_sc_hd__clkbuf_1 wire2919 (.A(net2920),
    .X(net2919));
 sky130_fd_sc_hd__clkbuf_1 wire2920 (.A(net2921),
    .X(net2920));
 sky130_fd_sc_hd__clkbuf_1 wire2921 (.A(net2930),
    .X(net2921));
 sky130_fd_sc_hd__clkbuf_1 max_length2922 (.A(net2923),
    .X(net2922));
 sky130_fd_sc_hd__buf_1 wire2923 (.A(net2924),
    .X(net2923));
 sky130_fd_sc_hd__clkbuf_1 wire2924 (.A(net2925),
    .X(net2924));
 sky130_fd_sc_hd__clkbuf_1 wire2925 (.A(net2926),
    .X(net2925));
 sky130_fd_sc_hd__clkbuf_1 wire2926 (.A(net2927),
    .X(net2926));
 sky130_fd_sc_hd__clkbuf_1 wire2927 (.A(net2928),
    .X(net2927));
 sky130_fd_sc_hd__clkbuf_1 wire2928 (.A(net2929),
    .X(net2928));
 sky130_fd_sc_hd__clkbuf_1 wire2929 (.A(net2930),
    .X(net2929));
 sky130_fd_sc_hd__buf_1 wire2930 (.A(_06514_),
    .X(net2930));
 sky130_fd_sc_hd__buf_2 wire2931 (.A(_06511_),
    .X(net2931));
 sky130_fd_sc_hd__clkbuf_2 wire2932 (.A(net2933),
    .X(net2932));
 sky130_fd_sc_hd__clkbuf_1 wire2933 (.A(net2934),
    .X(net2933));
 sky130_fd_sc_hd__clkbuf_1 wire2934 (.A(net2935),
    .X(net2934));
 sky130_fd_sc_hd__clkbuf_1 max_length2935 (.A(_06506_),
    .X(net2935));
 sky130_fd_sc_hd__clkbuf_2 wire2936 (.A(net2937),
    .X(net2936));
 sky130_fd_sc_hd__clkbuf_2 wire2937 (.A(net2938),
    .X(net2937));
 sky130_fd_sc_hd__clkbuf_1 wire2938 (.A(net2939),
    .X(net2938));
 sky130_fd_sc_hd__clkbuf_1 wire2939 (.A(net2940),
    .X(net2939));
 sky130_fd_sc_hd__clkbuf_1 wire2940 (.A(net2941),
    .X(net2940));
 sky130_fd_sc_hd__clkbuf_1 wire2941 (.A(_06501_),
    .X(net2941));
 sky130_fd_sc_hd__buf_1 wire2942 (.A(net2943),
    .X(net2942));
 sky130_fd_sc_hd__clkbuf_1 wire2943 (.A(_06501_),
    .X(net2943));
 sky130_fd_sc_hd__buf_1 wire2944 (.A(net2945),
    .X(net2944));
 sky130_fd_sc_hd__clkbuf_1 wire2945 (.A(_05689_),
    .X(net2945));
 sky130_fd_sc_hd__buf_1 wire2946 (.A(net2947),
    .X(net2946));
 sky130_fd_sc_hd__buf_1 wire2947 (.A(net2949),
    .X(net2947));
 sky130_fd_sc_hd__buf_1 wire2948 (.A(net2949),
    .X(net2948));
 sky130_fd_sc_hd__buf_1 wire2949 (.A(_05619_),
    .X(net2949));
 sky130_fd_sc_hd__buf_1 wire2950 (.A(net2951),
    .X(net2950));
 sky130_fd_sc_hd__clkbuf_1 wire2951 (.A(net2952),
    .X(net2951));
 sky130_fd_sc_hd__clkbuf_1 wire2952 (.A(net2953),
    .X(net2952));
 sky130_fd_sc_hd__clkbuf_1 wire2953 (.A(net2954),
    .X(net2953));
 sky130_fd_sc_hd__buf_1 wire2954 (.A(net2955),
    .X(net2954));
 sky130_fd_sc_hd__buf_1 wire2955 (.A(_05346_),
    .X(net2955));
 sky130_fd_sc_hd__clkbuf_1 max_length2956 (.A(_05346_),
    .X(net2956));
 sky130_fd_sc_hd__clkbuf_1 wire2957 (.A(net2958),
    .X(net2957));
 sky130_fd_sc_hd__buf_1 wire2958 (.A(net2960),
    .X(net2958));
 sky130_fd_sc_hd__buf_1 wire2959 (.A(net2960),
    .X(net2959));
 sky130_fd_sc_hd__buf_1 wire2960 (.A(net2961),
    .X(net2960));
 sky130_fd_sc_hd__buf_1 wire2961 (.A(net2962),
    .X(net2961));
 sky130_fd_sc_hd__clkbuf_1 wire2962 (.A(net2963),
    .X(net2962));
 sky130_fd_sc_hd__buf_1 wire2963 (.A(_05285_),
    .X(net2963));
 sky130_fd_sc_hd__buf_1 wire2964 (.A(net2965),
    .X(net2964));
 sky130_fd_sc_hd__buf_1 wire2965 (.A(_05190_),
    .X(net2965));
 sky130_fd_sc_hd__buf_1 wire2966 (.A(_05128_),
    .X(net2966));
 sky130_fd_sc_hd__buf_1 wire2967 (.A(net2968),
    .X(net2967));
 sky130_fd_sc_hd__buf_1 wire2968 (.A(net2969),
    .X(net2968));
 sky130_fd_sc_hd__clkbuf_1 wire2969 (.A(net2970),
    .X(net2969));
 sky130_fd_sc_hd__buf_1 wire2970 (.A(_05054_),
    .X(net2970));
 sky130_fd_sc_hd__buf_1 max_length2971 (.A(net2972),
    .X(net2971));
 sky130_fd_sc_hd__buf_1 wire2972 (.A(_04963_),
    .X(net2972));
 sky130_fd_sc_hd__buf_1 max_length2973 (.A(_04962_),
    .X(net2973));
 sky130_fd_sc_hd__buf_1 max_length2974 (.A(net2975),
    .X(net2974));
 sky130_fd_sc_hd__buf_1 wire2975 (.A(_04958_),
    .X(net2975));
 sky130_fd_sc_hd__clkbuf_1 max_length2976 (.A(_04956_),
    .X(net2976));
 sky130_fd_sc_hd__clkbuf_1 wire2977 (.A(net2978),
    .X(net2977));
 sky130_fd_sc_hd__buf_1 wire2978 (.A(net2979),
    .X(net2978));
 sky130_fd_sc_hd__clkbuf_1 wire2979 (.A(net2980),
    .X(net2979));
 sky130_fd_sc_hd__clkbuf_1 wire2980 (.A(_04929_),
    .X(net2980));
 sky130_fd_sc_hd__buf_1 wire2981 (.A(net2983),
    .X(net2981));
 sky130_fd_sc_hd__buf_1 max_length2982 (.A(net2983),
    .X(net2982));
 sky130_fd_sc_hd__buf_1 wire2983 (.A(net2984),
    .X(net2983));
 sky130_fd_sc_hd__buf_1 wire2984 (.A(net2985),
    .X(net2984));
 sky130_fd_sc_hd__clkbuf_1 wire2985 (.A(net2986),
    .X(net2985));
 sky130_fd_sc_hd__buf_1 wire2986 (.A(net2987),
    .X(net2986));
 sky130_fd_sc_hd__clkbuf_1 wire2987 (.A(_04909_),
    .X(net2987));
 sky130_fd_sc_hd__clkbuf_1 wire2988 (.A(_04909_),
    .X(net2988));
 sky130_fd_sc_hd__buf_1 wire2989 (.A(_04906_),
    .X(net2989));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length2990 (.A(net2991),
    .X(net2990));
 sky130_fd_sc_hd__buf_1 wire2991 (.A(_04890_),
    .X(net2991));
 sky130_fd_sc_hd__buf_1 wire2992 (.A(_04890_),
    .X(net2992));
 sky130_fd_sc_hd__buf_1 wire2993 (.A(net2994),
    .X(net2993));
 sky130_fd_sc_hd__clkbuf_2 wire2994 (.A(net2995),
    .X(net2994));
 sky130_fd_sc_hd__clkbuf_1 wire2995 (.A(net2996),
    .X(net2995));
 sky130_fd_sc_hd__clkbuf_1 wire2996 (.A(net2997),
    .X(net2996));
 sky130_fd_sc_hd__buf_1 wire2997 (.A(net2998),
    .X(net2997));
 sky130_fd_sc_hd__clkbuf_1 wire2998 (.A(net2999),
    .X(net2998));
 sky130_fd_sc_hd__clkbuf_1 wire2999 (.A(_00003_),
    .X(net2999));
 sky130_fd_sc_hd__clkbuf_1 max_length3000 (.A(_00003_),
    .X(net3000));
 sky130_fd_sc_hd__clkbuf_1 wire3001 (.A(net3002),
    .X(net3001));
 sky130_fd_sc_hd__clkbuf_1 wire3002 (.A(_00000_),
    .X(net3002));
 sky130_fd_sc_hd__buf_1 max_length3003 (.A(net3004),
    .X(net3003));
 sky130_fd_sc_hd__buf_1 wire3004 (.A(net3005),
    .X(net3004));
 sky130_fd_sc_hd__buf_1 wire3005 (.A(net3006),
    .X(net3005));
 sky130_fd_sc_hd__buf_1 max_length3006 (.A(_00000_),
    .X(net3006));
 sky130_fd_sc_hd__buf_1 wire3007 (.A(net3008),
    .X(net3007));
 sky130_fd_sc_hd__buf_1 max_length3008 (.A(_00008_),
    .X(net3008));
 sky130_fd_sc_hd__clkbuf_2 max_length3009 (.A(_00008_),
    .X(net3009));
 sky130_fd_sc_hd__buf_1 wire3010 (.A(net3011),
    .X(net3010));
 sky130_fd_sc_hd__clkbuf_1 wire3011 (.A(net3012),
    .X(net3011));
 sky130_fd_sc_hd__clkbuf_1 wire3012 (.A(net3013),
    .X(net3012));
 sky130_fd_sc_hd__clkbuf_1 wire3013 (.A(net3014),
    .X(net3013));
 sky130_fd_sc_hd__clkbuf_1 wire3014 (.A(net3015),
    .X(net3014));
 sky130_fd_sc_hd__clkbuf_1 wire3015 (.A(net3018),
    .X(net3015));
 sky130_fd_sc_hd__buf_1 wire3016 (.A(net3017),
    .X(net3016));
 sky130_fd_sc_hd__buf_1 max_length3017 (.A(net3018),
    .X(net3017));
 sky130_fd_sc_hd__buf_1 wire3018 (.A(_04874_),
    .X(net3018));
 sky130_fd_sc_hd__clkbuf_1 wire3019 (.A(net3020),
    .X(net3019));
 sky130_fd_sc_hd__buf_1 wire3020 (.A(net3021),
    .X(net3020));
 sky130_fd_sc_hd__buf_1 wire3021 (.A(net3027),
    .X(net3021));
 sky130_fd_sc_hd__buf_1 wire3022 (.A(net3023),
    .X(net3022));
 sky130_fd_sc_hd__clkbuf_1 wire3023 (.A(net3024),
    .X(net3023));
 sky130_fd_sc_hd__clkbuf_1 wire3024 (.A(net3025),
    .X(net3024));
 sky130_fd_sc_hd__clkbuf_1 wire3025 (.A(net3026),
    .X(net3025));
 sky130_fd_sc_hd__clkbuf_1 wire3026 (.A(_04870_),
    .X(net3026));
 sky130_fd_sc_hd__clkbuf_1 max_length3027 (.A(_04870_),
    .X(net3027));
 sky130_fd_sc_hd__buf_1 wire3028 (.A(net3029),
    .X(net3028));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3029 (.A(_04857_),
    .X(net3029));
 sky130_fd_sc_hd__buf_1 wire3030 (.A(_04857_),
    .X(net3030));
 sky130_fd_sc_hd__buf_1 wire3031 (.A(net3032),
    .X(net3031));
 sky130_fd_sc_hd__buf_1 wire3032 (.A(_04857_),
    .X(net3032));
 sky130_fd_sc_hd__buf_1 wire3033 (.A(_04849_),
    .X(net3033));
 sky130_fd_sc_hd__clkbuf_1 wire3034 (.A(net3035),
    .X(net3034));
 sky130_fd_sc_hd__clkbuf_1 wire3035 (.A(net3036),
    .X(net3035));
 sky130_fd_sc_hd__clkbuf_1 wire3036 (.A(_04532_),
    .X(net3036));
 sky130_fd_sc_hd__clkbuf_1 wire3037 (.A(net3038),
    .X(net3037));
 sky130_fd_sc_hd__clkbuf_1 wire3038 (.A(net3039),
    .X(net3038));
 sky130_fd_sc_hd__clkbuf_1 wire3039 (.A(_04348_),
    .X(net3039));
 sky130_fd_sc_hd__clkbuf_2 wire3040 (.A(net3041),
    .X(net3040));
 sky130_fd_sc_hd__clkbuf_2 wire3041 (.A(_03971_),
    .X(net3041));
 sky130_fd_sc_hd__clkbuf_1 wire3042 (.A(_03791_),
    .X(net3042));
 sky130_fd_sc_hd__clkbuf_1 wire3043 (.A(net3048),
    .X(net3043));
 sky130_fd_sc_hd__buf_1 wire3044 (.A(net3045),
    .X(net3044));
 sky130_fd_sc_hd__buf_1 wire3045 (.A(net3046),
    .X(net3045));
 sky130_fd_sc_hd__buf_1 wire3046 (.A(net3047),
    .X(net3046));
 sky130_fd_sc_hd__clkbuf_1 max_length3047 (.A(net3048),
    .X(net3047));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3048 (.A(_03739_),
    .X(net3048));
 sky130_fd_sc_hd__buf_1 wire3049 (.A(_03644_),
    .X(net3049));
 sky130_fd_sc_hd__clkbuf_1 wire3050 (.A(net3051),
    .X(net3050));
 sky130_fd_sc_hd__clkbuf_1 wire3051 (.A(_03373_),
    .X(net3051));
 sky130_fd_sc_hd__buf_1 wire3052 (.A(net3053),
    .X(net3052));
 sky130_fd_sc_hd__buf_1 wire3053 (.A(net3054),
    .X(net3053));
 sky130_fd_sc_hd__buf_1 wire3054 (.A(net3055),
    .X(net3054));
 sky130_fd_sc_hd__clkbuf_1 max_length3055 (.A(_03373_),
    .X(net3055));
 sky130_fd_sc_hd__clkbuf_1 wire3056 (.A(net3057),
    .X(net3056));
 sky130_fd_sc_hd__clkbuf_1 wire3057 (.A(net3058),
    .X(net3057));
 sky130_fd_sc_hd__clkbuf_1 wire3058 (.A(_03313_),
    .X(net3058));
 sky130_fd_sc_hd__buf_1 wire3059 (.A(_03198_),
    .X(net3059));
 sky130_fd_sc_hd__buf_1 wire3060 (.A(_03108_),
    .X(net3060));
 sky130_fd_sc_hd__buf_1 wire3061 (.A(net3062),
    .X(net3061));
 sky130_fd_sc_hd__buf_1 wire3062 (.A(net3063),
    .X(net3062));
 sky130_fd_sc_hd__buf_1 wire3063 (.A(_02867_),
    .X(net3063));
 sky130_fd_sc_hd__buf_1 wire3064 (.A(net3067),
    .X(net3064));
 sky130_fd_sc_hd__buf_1 wire3065 (.A(net3066),
    .X(net3065));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3066 (.A(net3067),
    .X(net3066));
 sky130_fd_sc_hd__clkbuf_1 wire3067 (.A(_02722_),
    .X(net3067));
 sky130_fd_sc_hd__buf_1 wire3068 (.A(_02684_),
    .X(net3068));
 sky130_fd_sc_hd__clkbuf_1 wire3069 (.A(_02682_),
    .X(net3069));
 sky130_fd_sc_hd__buf_1 wire3070 (.A(net3071),
    .X(net3070));
 sky130_fd_sc_hd__clkbuf_1 wire3071 (.A(_02680_),
    .X(net3071));
 sky130_fd_sc_hd__buf_1 wire3072 (.A(net3073),
    .X(net3072));
 sky130_fd_sc_hd__clkbuf_1 wire3073 (.A(net3074),
    .X(net3073));
 sky130_fd_sc_hd__clkbuf_1 wire3074 (.A(net3075),
    .X(net3074));
 sky130_fd_sc_hd__clkbuf_1 wire3075 (.A(_02678_),
    .X(net3075));
 sky130_fd_sc_hd__buf_1 wire3076 (.A(net3077),
    .X(net3076));
 sky130_fd_sc_hd__clkbuf_2 wire3077 (.A(net3078),
    .X(net3077));
 sky130_fd_sc_hd__buf_1 wire3078 (.A(_02604_),
    .X(net3078));
 sky130_fd_sc_hd__buf_1 max_length3079 (.A(_02604_),
    .X(net3079));
 sky130_fd_sc_hd__buf_1 wire3080 (.A(net3081),
    .X(net3080));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3081 (.A(_02600_),
    .X(net3081));
 sky130_fd_sc_hd__buf_1 wire3082 (.A(net3086),
    .X(net3082));
 sky130_fd_sc_hd__buf_1 wire3083 (.A(net3084),
    .X(net3083));
 sky130_fd_sc_hd__clkbuf_1 max_length3084 (.A(net3085),
    .X(net3084));
 sky130_fd_sc_hd__buf_1 wire3085 (.A(_02599_),
    .X(net3085));
 sky130_fd_sc_hd__buf_1 max_length3086 (.A(_02599_),
    .X(net3086));
 sky130_fd_sc_hd__buf_1 wire3087 (.A(net3088),
    .X(net3087));
 sky130_fd_sc_hd__buf_1 wire3088 (.A(_02561_),
    .X(net3088));
 sky130_fd_sc_hd__buf_1 wire3089 (.A(_02553_),
    .X(net3089));
 sky130_fd_sc_hd__buf_1 wire3090 (.A(net3091),
    .X(net3090));
 sky130_fd_sc_hd__buf_1 max_length3091 (.A(_02553_),
    .X(net3091));
 sky130_fd_sc_hd__buf_1 wire3092 (.A(_02552_),
    .X(net3092));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3093 (.A(_02546_),
    .X(net3093));
 sky130_fd_sc_hd__clkbuf_2 wire3094 (.A(net3095),
    .X(net3094));
 sky130_fd_sc_hd__buf_1 wire3095 (.A(net3096),
    .X(net3095));
 sky130_fd_sc_hd__clkbuf_1 wire3096 (.A(net3097),
    .X(net3096));
 sky130_fd_sc_hd__clkbuf_1 wire3097 (.A(net3098),
    .X(net3097));
 sky130_fd_sc_hd__buf_1 wire3098 (.A(net3099),
    .X(net3098));
 sky130_fd_sc_hd__clkbuf_1 wire3099 (.A(net3100),
    .X(net3099));
 sky130_fd_sc_hd__clkbuf_1 wire3100 (.A(_02542_),
    .X(net3100));
 sky130_fd_sc_hd__clkbuf_1 wire3101 (.A(net3102),
    .X(net3101));
 sky130_fd_sc_hd__buf_1 wire3102 (.A(net3105),
    .X(net3102));
 sky130_fd_sc_hd__clkbuf_2 wire3103 (.A(net3104),
    .X(net3103));
 sky130_fd_sc_hd__buf_1 wire3104 (.A(_02519_),
    .X(net3104));
 sky130_fd_sc_hd__buf_1 max_length3105 (.A(_02519_),
    .X(net3105));
 sky130_fd_sc_hd__clkbuf_1 wire3106 (.A(net3107),
    .X(net3106));
 sky130_fd_sc_hd__buf_1 wire3107 (.A(net3108),
    .X(net3107));
 sky130_fd_sc_hd__buf_1 wire3108 (.A(net3109),
    .X(net3108));
 sky130_fd_sc_hd__clkbuf_1 wire3109 (.A(net3110),
    .X(net3109));
 sky130_fd_sc_hd__clkbuf_1 wire3110 (.A(_01609_),
    .X(net3110));
 sky130_fd_sc_hd__buf_1 wire3111 (.A(net3112),
    .X(net3111));
 sky130_fd_sc_hd__clkbuf_1 wire3112 (.A(net3113),
    .X(net3112));
 sky130_fd_sc_hd__clkbuf_1 wire3113 (.A(_00961_),
    .X(net3113));
 sky130_fd_sc_hd__clkbuf_1 wire3114 (.A(net3116),
    .X(net3114));
 sky130_fd_sc_hd__clkbuf_1 max_length3115 (.A(net3116),
    .X(net3115));
 sky130_fd_sc_hd__buf_1 wire3116 (.A(net3117),
    .X(net3116));
 sky130_fd_sc_hd__clkbuf_1 wire3117 (.A(net3118),
    .X(net3117));
 sky130_fd_sc_hd__buf_1 wire3118 (.A(net3119),
    .X(net3118));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3119 (.A(net3120),
    .X(net3119));
 sky130_fd_sc_hd__clkbuf_1 wire3120 (.A(_00872_),
    .X(net3120));
 sky130_fd_sc_hd__buf_1 max_length3121 (.A(_00872_),
    .X(net3121));
 sky130_fd_sc_hd__clkbuf_2 wire3122 (.A(net3123),
    .X(net3122));
 sky130_fd_sc_hd__clkbuf_2 wire3123 (.A(_12500_),
    .X(net3123));
 sky130_fd_sc_hd__buf_1 wire3124 (.A(_12313_),
    .X(net3124));
 sky130_fd_sc_hd__clkbuf_2 max_length3125 (.A(_11754_),
    .X(net3125));
 sky130_fd_sc_hd__clkbuf_2 wire3126 (.A(net3127),
    .X(net3126));
 sky130_fd_sc_hd__buf_1 wire3127 (.A(_11620_),
    .X(net3127));
 sky130_fd_sc_hd__clkbuf_1 max_length3128 (.A(net3129),
    .X(net3128));
 sky130_fd_sc_hd__buf_1 wire3129 (.A(_11572_),
    .X(net3129));
 sky130_fd_sc_hd__buf_1 max_length3130 (.A(net3131),
    .X(net3130));
 sky130_fd_sc_hd__buf_1 wire3131 (.A(_11489_),
    .X(net3131));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3132 (.A(net3134),
    .X(net3132));
 sky130_fd_sc_hd__clkbuf_1 max_length3133 (.A(net3134),
    .X(net3133));
 sky130_fd_sc_hd__buf_1 max_length3134 (.A(_11489_),
    .X(net3134));
 sky130_fd_sc_hd__buf_1 wire3135 (.A(net3136),
    .X(net3135));
 sky130_fd_sc_hd__clkbuf_2 wire3136 (.A(_11447_),
    .X(net3136));
 sky130_fd_sc_hd__buf_1 wire3137 (.A(net3138),
    .X(net3137));
 sky130_fd_sc_hd__buf_1 wire3138 (.A(_11431_),
    .X(net3138));
 sky130_fd_sc_hd__clkbuf_1 wire3139 (.A(net3140),
    .X(net3139));
 sky130_fd_sc_hd__buf_1 wire3140 (.A(_11410_),
    .X(net3140));
 sky130_fd_sc_hd__buf_1 wire3141 (.A(net3142),
    .X(net3141));
 sky130_fd_sc_hd__buf_1 wire3142 (.A(_11410_),
    .X(net3142));
 sky130_fd_sc_hd__buf_1 max_length3143 (.A(net3144),
    .X(net3143));
 sky130_fd_sc_hd__buf_1 wire3144 (.A(net3145),
    .X(net3144));
 sky130_fd_sc_hd__buf_1 max_length3145 (.A(net3146),
    .X(net3145));
 sky130_fd_sc_hd__buf_1 wire3146 (.A(_11409_),
    .X(net3146));
 sky130_fd_sc_hd__buf_1 wire3147 (.A(net3148),
    .X(net3147));
 sky130_fd_sc_hd__clkbuf_1 wire3148 (.A(net3149),
    .X(net3148));
 sky130_fd_sc_hd__buf_1 max_length3149 (.A(net3150),
    .X(net3149));
 sky130_fd_sc_hd__buf_1 wire3150 (.A(net3151),
    .X(net3150));
 sky130_fd_sc_hd__buf_1 wire3151 (.A(_11382_),
    .X(net3151));
 sky130_fd_sc_hd__buf_1 wire3152 (.A(net3153),
    .X(net3152));
 sky130_fd_sc_hd__clkbuf_2 wire3153 (.A(net3154),
    .X(net3153));
 sky130_fd_sc_hd__buf_1 wire3154 (.A(_11376_),
    .X(net3154));
 sky130_fd_sc_hd__buf_1 wire3155 (.A(net3156),
    .X(net3155));
 sky130_fd_sc_hd__clkbuf_1 wire3156 (.A(_11349_),
    .X(net3156));
 sky130_fd_sc_hd__clkbuf_2 wire3157 (.A(_11330_),
    .X(net3157));
 sky130_fd_sc_hd__clkbuf_2 wire3158 (.A(net3159),
    .X(net3158));
 sky130_fd_sc_hd__clkbuf_1 wire3159 (.A(net3160),
    .X(net3159));
 sky130_fd_sc_hd__clkbuf_1 wire3160 (.A(_11293_),
    .X(net3160));
 sky130_fd_sc_hd__clkbuf_2 wire3161 (.A(_11273_),
    .X(net3161));
 sky130_fd_sc_hd__clkbuf_2 wire3162 (.A(_11269_),
    .X(net3162));
 sky130_fd_sc_hd__clkbuf_1 wire3163 (.A(net3164),
    .X(net3163));
 sky130_fd_sc_hd__buf_1 wire3164 (.A(net3165),
    .X(net3164));
 sky130_fd_sc_hd__buf_1 wire3165 (.A(net3168),
    .X(net3165));
 sky130_fd_sc_hd__buf_1 wire3166 (.A(net3167),
    .X(net3166));
 sky130_fd_sc_hd__clkbuf_2 wire3167 (.A(_11132_),
    .X(net3167));
 sky130_fd_sc_hd__clkbuf_1 max_length3168 (.A(_11132_),
    .X(net3168));
 sky130_fd_sc_hd__buf_1 wire3169 (.A(net3170),
    .X(net3169));
 sky130_fd_sc_hd__buf_1 wire3170 (.A(net3171),
    .X(net3170));
 sky130_fd_sc_hd__clkbuf_1 wire3171 (.A(net3172),
    .X(net3171));
 sky130_fd_sc_hd__clkbuf_1 wire3172 (.A(net3173),
    .X(net3172));
 sky130_fd_sc_hd__buf_1 wire3173 (.A(_11122_),
    .X(net3173));
 sky130_fd_sc_hd__buf_1 wire3174 (.A(net3175),
    .X(net3174));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3175 (.A(_11061_),
    .X(net3175));
 sky130_fd_sc_hd__buf_1 wire3176 (.A(net3177),
    .X(net3176));
 sky130_fd_sc_hd__buf_1 wire3177 (.A(_11061_),
    .X(net3177));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3178 (.A(net3179),
    .X(net3178));
 sky130_fd_sc_hd__clkbuf_1 wire3179 (.A(_11055_),
    .X(net3179));
 sky130_fd_sc_hd__buf_1 wire3180 (.A(net3181),
    .X(net3180));
 sky130_fd_sc_hd__clkbuf_1 wire3181 (.A(net3182),
    .X(net3181));
 sky130_fd_sc_hd__clkbuf_1 wire3182 (.A(_11037_),
    .X(net3182));
 sky130_fd_sc_hd__buf_1 wire3183 (.A(_11027_),
    .X(net3183));
 sky130_fd_sc_hd__clkbuf_1 wire3184 (.A(_10990_),
    .X(net3184));
 sky130_fd_sc_hd__clkbuf_2 wire3185 (.A(net3186),
    .X(net3185));
 sky130_fd_sc_hd__clkbuf_2 wire3186 (.A(_10973_),
    .X(net3186));
 sky130_fd_sc_hd__clkbuf_2 wire3187 (.A(net3188),
    .X(net3187));
 sky130_fd_sc_hd__clkbuf_1 wire3188 (.A(_10962_),
    .X(net3188));
 sky130_fd_sc_hd__buf_1 wire3189 (.A(_10942_),
    .X(net3189));
 sky130_fd_sc_hd__clkbuf_2 wire3190 (.A(_10938_),
    .X(net3190));
 sky130_fd_sc_hd__buf_1 wire3191 (.A(_10923_),
    .X(net3191));
 sky130_fd_sc_hd__buf_1 wire3192 (.A(_10919_),
    .X(net3192));
 sky130_fd_sc_hd__buf_1 wire3193 (.A(net3194),
    .X(net3193));
 sky130_fd_sc_hd__clkbuf_1 wire3194 (.A(net3195),
    .X(net3194));
 sky130_fd_sc_hd__buf_1 wire3195 (.A(net3197),
    .X(net3195));
 sky130_fd_sc_hd__clkbuf_1 max_length3196 (.A(net3197),
    .X(net3196));
 sky130_fd_sc_hd__buf_1 wire3197 (.A(net3198),
    .X(net3197));
 sky130_fd_sc_hd__buf_1 max_length3198 (.A(_10911_),
    .X(net3198));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3199 (.A(net3200),
    .X(net3199));
 sky130_fd_sc_hd__buf_1 wire3200 (.A(net3201),
    .X(net3200));
 sky130_fd_sc_hd__buf_1 wire3201 (.A(_10871_),
    .X(net3201));
 sky130_fd_sc_hd__buf_1 wire3202 (.A(net3203),
    .X(net3202));
 sky130_fd_sc_hd__buf_1 max_length3203 (.A(_10843_),
    .X(net3203));
 sky130_fd_sc_hd__clkbuf_1 max_length3204 (.A(net3205),
    .X(net3204));
 sky130_fd_sc_hd__buf_1 wire3205 (.A(net3206),
    .X(net3205));
 sky130_fd_sc_hd__buf_1 wire3206 (.A(_10836_),
    .X(net3206));
 sky130_fd_sc_hd__clkbuf_1 wire3207 (.A(net3208),
    .X(net3207));
 sky130_fd_sc_hd__buf_1 wire3208 (.A(_10836_),
    .X(net3208));
 sky130_fd_sc_hd__buf_1 wire3209 (.A(_10829_),
    .X(net3209));
 sky130_fd_sc_hd__buf_1 wire3210 (.A(_10829_),
    .X(net3210));
 sky130_fd_sc_hd__buf_1 wire3211 (.A(net3212),
    .X(net3211));
 sky130_fd_sc_hd__buf_1 wire3212 (.A(_10821_),
    .X(net3212));
 sky130_fd_sc_hd__buf_1 wire3213 (.A(_10811_),
    .X(net3213));
 sky130_fd_sc_hd__clkbuf_2 wire3214 (.A(_10805_),
    .X(net3214));
 sky130_fd_sc_hd__buf_1 wire3215 (.A(_10792_),
    .X(net3215));
 sky130_fd_sc_hd__clkbuf_2 wire3216 (.A(net3217),
    .X(net3216));
 sky130_fd_sc_hd__clkbuf_1 wire3217 (.A(net3218),
    .X(net3217));
 sky130_fd_sc_hd__clkbuf_1 wire3218 (.A(net3219),
    .X(net3218));
 sky130_fd_sc_hd__clkbuf_1 wire3219 (.A(net3220),
    .X(net3219));
 sky130_fd_sc_hd__clkbuf_1 wire3220 (.A(_10789_),
    .X(net3220));
 sky130_fd_sc_hd__buf_1 wire3221 (.A(net3222),
    .X(net3221));
 sky130_fd_sc_hd__buf_1 wire3222 (.A(net3224),
    .X(net3222));
 sky130_fd_sc_hd__buf_1 wire3223 (.A(net3224),
    .X(net3223));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3224 (.A(_10391_),
    .X(net3224));
 sky130_fd_sc_hd__clkbuf_2 max_length3225 (.A(_10223_),
    .X(net3225));
 sky130_fd_sc_hd__clkbuf_1 wire3226 (.A(net3227),
    .X(net3226));
 sky130_fd_sc_hd__clkbuf_1 wire3227 (.A(_10165_),
    .X(net3227));
 sky130_fd_sc_hd__buf_1 wire3228 (.A(_10124_),
    .X(net3228));
 sky130_fd_sc_hd__clkbuf_2 wire3229 (.A(_10104_),
    .X(net3229));
 sky130_fd_sc_hd__clkbuf_1 wire3230 (.A(_10063_),
    .X(net3230));
 sky130_fd_sc_hd__clkbuf_2 wire3231 (.A(net3232),
    .X(net3231));
 sky130_fd_sc_hd__buf_1 max_length3232 (.A(_10063_),
    .X(net3232));
 sky130_fd_sc_hd__buf_1 wire3233 (.A(_10047_),
    .X(net3233));
 sky130_fd_sc_hd__buf_1 wire3234 (.A(_09955_),
    .X(net3234));
 sky130_fd_sc_hd__clkbuf_2 wire3235 (.A(net3236),
    .X(net3235));
 sky130_fd_sc_hd__clkbuf_1 wire3236 (.A(_09880_),
    .X(net3236));
 sky130_fd_sc_hd__buf_1 wire3237 (.A(_09851_),
    .X(net3237));
 sky130_fd_sc_hd__buf_1 wire3238 (.A(_09802_),
    .X(net3238));
 sky130_fd_sc_hd__buf_1 wire3239 (.A(_09801_),
    .X(net3239));
 sky130_fd_sc_hd__buf_1 max_length3240 (.A(net3241),
    .X(net3240));
 sky130_fd_sc_hd__clkbuf_2 wire3241 (.A(_09792_),
    .X(net3241));
 sky130_fd_sc_hd__buf_1 wire3242 (.A(net3243),
    .X(net3242));
 sky130_fd_sc_hd__clkbuf_1 wire3243 (.A(net3244),
    .X(net3243));
 sky130_fd_sc_hd__clkbuf_1 wire3244 (.A(_09737_),
    .X(net3244));
 sky130_fd_sc_hd__clkbuf_2 wire3245 (.A(_09730_),
    .X(net3245));
 sky130_fd_sc_hd__clkbuf_1 wire3246 (.A(net3247),
    .X(net3246));
 sky130_fd_sc_hd__buf_1 wire3247 (.A(_09675_),
    .X(net3247));
 sky130_fd_sc_hd__buf_1 wire3248 (.A(net3249),
    .X(net3248));
 sky130_fd_sc_hd__clkbuf_1 wire3249 (.A(net3250),
    .X(net3249));
 sky130_fd_sc_hd__clkbuf_1 wire3250 (.A(net3251),
    .X(net3250));
 sky130_fd_sc_hd__clkbuf_1 wire3251 (.A(net3252),
    .X(net3251));
 sky130_fd_sc_hd__clkbuf_1 wire3252 (.A(_09662_),
    .X(net3252));
 sky130_fd_sc_hd__buf_1 max_length3253 (.A(net3254),
    .X(net3253));
 sky130_fd_sc_hd__buf_1 wire3254 (.A(_09649_),
    .X(net3254));
 sky130_fd_sc_hd__buf_1 wire3255 (.A(net3256),
    .X(net3255));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3256 (.A(_09649_),
    .X(net3256));
 sky130_fd_sc_hd__buf_1 wire3257 (.A(_09643_),
    .X(net3257));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3258 (.A(_09643_),
    .X(net3258));
 sky130_fd_sc_hd__buf_1 wire3259 (.A(_09638_),
    .X(net3259));
 sky130_fd_sc_hd__clkbuf_2 wire3260 (.A(_09633_),
    .X(net3260));
 sky130_fd_sc_hd__buf_1 max_length3261 (.A(net3262),
    .X(net3261));
 sky130_fd_sc_hd__buf_1 max_length3262 (.A(net3263),
    .X(net3262));
 sky130_fd_sc_hd__clkbuf_2 max_length3263 (.A(_09620_),
    .X(net3263));
 sky130_fd_sc_hd__buf_1 wire3264 (.A(_09615_),
    .X(net3264));
 sky130_fd_sc_hd__clkbuf_2 wire3265 (.A(net3266),
    .X(net3265));
 sky130_fd_sc_hd__buf_1 max_length3266 (.A(_09615_),
    .X(net3266));
 sky130_fd_sc_hd__buf_1 wire3267 (.A(net3268),
    .X(net3267));
 sky130_fd_sc_hd__clkbuf_2 wire3268 (.A(_09600_),
    .X(net3268));
 sky130_fd_sc_hd__buf_1 wire3269 (.A(_09575_),
    .X(net3269));
 sky130_fd_sc_hd__buf_1 wire3270 (.A(_09575_),
    .X(net3270));
 sky130_fd_sc_hd__buf_1 wire3271 (.A(net3272),
    .X(net3271));
 sky130_fd_sc_hd__buf_1 wire3272 (.A(_09393_),
    .X(net3272));
 sky130_fd_sc_hd__buf_1 wire3273 (.A(net3274),
    .X(net3273));
 sky130_fd_sc_hd__buf_1 wire3274 (.A(_09332_),
    .X(net3274));
 sky130_fd_sc_hd__buf_1 wire3275 (.A(_09332_),
    .X(net3275));
 sky130_fd_sc_hd__buf_1 wire3276 (.A(net3277),
    .X(net3276));
 sky130_fd_sc_hd__clkbuf_1 max_length3277 (.A(_09268_),
    .X(net3277));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3278 (.A(net3279),
    .X(net3278));
 sky130_fd_sc_hd__buf_1 wire3279 (.A(_09258_),
    .X(net3279));
 sky130_fd_sc_hd__buf_1 wire3280 (.A(net3281),
    .X(net3280));
 sky130_fd_sc_hd__buf_1 wire3281 (.A(net3283),
    .X(net3281));
 sky130_fd_sc_hd__clkbuf_2 max_length3282 (.A(net3283),
    .X(net3282));
 sky130_fd_sc_hd__buf_1 wire3283 (.A(_09177_),
    .X(net3283));
 sky130_fd_sc_hd__clkbuf_2 max_length3284 (.A(net3285),
    .X(net3284));
 sky130_fd_sc_hd__buf_1 max_length3285 (.A(net3286),
    .X(net3285));
 sky130_fd_sc_hd__buf_1 max_length3286 (.A(net3287),
    .X(net3286));
 sky130_fd_sc_hd__buf_1 wire3287 (.A(net3288),
    .X(net3287));
 sky130_fd_sc_hd__clkbuf_1 wire3288 (.A(net3289),
    .X(net3288));
 sky130_fd_sc_hd__clkbuf_1 max_length3289 (.A(_09157_),
    .X(net3289));
 sky130_fd_sc_hd__buf_1 wire3290 (.A(net3295),
    .X(net3290));
 sky130_fd_sc_hd__buf_1 wire3291 (.A(net3292),
    .X(net3291));
 sky130_fd_sc_hd__buf_1 wire3292 (.A(net3293),
    .X(net3292));
 sky130_fd_sc_hd__clkbuf_1 wire3293 (.A(net3294),
    .X(net3293));
 sky130_fd_sc_hd__buf_1 wire3294 (.A(net3295),
    .X(net3294));
 sky130_fd_sc_hd__buf_1 max_length3295 (.A(_09097_),
    .X(net3295));
 sky130_fd_sc_hd__buf_1 wire3296 (.A(net3297),
    .X(net3296));
 sky130_fd_sc_hd__buf_1 wire3297 (.A(net3299),
    .X(net3297));
 sky130_fd_sc_hd__buf_1 wire3298 (.A(net3299),
    .X(net3298));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3299 (.A(net3300),
    .X(net3299));
 sky130_fd_sc_hd__clkbuf_1 wire3300 (.A(net3301),
    .X(net3300));
 sky130_fd_sc_hd__buf_1 wire3301 (.A(net3302),
    .X(net3301));
 sky130_fd_sc_hd__clkbuf_1 wire3302 (.A(net3303),
    .X(net3302));
 sky130_fd_sc_hd__clkbuf_1 wire3303 (.A(net3304),
    .X(net3303));
 sky130_fd_sc_hd__clkbuf_1 wire3304 (.A(_09093_),
    .X(net3304));
 sky130_fd_sc_hd__buf_2 wire3305 (.A(_09082_),
    .X(net3305));
 sky130_fd_sc_hd__clkbuf_1 wire3306 (.A(net3312),
    .X(net3306));
 sky130_fd_sc_hd__buf_1 wire3307 (.A(net3309),
    .X(net3307));
 sky130_fd_sc_hd__buf_1 max_length3308 (.A(net3309),
    .X(net3308));
 sky130_fd_sc_hd__buf_1 max_length3309 (.A(net3310),
    .X(net3309));
 sky130_fd_sc_hd__buf_1 wire3310 (.A(net3311),
    .X(net3310));
 sky130_fd_sc_hd__buf_1 max_length3311 (.A(net3312),
    .X(net3311));
 sky130_fd_sc_hd__buf_1 wire3312 (.A(_09051_),
    .X(net3312));
 sky130_fd_sc_hd__clkbuf_2 wire3313 (.A(net3314),
    .X(net3313));
 sky130_fd_sc_hd__clkbuf_2 wire3314 (.A(_09031_),
    .X(net3314));
 sky130_fd_sc_hd__clkbuf_1 wire3315 (.A(net3316),
    .X(net3315));
 sky130_fd_sc_hd__buf_1 wire3316 (.A(net3317),
    .X(net3316));
 sky130_fd_sc_hd__buf_1 wire3317 (.A(net3318),
    .X(net3317));
 sky130_fd_sc_hd__clkbuf_1 wire3318 (.A(net3319),
    .X(net3318));
 sky130_fd_sc_hd__clkbuf_1 wire3319 (.A(_09023_),
    .X(net3319));
 sky130_fd_sc_hd__clkbuf_1 wire3320 (.A(net3321),
    .X(net3320));
 sky130_fd_sc_hd__clkbuf_1 wire3321 (.A(net3322),
    .X(net3321));
 sky130_fd_sc_hd__buf_1 wire3322 (.A(net3323),
    .X(net3322));
 sky130_fd_sc_hd__buf_1 wire3323 (.A(net3324),
    .X(net3323));
 sky130_fd_sc_hd__buf_1 wire3324 (.A(_09023_),
    .X(net3324));
 sky130_fd_sc_hd__clkbuf_2 wire3325 (.A(net3326),
    .X(net3325));
 sky130_fd_sc_hd__buf_1 max_length3326 (.A(net3327),
    .X(net3326));
 sky130_fd_sc_hd__buf_1 wire3327 (.A(_09006_),
    .X(net3327));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3328 (.A(net3329),
    .X(net3328));
 sky130_fd_sc_hd__clkbuf_1 wire3329 (.A(net3330),
    .X(net3329));
 sky130_fd_sc_hd__buf_1 max_length3330 (.A(net3331),
    .X(net3330));
 sky130_fd_sc_hd__buf_1 wire3331 (.A(_08985_),
    .X(net3331));
 sky130_fd_sc_hd__buf_1 wire3332 (.A(_08971_),
    .X(net3332));
 sky130_fd_sc_hd__buf_1 max_length3333 (.A(_08971_),
    .X(net3333));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3334 (.A(net3335),
    .X(net3334));
 sky130_fd_sc_hd__clkbuf_2 wire3335 (.A(_08969_),
    .X(net3335));
 sky130_fd_sc_hd__buf_1 wire3336 (.A(net3337),
    .X(net3336));
 sky130_fd_sc_hd__buf_1 wire3337 (.A(net3338),
    .X(net3337));
 sky130_fd_sc_hd__clkbuf_1 wire3338 (.A(net3339),
    .X(net3338));
 sky130_fd_sc_hd__buf_1 wire3339 (.A(net3340),
    .X(net3339));
 sky130_fd_sc_hd__buf_1 max_length3340 (.A(_08967_),
    .X(net3340));
 sky130_fd_sc_hd__clkbuf_1 max_length3341 (.A(net3342),
    .X(net3341));
 sky130_fd_sc_hd__buf_1 wire3342 (.A(_08948_),
    .X(net3342));
 sky130_fd_sc_hd__buf_1 max_length3343 (.A(_08946_),
    .X(net3343));
 sky130_fd_sc_hd__clkbuf_1 wire3344 (.A(_08927_),
    .X(net3344));
 sky130_fd_sc_hd__clkbuf_2 max_length3345 (.A(_08924_),
    .X(net3345));
 sky130_fd_sc_hd__buf_1 wire3346 (.A(net3348),
    .X(net3346));
 sky130_fd_sc_hd__buf_1 wire3347 (.A(net3348),
    .X(net3347));
 sky130_fd_sc_hd__buf_1 wire3348 (.A(_08914_),
    .X(net3348));
 sky130_fd_sc_hd__buf_1 wire3349 (.A(_08914_),
    .X(net3349));
 sky130_fd_sc_hd__clkbuf_1 wire3350 (.A(net3351),
    .X(net3350));
 sky130_fd_sc_hd__buf_1 wire3351 (.A(net3352),
    .X(net3351));
 sky130_fd_sc_hd__clkbuf_1 wire3352 (.A(net3353),
    .X(net3352));
 sky130_fd_sc_hd__buf_1 wire3353 (.A(net3354),
    .X(net3353));
 sky130_fd_sc_hd__buf_1 max_length3354 (.A(net3355),
    .X(net3354));
 sky130_fd_sc_hd__buf_1 wire3355 (.A(net3356),
    .X(net3355));
 sky130_fd_sc_hd__clkbuf_1 wire3356 (.A(_08909_),
    .X(net3356));
 sky130_fd_sc_hd__clkbuf_1 wire3357 (.A(net3358),
    .X(net3357));
 sky130_fd_sc_hd__clkbuf_1 wire3358 (.A(net3359),
    .X(net3358));
 sky130_fd_sc_hd__buf_1 wire3359 (.A(_08909_),
    .X(net3359));
 sky130_fd_sc_hd__clkbuf_1 max_cap3360 (.A(net9246),
    .X(net3360));
 sky130_fd_sc_hd__clkbuf_1 wire3361 (.A(net3362),
    .X(net3361));
 sky130_fd_sc_hd__buf_1 wire3362 (.A(_08843_),
    .X(net3362));
 sky130_fd_sc_hd__buf_1 wire3363 (.A(_08829_),
    .X(net3363));
 sky130_fd_sc_hd__clkbuf_1 wire3364 (.A(_08826_),
    .X(net3364));
 sky130_fd_sc_hd__clkbuf_2 max_length3365 (.A(net3366),
    .X(net3365));
 sky130_fd_sc_hd__clkbuf_2 max_length3366 (.A(_08803_),
    .X(net3366));
 sky130_fd_sc_hd__clkbuf_2 wire3367 (.A(_08792_),
    .X(net3367));
 sky130_fd_sc_hd__clkbuf_2 wire3368 (.A(_08792_),
    .X(net3368));
 sky130_fd_sc_hd__buf_1 wire3369 (.A(net3370),
    .X(net3369));
 sky130_fd_sc_hd__clkbuf_2 wire3370 (.A(net3371),
    .X(net3370));
 sky130_fd_sc_hd__clkbuf_1 wire3371 (.A(net3377),
    .X(net3371));
 sky130_fd_sc_hd__buf_1 max_length3372 (.A(net3373),
    .X(net3372));
 sky130_fd_sc_hd__clkbuf_2 wire3373 (.A(net3374),
    .X(net3373));
 sky130_fd_sc_hd__clkbuf_1 wire3374 (.A(net3375),
    .X(net3374));
 sky130_fd_sc_hd__clkbuf_1 wire3375 (.A(net3376),
    .X(net3375));
 sky130_fd_sc_hd__clkbuf_1 wire3376 (.A(_08781_),
    .X(net3376));
 sky130_fd_sc_hd__clkbuf_1 max_length3377 (.A(_08781_),
    .X(net3377));
 sky130_fd_sc_hd__clkbuf_2 wire3378 (.A(_08770_),
    .X(net3378));
 sky130_fd_sc_hd__buf_1 wire3379 (.A(_08770_),
    .X(net3379));
 sky130_fd_sc_hd__clkbuf_2 wire3380 (.A(net3381),
    .X(net3380));
 sky130_fd_sc_hd__clkbuf_2 wire3381 (.A(net3382),
    .X(net3381));
 sky130_fd_sc_hd__buf_1 wire3382 (.A(_08759_),
    .X(net3382));
 sky130_fd_sc_hd__buf_1 wire3383 (.A(_08663_),
    .X(net3383));
 sky130_fd_sc_hd__buf_1 wire3384 (.A(net3385),
    .X(net3384));
 sky130_fd_sc_hd__clkbuf_1 wire3385 (.A(net3386),
    .X(net3385));
 sky130_fd_sc_hd__buf_1 wire3386 (.A(_08647_),
    .X(net3386));
 sky130_fd_sc_hd__buf_1 max_length3387 (.A(net3388),
    .X(net3387));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3388 (.A(_08647_),
    .X(net3388));
 sky130_fd_sc_hd__buf_1 wire3389 (.A(_08645_),
    .X(net3389));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3390 (.A(net3391),
    .X(net3390));
 sky130_fd_sc_hd__clkbuf_1 wire3391 (.A(_07847_),
    .X(net3391));
 sky130_fd_sc_hd__buf_1 wire3392 (.A(net3393),
    .X(net3392));
 sky130_fd_sc_hd__buf_1 wire3393 (.A(_07723_),
    .X(net3393));
 sky130_fd_sc_hd__buf_1 wire3394 (.A(_07688_),
    .X(net3394));
 sky130_fd_sc_hd__buf_1 max_length3395 (.A(_07688_),
    .X(net3395));
 sky130_fd_sc_hd__buf_1 wire3396 (.A(_07686_),
    .X(net3396));
 sky130_fd_sc_hd__buf_1 wire3397 (.A(_07684_),
    .X(net3397));
 sky130_fd_sc_hd__clkbuf_2 wire3398 (.A(_07654_),
    .X(net3398));
 sky130_fd_sc_hd__buf_1 wire3399 (.A(net3400),
    .X(net3399));
 sky130_fd_sc_hd__buf_1 wire3400 (.A(_07603_),
    .X(net3400));
 sky130_fd_sc_hd__clkbuf_1 wire3401 (.A(net3402),
    .X(net3401));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3402 (.A(net3403),
    .X(net3402));
 sky130_fd_sc_hd__clkbuf_1 wire3403 (.A(_07598_),
    .X(net3403));
 sky130_fd_sc_hd__buf_1 wire3404 (.A(net3406),
    .X(net3404));
 sky130_fd_sc_hd__clkbuf_1 max_length3405 (.A(net3406),
    .X(net3405));
 sky130_fd_sc_hd__buf_1 wire3406 (.A(_07574_),
    .X(net3406));
 sky130_fd_sc_hd__buf_1 wire3407 (.A(net3408),
    .X(net3407));
 sky130_fd_sc_hd__clkbuf_1 wire3408 (.A(_07571_),
    .X(net3408));
 sky130_fd_sc_hd__buf_1 wire3409 (.A(net3410),
    .X(net3409));
 sky130_fd_sc_hd__clkbuf_1 wire3410 (.A(net3411),
    .X(net3410));
 sky130_fd_sc_hd__buf_1 wire3411 (.A(net3412),
    .X(net3411));
 sky130_fd_sc_hd__buf_1 wire3412 (.A(_07528_),
    .X(net3412));
 sky130_fd_sc_hd__buf_1 wire3413 (.A(net3414),
    .X(net3413));
 sky130_fd_sc_hd__buf_1 wire3414 (.A(net3419),
    .X(net3414));
 sky130_fd_sc_hd__buf_1 max_length3415 (.A(net3416),
    .X(net3415));
 sky130_fd_sc_hd__buf_1 wire3416 (.A(net3417),
    .X(net3416));
 sky130_fd_sc_hd__buf_1 wire3417 (.A(net3418),
    .X(net3417));
 sky130_fd_sc_hd__buf_1 wire3418 (.A(net3419),
    .X(net3418));
 sky130_fd_sc_hd__buf_1 wire3419 (.A(_07516_),
    .X(net3419));
 sky130_fd_sc_hd__buf_1 wire3420 (.A(net3421),
    .X(net3420));
 sky130_fd_sc_hd__buf_1 wire3421 (.A(net3422),
    .X(net3421));
 sky130_fd_sc_hd__buf_1 wire3422 (.A(_07511_),
    .X(net3422));
 sky130_fd_sc_hd__buf_1 wire3423 (.A(_07507_),
    .X(net3423));
 sky130_fd_sc_hd__buf_1 wire3424 (.A(_07486_),
    .X(net3424));
 sky130_fd_sc_hd__buf_1 wire3425 (.A(net3426),
    .X(net3425));
 sky130_fd_sc_hd__buf_1 wire3426 (.A(_07486_),
    .X(net3426));
 sky130_fd_sc_hd__buf_1 wire3427 (.A(net3428),
    .X(net3427));
 sky130_fd_sc_hd__buf_1 wire3428 (.A(net3430),
    .X(net3428));
 sky130_fd_sc_hd__buf_1 wire3429 (.A(net3430),
    .X(net3429));
 sky130_fd_sc_hd__buf_1 wire3430 (.A(_07485_),
    .X(net3430));
 sky130_fd_sc_hd__buf_1 wire3431 (.A(net3432),
    .X(net3431));
 sky130_fd_sc_hd__buf_1 wire3432 (.A(net3433),
    .X(net3432));
 sky130_fd_sc_hd__clkbuf_1 wire3433 (.A(_07378_),
    .X(net3433));
 sky130_fd_sc_hd__buf_1 wire3434 (.A(net3437),
    .X(net3434));
 sky130_fd_sc_hd__buf_1 wire3435 (.A(net3436),
    .X(net3435));
 sky130_fd_sc_hd__buf_1 wire3436 (.A(net3437),
    .X(net3436));
 sky130_fd_sc_hd__buf_1 wire3437 (.A(net3438),
    .X(net3437));
 sky130_fd_sc_hd__buf_1 wire3438 (.A(_07371_),
    .X(net3438));
 sky130_fd_sc_hd__buf_1 max_length3439 (.A(net3440),
    .X(net3439));
 sky130_fd_sc_hd__buf_1 wire3440 (.A(net3441),
    .X(net3440));
 sky130_fd_sc_hd__buf_1 wire3441 (.A(_07353_),
    .X(net3441));
 sky130_fd_sc_hd__buf_1 wire3442 (.A(_07353_),
    .X(net3442));
 sky130_fd_sc_hd__buf_1 wire3443 (.A(_07303_),
    .X(net3443));
 sky130_fd_sc_hd__buf_1 wire3444 (.A(_07245_),
    .X(net3444));
 sky130_fd_sc_hd__clkbuf_1 wire3445 (.A(net3446),
    .X(net3445));
 sky130_fd_sc_hd__buf_1 wire3446 (.A(_07245_),
    .X(net3446));
 sky130_fd_sc_hd__buf_1 wire3447 (.A(net3448),
    .X(net3447));
 sky130_fd_sc_hd__buf_1 max_length3448 (.A(net3449),
    .X(net3448));
 sky130_fd_sc_hd__buf_1 max_length3449 (.A(net3450),
    .X(net3449));
 sky130_fd_sc_hd__buf_1 wire3450 (.A(_07230_),
    .X(net3450));
 sky130_fd_sc_hd__buf_1 wire3451 (.A(net3452),
    .X(net3451));
 sky130_fd_sc_hd__clkbuf_1 max_length3452 (.A(_07230_),
    .X(net3452));
 sky130_fd_sc_hd__buf_1 wire3453 (.A(_07194_),
    .X(net3453));
 sky130_fd_sc_hd__clkbuf_1 wire3454 (.A(net3455),
    .X(net3454));
 sky130_fd_sc_hd__buf_1 wire3455 (.A(net3456),
    .X(net3455));
 sky130_fd_sc_hd__buf_1 wire3456 (.A(net3457),
    .X(net3456));
 sky130_fd_sc_hd__clkbuf_1 wire3457 (.A(_07192_),
    .X(net3457));
 sky130_fd_sc_hd__buf_1 wire3458 (.A(net3460),
    .X(net3458));
 sky130_fd_sc_hd__clkbuf_1 max_length3459 (.A(net3460),
    .X(net3459));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3460 (.A(net3463),
    .X(net3460));
 sky130_fd_sc_hd__clkbuf_1 wire3461 (.A(net3462),
    .X(net3461));
 sky130_fd_sc_hd__buf_1 wire3462 (.A(_07189_),
    .X(net3462));
 sky130_fd_sc_hd__clkbuf_1 max_length3463 (.A(_07189_),
    .X(net3463));
 sky130_fd_sc_hd__buf_1 wire3464 (.A(_07179_),
    .X(net3464));
 sky130_fd_sc_hd__buf_1 wire3465 (.A(net3466),
    .X(net3465));
 sky130_fd_sc_hd__buf_1 wire3466 (.A(_07157_),
    .X(net3466));
 sky130_fd_sc_hd__buf_1 max_length3467 (.A(net3468),
    .X(net3467));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3468 (.A(net3469),
    .X(net3468));
 sky130_fd_sc_hd__clkbuf_1 wire3469 (.A(net3470),
    .X(net3469));
 sky130_fd_sc_hd__clkbuf_1 wire3470 (.A(_07152_),
    .X(net3470));
 sky130_fd_sc_hd__buf_1 wire3471 (.A(net3472),
    .X(net3471));
 sky130_fd_sc_hd__clkbuf_1 wire3472 (.A(net3473),
    .X(net3472));
 sky130_fd_sc_hd__clkbuf_1 max_length3473 (.A(_07152_),
    .X(net3473));
 sky130_fd_sc_hd__buf_1 max_length3474 (.A(net3475),
    .X(net3474));
 sky130_fd_sc_hd__buf_1 wire3475 (.A(net3476),
    .X(net3475));
 sky130_fd_sc_hd__clkbuf_1 wire3476 (.A(net3477),
    .X(net3476));
 sky130_fd_sc_hd__clkbuf_1 wire3477 (.A(_07151_),
    .X(net3477));
 sky130_fd_sc_hd__buf_1 wire3478 (.A(net3479),
    .X(net3478));
 sky130_fd_sc_hd__clkbuf_1 wire3479 (.A(net3480),
    .X(net3479));
 sky130_fd_sc_hd__clkbuf_1 max_length3480 (.A(_07151_),
    .X(net3480));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3481 (.A(net3482),
    .X(net3481));
 sky130_fd_sc_hd__buf_1 max_length3482 (.A(net3483),
    .X(net3482));
 sky130_fd_sc_hd__buf_1 wire3483 (.A(_07150_),
    .X(net3483));
 sky130_fd_sc_hd__clkbuf_1 wire3484 (.A(net3485),
    .X(net3484));
 sky130_fd_sc_hd__clkbuf_1 wire3485 (.A(_07150_),
    .X(net3485));
 sky130_fd_sc_hd__buf_1 wire3486 (.A(net3487),
    .X(net3486));
 sky130_fd_sc_hd__buf_1 wire3487 (.A(_07141_),
    .X(net3487));
 sky130_fd_sc_hd__buf_1 max_length3488 (.A(net3489),
    .X(net3488));
 sky130_fd_sc_hd__buf_1 wire3489 (.A(net3490),
    .X(net3489));
 sky130_fd_sc_hd__clkbuf_1 wire3490 (.A(net3491),
    .X(net3490));
 sky130_fd_sc_hd__clkbuf_1 wire3491 (.A(_07137_),
    .X(net3491));
 sky130_fd_sc_hd__buf_1 wire3492 (.A(net3493),
    .X(net3492));
 sky130_fd_sc_hd__clkbuf_1 wire3493 (.A(net3494),
    .X(net3493));
 sky130_fd_sc_hd__buf_1 wire3494 (.A(_07118_),
    .X(net3494));
 sky130_fd_sc_hd__buf_1 wire3495 (.A(_07107_),
    .X(net3495));
 sky130_fd_sc_hd__clkbuf_1 max_length3496 (.A(net3501),
    .X(net3496));
 sky130_fd_sc_hd__buf_1 wire3497 (.A(net3498),
    .X(net3497));
 sky130_fd_sc_hd__buf_1 wire3498 (.A(net3499),
    .X(net3498));
 sky130_fd_sc_hd__clkbuf_2 wire3499 (.A(net3500),
    .X(net3499));
 sky130_fd_sc_hd__clkbuf_1 wire3500 (.A(net3501),
    .X(net3500));
 sky130_fd_sc_hd__buf_1 wire3501 (.A(_07106_),
    .X(net3501));
 sky130_fd_sc_hd__buf_1 wire3502 (.A(net3503),
    .X(net3502));
 sky130_fd_sc_hd__buf_1 max_length3503 (.A(_07101_),
    .X(net3503));
 sky130_fd_sc_hd__clkbuf_1 wire3504 (.A(net3505),
    .X(net3504));
 sky130_fd_sc_hd__buf_1 wire3505 (.A(net3508),
    .X(net3505));
 sky130_fd_sc_hd__buf_1 max_length3506 (.A(net3507),
    .X(net3506));
 sky130_fd_sc_hd__buf_1 wire3507 (.A(_07096_),
    .X(net3507));
 sky130_fd_sc_hd__buf_1 max_length3508 (.A(_07096_),
    .X(net3508));
 sky130_fd_sc_hd__clkbuf_1 wire3509 (.A(net3510),
    .X(net3509));
 sky130_fd_sc_hd__buf_1 wire3510 (.A(net3513),
    .X(net3510));
 sky130_fd_sc_hd__buf_1 max_length3511 (.A(net3512),
    .X(net3511));
 sky130_fd_sc_hd__buf_1 wire3512 (.A(_07095_),
    .X(net3512));
 sky130_fd_sc_hd__buf_1 max_length3513 (.A(_07095_),
    .X(net3513));
 sky130_fd_sc_hd__clkbuf_1 wire3514 (.A(net3518),
    .X(net3514));
 sky130_fd_sc_hd__clkbuf_1 wire3515 (.A(net3517),
    .X(net3515));
 sky130_fd_sc_hd__buf_1 wire3516 (.A(net3517),
    .X(net3516));
 sky130_fd_sc_hd__buf_1 wire3517 (.A(net3518),
    .X(net3517));
 sky130_fd_sc_hd__buf_1 wire3518 (.A(net3519),
    .X(net3518));
 sky130_fd_sc_hd__clkbuf_1 wire3519 (.A(net3520),
    .X(net3519));
 sky130_fd_sc_hd__clkbuf_1 wire3520 (.A(_07066_),
    .X(net3520));
 sky130_fd_sc_hd__buf_1 max_length3521 (.A(_07066_),
    .X(net3521));
 sky130_fd_sc_hd__buf_1 wire3522 (.A(net3523),
    .X(net3522));
 sky130_fd_sc_hd__buf_1 wire3523 (.A(net3524),
    .X(net3523));
 sky130_fd_sc_hd__clkbuf_1 wire3524 (.A(net3525),
    .X(net3524));
 sky130_fd_sc_hd__buf_1 wire3525 (.A(_07063_),
    .X(net3525));
 sky130_fd_sc_hd__buf_1 wire3526 (.A(net3527),
    .X(net3526));
 sky130_fd_sc_hd__buf_1 wire3527 (.A(_07062_),
    .X(net3527));
 sky130_fd_sc_hd__buf_1 wire3528 (.A(net3529),
    .X(net3528));
 sky130_fd_sc_hd__buf_1 wire3529 (.A(_07062_),
    .X(net3529));
 sky130_fd_sc_hd__clkbuf_1 wire3530 (.A(net3531),
    .X(net3530));
 sky130_fd_sc_hd__buf_1 max_length3531 (.A(net3532),
    .X(net3531));
 sky130_fd_sc_hd__buf_1 wire3532 (.A(net3534),
    .X(net3532));
 sky130_fd_sc_hd__clkbuf_1 wire3533 (.A(net3535),
    .X(net3533));
 sky130_fd_sc_hd__buf_1 max_length3534 (.A(net3535),
    .X(net3534));
 sky130_fd_sc_hd__buf_1 wire3535 (.A(net3536),
    .X(net3535));
 sky130_fd_sc_hd__buf_1 wire3536 (.A(_07061_),
    .X(net3536));
 sky130_fd_sc_hd__buf_1 wire3537 (.A(net3538),
    .X(net3537));
 sky130_fd_sc_hd__clkbuf_1 wire3538 (.A(_07055_),
    .X(net3538));
 sky130_fd_sc_hd__buf_1 wire3539 (.A(net3540),
    .X(net3539));
 sky130_fd_sc_hd__clkbuf_1 wire3540 (.A(_07049_),
    .X(net3540));
 sky130_fd_sc_hd__buf_1 wire3541 (.A(net3542),
    .X(net3541));
 sky130_fd_sc_hd__clkbuf_1 wire3542 (.A(net3543),
    .X(net3542));
 sky130_fd_sc_hd__clkbuf_1 wire3543 (.A(_07048_),
    .X(net3543));
 sky130_fd_sc_hd__clkbuf_2 wire3544 (.A(_07047_),
    .X(net3544));
 sky130_fd_sc_hd__buf_1 wire3545 (.A(net3549),
    .X(net3545));
 sky130_fd_sc_hd__buf_1 wire3546 (.A(net3547),
    .X(net3546));
 sky130_fd_sc_hd__clkbuf_1 wire3547 (.A(net3548),
    .X(net3547));
 sky130_fd_sc_hd__clkbuf_1 wire3548 (.A(net3549),
    .X(net3548));
 sky130_fd_sc_hd__buf_1 wire3549 (.A(_07044_),
    .X(net3549));
 sky130_fd_sc_hd__buf_1 wire3550 (.A(net3551),
    .X(net3550));
 sky130_fd_sc_hd__buf_1 wire3551 (.A(net3552),
    .X(net3551));
 sky130_fd_sc_hd__buf_1 wire3552 (.A(net3553),
    .X(net3552));
 sky130_fd_sc_hd__buf_1 wire3553 (.A(_07043_),
    .X(net3553));
 sky130_fd_sc_hd__buf_1 wire3554 (.A(net3555),
    .X(net3554));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length3555 (.A(_07042_),
    .X(net3555));
 sky130_fd_sc_hd__buf_1 wire3556 (.A(net3557),
    .X(net3556));
 sky130_fd_sc_hd__buf_1 wire3557 (.A(net3558),
    .X(net3557));
 sky130_fd_sc_hd__buf_1 wire3558 (.A(_07039_),
    .X(net3558));
 sky130_fd_sc_hd__buf_1 wire3559 (.A(net3560),
    .X(net3559));
 sky130_fd_sc_hd__buf_1 max_length3560 (.A(_07038_),
    .X(net3560));
 sky130_fd_sc_hd__buf_1 wire3561 (.A(_07035_),
    .X(net3561));
 sky130_fd_sc_hd__buf_1 wire3562 (.A(net3563),
    .X(net3562));
 sky130_fd_sc_hd__clkbuf_1 wire3563 (.A(net3564),
    .X(net3563));
 sky130_fd_sc_hd__clkbuf_1 max_length3564 (.A(_07035_),
    .X(net3564));
 sky130_fd_sc_hd__clkbuf_1 wire3565 (.A(net3566),
    .X(net3565));
 sky130_fd_sc_hd__buf_1 wire3566 (.A(net3567),
    .X(net3566));
 sky130_fd_sc_hd__buf_1 wire3567 (.A(net3568),
    .X(net3567));
 sky130_fd_sc_hd__buf_1 wire3568 (.A(_07034_),
    .X(net3568));
 sky130_fd_sc_hd__buf_1 wire3569 (.A(net3570),
    .X(net3569));
 sky130_fd_sc_hd__buf_1 wire3570 (.A(net3572),
    .X(net3570));
 sky130_fd_sc_hd__clkbuf_1 max_length3571 (.A(net3572),
    .X(net3571));
 sky130_fd_sc_hd__buf_1 wire3572 (.A(_07028_),
    .X(net3572));
 sky130_fd_sc_hd__buf_1 wire3573 (.A(net3574),
    .X(net3573));
 sky130_fd_sc_hd__buf_1 wire3574 (.A(net3576),
    .X(net3574));
 sky130_fd_sc_hd__clkbuf_1 max_length3575 (.A(net3576),
    .X(net3575));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3576 (.A(_07026_),
    .X(net3576));
 sky130_fd_sc_hd__buf_1 max_length3577 (.A(net3578),
    .X(net3577));
 sky130_fd_sc_hd__buf_1 wire3578 (.A(net3579),
    .X(net3578));
 sky130_fd_sc_hd__buf_1 wire3579 (.A(_07021_),
    .X(net3579));
 sky130_fd_sc_hd__buf_1 wire3580 (.A(net3581),
    .X(net3580));
 sky130_fd_sc_hd__buf_1 wire3581 (.A(_07021_),
    .X(net3581));
 sky130_fd_sc_hd__buf_1 wire3582 (.A(net3583),
    .X(net3582));
 sky130_fd_sc_hd__buf_1 wire3583 (.A(_07019_),
    .X(net3583));
 sky130_fd_sc_hd__buf_1 max_length3584 (.A(net3585),
    .X(net3584));
 sky130_fd_sc_hd__buf_1 wire3585 (.A(net3586),
    .X(net3585));
 sky130_fd_sc_hd__buf_1 wire3586 (.A(_07019_),
    .X(net3586));
 sky130_fd_sc_hd__buf_1 wire3587 (.A(net3588),
    .X(net3587));
 sky130_fd_sc_hd__clkbuf_1 wire3588 (.A(net3589),
    .X(net3588));
 sky130_fd_sc_hd__clkbuf_1 wire3589 (.A(_06989_),
    .X(net3589));
 sky130_fd_sc_hd__clkbuf_1 max_length3590 (.A(net3591),
    .X(net3590));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3591 (.A(net3593),
    .X(net3591));
 sky130_fd_sc_hd__buf_1 wire3592 (.A(net3593),
    .X(net3592));
 sky130_fd_sc_hd__buf_1 wire3593 (.A(_06985_),
    .X(net3593));
 sky130_fd_sc_hd__buf_1 wire3594 (.A(net3595),
    .X(net3594));
 sky130_fd_sc_hd__buf_1 wire3595 (.A(_06984_),
    .X(net3595));
 sky130_fd_sc_hd__clkbuf_1 max_length3596 (.A(net3597),
    .X(net3596));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3597 (.A(_06984_),
    .X(net3597));
 sky130_fd_sc_hd__buf_1 wire3598 (.A(_06973_),
    .X(net3598));
 sky130_fd_sc_hd__buf_1 wire3599 (.A(net3600),
    .X(net3599));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3600 (.A(net3601),
    .X(net3600));
 sky130_fd_sc_hd__buf_1 wire3601 (.A(_06967_),
    .X(net3601));
 sky130_fd_sc_hd__buf_1 wire3602 (.A(net3603),
    .X(net3602));
 sky130_fd_sc_hd__buf_1 max_length3603 (.A(_06964_),
    .X(net3603));
 sky130_fd_sc_hd__clkbuf_2 wire3604 (.A(net3605),
    .X(net3604));
 sky130_fd_sc_hd__buf_1 max_length3605 (.A(net3606),
    .X(net3605));
 sky130_fd_sc_hd__clkbuf_2 wire3606 (.A(_06950_),
    .X(net3606));
 sky130_fd_sc_hd__clkbuf_2 wire3607 (.A(net3608),
    .X(net3607));
 sky130_fd_sc_hd__clkbuf_2 max_length3608 (.A(net3609),
    .X(net3608));
 sky130_fd_sc_hd__buf_1 max_length3609 (.A(_06939_),
    .X(net3609));
 sky130_fd_sc_hd__clkbuf_2 wire3610 (.A(net3611),
    .X(net3610));
 sky130_fd_sc_hd__buf_1 wire3611 (.A(_06928_),
    .X(net3611));
 sky130_fd_sc_hd__buf_1 max_length3612 (.A(_06928_),
    .X(net3612));
 sky130_fd_sc_hd__buf_1 max_length3613 (.A(net3614),
    .X(net3613));
 sky130_fd_sc_hd__buf_1 wire3614 (.A(net3615),
    .X(net3614));
 sky130_fd_sc_hd__buf_1 wire3615 (.A(_06862_),
    .X(net3615));
 sky130_fd_sc_hd__buf_1 wire3616 (.A(_06862_),
    .X(net3616));
 sky130_fd_sc_hd__clkbuf_1 wire3617 (.A(_06831_),
    .X(net3617));
 sky130_fd_sc_hd__buf_1 wire3618 (.A(net3619),
    .X(net3618));
 sky130_fd_sc_hd__buf_1 wire3619 (.A(net3620),
    .X(net3619));
 sky130_fd_sc_hd__buf_1 wire3620 (.A(net3621),
    .X(net3620));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3621 (.A(_06823_),
    .X(net3621));
 sky130_fd_sc_hd__clkbuf_1 wire3622 (.A(_06823_),
    .X(net3622));
 sky130_fd_sc_hd__clkbuf_1 max_length3623 (.A(_06823_),
    .X(net3623));
 sky130_fd_sc_hd__buf_1 wire3624 (.A(net3625),
    .X(net3624));
 sky130_fd_sc_hd__buf_1 wire3625 (.A(_06818_),
    .X(net3625));
 sky130_fd_sc_hd__clkbuf_1 wire3626 (.A(_06818_),
    .X(net3626));
 sky130_fd_sc_hd__buf_1 wire3627 (.A(net3628),
    .X(net3627));
 sky130_fd_sc_hd__buf_1 wire3628 (.A(net3629),
    .X(net3628));
 sky130_fd_sc_hd__buf_1 wire3629 (.A(_06800_),
    .X(net3629));
 sky130_fd_sc_hd__buf_1 max_length3630 (.A(_06800_),
    .X(net3630));
 sky130_fd_sc_hd__buf_1 wire3631 (.A(net3632),
    .X(net3631));
 sky130_fd_sc_hd__buf_1 wire3632 (.A(net3634),
    .X(net3632));
 sky130_fd_sc_hd__buf_1 wire3633 (.A(net3634),
    .X(net3633));
 sky130_fd_sc_hd__buf_1 wire3634 (.A(_06609_),
    .X(net3634));
 sky130_fd_sc_hd__buf_1 wire3635 (.A(net3636),
    .X(net3635));
 sky130_fd_sc_hd__buf_1 wire3636 (.A(_06575_),
    .X(net3636));
 sky130_fd_sc_hd__buf_1 wire3637 (.A(_06575_),
    .X(net3637));
 sky130_fd_sc_hd__clkbuf_1 wire3638 (.A(net3639),
    .X(net3638));
 sky130_fd_sc_hd__buf_1 wire3639 (.A(net3640),
    .X(net3639));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3640 (.A(net3641),
    .X(net3640));
 sky130_fd_sc_hd__buf_1 wire3641 (.A(_06533_),
    .X(net3641));
 sky130_fd_sc_hd__buf_1 max_length3642 (.A(net3643),
    .X(net3642));
 sky130_fd_sc_hd__buf_1 wire3643 (.A(net3644),
    .X(net3643));
 sky130_fd_sc_hd__clkbuf_1 wire3644 (.A(net3645),
    .X(net3644));
 sky130_fd_sc_hd__buf_1 wire3645 (.A(net3646),
    .X(net3645));
 sky130_fd_sc_hd__buf_1 wire3646 (.A(_06527_),
    .X(net3646));
 sky130_fd_sc_hd__buf_1 wire3647 (.A(net3648),
    .X(net3647));
 sky130_fd_sc_hd__buf_1 wire3648 (.A(_06524_),
    .X(net3648));
 sky130_fd_sc_hd__buf_1 wire3649 (.A(net3650),
    .X(net3649));
 sky130_fd_sc_hd__clkbuf_1 wire3650 (.A(net3651),
    .X(net3650));
 sky130_fd_sc_hd__clkbuf_1 wire3651 (.A(net3652),
    .X(net3651));
 sky130_fd_sc_hd__clkbuf_1 wire3652 (.A(net3653),
    .X(net3652));
 sky130_fd_sc_hd__clkbuf_1 wire3653 (.A(net3654),
    .X(net3653));
 sky130_fd_sc_hd__clkbuf_1 wire3654 (.A(net3655),
    .X(net3654));
 sky130_fd_sc_hd__clkbuf_1 wire3655 (.A(net3656),
    .X(net3655));
 sky130_fd_sc_hd__clkbuf_1 wire3656 (.A(net3666),
    .X(net3656));
 sky130_fd_sc_hd__clkbuf_1 wire3657 (.A(net3658),
    .X(net3657));
 sky130_fd_sc_hd__buf_1 wire3658 (.A(net3659),
    .X(net3658));
 sky130_fd_sc_hd__clkbuf_1 wire3659 (.A(net3660),
    .X(net3659));
 sky130_fd_sc_hd__clkbuf_1 wire3660 (.A(net3661),
    .X(net3660));
 sky130_fd_sc_hd__clkbuf_1 wire3661 (.A(net3662),
    .X(net3661));
 sky130_fd_sc_hd__clkbuf_1 wire3662 (.A(net3663),
    .X(net3662));
 sky130_fd_sc_hd__clkbuf_1 wire3663 (.A(net3664),
    .X(net3663));
 sky130_fd_sc_hd__clkbuf_1 wire3664 (.A(net3665),
    .X(net3664));
 sky130_fd_sc_hd__clkbuf_1 wire3665 (.A(_06510_),
    .X(net3665));
 sky130_fd_sc_hd__clkbuf_1 max_length3666 (.A(_06510_),
    .X(net3666));
 sky130_fd_sc_hd__buf_1 max_length3667 (.A(net3668),
    .X(net3667));
 sky130_fd_sc_hd__buf_1 wire3668 (.A(_06505_),
    .X(net3668));
 sky130_fd_sc_hd__buf_1 wire3669 (.A(net3670),
    .X(net3669));
 sky130_fd_sc_hd__buf_1 wire3670 (.A(net3671),
    .X(net3670));
 sky130_fd_sc_hd__clkbuf_1 wire3671 (.A(net3672),
    .X(net3671));
 sky130_fd_sc_hd__clkbuf_1 wire3672 (.A(net3673),
    .X(net3672));
 sky130_fd_sc_hd__buf_1 wire3673 (.A(net3674),
    .X(net3673));
 sky130_fd_sc_hd__buf_1 wire3674 (.A(_05709_),
    .X(net3674));
 sky130_fd_sc_hd__buf_1 wire3675 (.A(_05616_),
    .X(net3675));
 sky130_fd_sc_hd__buf_1 max_length3676 (.A(net3677),
    .X(net3676));
 sky130_fd_sc_hd__buf_1 wire3677 (.A(net3678),
    .X(net3677));
 sky130_fd_sc_hd__buf_1 wire3678 (.A(net3679),
    .X(net3678));
 sky130_fd_sc_hd__buf_1 wire3679 (.A(net3680),
    .X(net3679));
 sky130_fd_sc_hd__clkbuf_1 wire3680 (.A(net3681),
    .X(net3680));
 sky130_fd_sc_hd__clkbuf_1 wire3681 (.A(_05615_),
    .X(net3681));
 sky130_fd_sc_hd__buf_1 wire3682 (.A(net3683),
    .X(net3682));
 sky130_fd_sc_hd__clkbuf_1 wire3683 (.A(_05531_),
    .X(net3683));
 sky130_fd_sc_hd__clkbuf_1 wire3684 (.A(_05345_),
    .X(net3684));
 sky130_fd_sc_hd__buf_1 wire3685 (.A(net3686),
    .X(net3685));
 sky130_fd_sc_hd__buf_1 wire3686 (.A(net3687),
    .X(net3686));
 sky130_fd_sc_hd__buf_1 wire3687 (.A(_05053_),
    .X(net3687));
 sky130_fd_sc_hd__buf_1 wire3688 (.A(net3692),
    .X(net3688));
 sky130_fd_sc_hd__buf_1 wire3689 (.A(net3690),
    .X(net3689));
 sky130_fd_sc_hd__clkbuf_1 wire3690 (.A(net3691),
    .X(net3690));
 sky130_fd_sc_hd__clkbuf_1 wire3691 (.A(net3692),
    .X(net3691));
 sky130_fd_sc_hd__clkbuf_1 wire3692 (.A(_05022_),
    .X(net3692));
 sky130_fd_sc_hd__buf_1 wire3693 (.A(_04897_),
    .X(net3693));
 sky130_fd_sc_hd__buf_1 wire3694 (.A(_04897_),
    .X(net3694));
 sky130_fd_sc_hd__clkbuf_2 wire3695 (.A(_04894_),
    .X(net3695));
 sky130_fd_sc_hd__buf_1 wire3696 (.A(_04886_),
    .X(net3696));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3697 (.A(_04884_),
    .X(net3697));
 sky130_fd_sc_hd__clkbuf_1 max_length3698 (.A(_04884_),
    .X(net3698));
 sky130_fd_sc_hd__buf_1 wire3699 (.A(net3700),
    .X(net3699));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3700 (.A(net3701),
    .X(net3700));
 sky130_fd_sc_hd__buf_1 wire3701 (.A(_04882_),
    .X(net3701));
 sky130_fd_sc_hd__clkbuf_2 wire3702 (.A(net3703),
    .X(net3702));
 sky130_fd_sc_hd__buf_1 wire3703 (.A(net3704),
    .X(net3703));
 sky130_fd_sc_hd__buf_1 wire3704 (.A(_04877_),
    .X(net3704));
 sky130_fd_sc_hd__clkbuf_2 wire3705 (.A(net3706),
    .X(net3705));
 sky130_fd_sc_hd__clkbuf_1 wire3706 (.A(net3707),
    .X(net3706));
 sky130_fd_sc_hd__clkbuf_1 wire3707 (.A(net3708),
    .X(net3707));
 sky130_fd_sc_hd__clkbuf_1 wire3708 (.A(net3709),
    .X(net3708));
 sky130_fd_sc_hd__buf_1 wire3709 (.A(_04873_),
    .X(net3709));
 sky130_fd_sc_hd__buf_1 wire3710 (.A(net3711),
    .X(net3710));
 sky130_fd_sc_hd__clkbuf_2 wire3711 (.A(net3712),
    .X(net3711));
 sky130_fd_sc_hd__clkbuf_1 wire3712 (.A(net3713),
    .X(net3712));
 sky130_fd_sc_hd__clkbuf_1 wire3713 (.A(net3714),
    .X(net3713));
 sky130_fd_sc_hd__clkbuf_1 wire3714 (.A(net3715),
    .X(net3714));
 sky130_fd_sc_hd__buf_1 wire3715 (.A(_04869_),
    .X(net3715));
 sky130_fd_sc_hd__clkbuf_1 max_length3716 (.A(_04869_),
    .X(net3716));
 sky130_fd_sc_hd__clkbuf_1 wire3717 (.A(_04867_),
    .X(net3717));
 sky130_fd_sc_hd__buf_1 wire3718 (.A(net3719),
    .X(net3718));
 sky130_fd_sc_hd__buf_1 wire3719 (.A(net3720),
    .X(net3719));
 sky130_fd_sc_hd__clkbuf_1 wire3720 (.A(net3721),
    .X(net3720));
 sky130_fd_sc_hd__clkbuf_1 wire3721 (.A(net3722),
    .X(net3721));
 sky130_fd_sc_hd__clkbuf_1 wire3722 (.A(net3723),
    .X(net3722));
 sky130_fd_sc_hd__clkbuf_1 wire3723 (.A(net3724),
    .X(net3723));
 sky130_fd_sc_hd__clkbuf_1 wire3724 (.A(net3725),
    .X(net3724));
 sky130_fd_sc_hd__clkbuf_1 wire3725 (.A(net3726),
    .X(net3725));
 sky130_fd_sc_hd__clkbuf_1 wire3726 (.A(_04867_),
    .X(net3726));
 sky130_fd_sc_hd__buf_1 wire3727 (.A(net3728),
    .X(net3727));
 sky130_fd_sc_hd__clkbuf_1 wire3728 (.A(net3729),
    .X(net3728));
 sky130_fd_sc_hd__clkbuf_1 wire3729 (.A(_04531_),
    .X(net3729));
 sky130_fd_sc_hd__buf_1 max_length3730 (.A(_04531_),
    .X(net3730));
 sky130_fd_sc_hd__buf_1 wire3731 (.A(_04502_),
    .X(net3731));
 sky130_fd_sc_hd__buf_1 wire3732 (.A(net3733),
    .X(net3732));
 sky130_fd_sc_hd__clkbuf_1 wire3733 (.A(_04172_),
    .X(net3733));
 sky130_fd_sc_hd__buf_1 wire3734 (.A(net3735),
    .X(net3734));
 sky130_fd_sc_hd__clkbuf_1 wire3735 (.A(net3736),
    .X(net3735));
 sky130_fd_sc_hd__buf_1 max_length3736 (.A(_04117_),
    .X(net3736));
 sky130_fd_sc_hd__buf_1 wire3737 (.A(_04038_),
    .X(net3737));
 sky130_fd_sc_hd__buf_1 wire3738 (.A(_03861_),
    .X(net3738));
 sky130_fd_sc_hd__buf_1 wire3739 (.A(net3740),
    .X(net3739));
 sky130_fd_sc_hd__clkbuf_1 wire3740 (.A(_03771_),
    .X(net3740));
 sky130_fd_sc_hd__buf_1 wire3741 (.A(net3742),
    .X(net3741));
 sky130_fd_sc_hd__buf_1 max_length3742 (.A(_03705_),
    .X(net3742));
 sky130_fd_sc_hd__clkbuf_2 wire3743 (.A(_03608_),
    .X(net3743));
 sky130_fd_sc_hd__buf_1 wire3744 (.A(net3745),
    .X(net3744));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3745 (.A(_03605_),
    .X(net3745));
 sky130_fd_sc_hd__clkbuf_1 wire3746 (.A(_03456_),
    .X(net3746));
 sky130_fd_sc_hd__buf_1 wire3747 (.A(_03456_),
    .X(net3747));
 sky130_fd_sc_hd__buf_1 max_length3748 (.A(_03456_),
    .X(net3748));
 sky130_fd_sc_hd__clkbuf_2 wire3749 (.A(_03074_),
    .X(net3749));
 sky130_fd_sc_hd__clkbuf_1 wire3750 (.A(net3751),
    .X(net3750));
 sky130_fd_sc_hd__clkbuf_1 wire3751 (.A(net3752),
    .X(net3751));
 sky130_fd_sc_hd__buf_1 wire3752 (.A(_03065_),
    .X(net3752));
 sky130_fd_sc_hd__buf_1 wire3753 (.A(net3754),
    .X(net3753));
 sky130_fd_sc_hd__clkbuf_1 wire3754 (.A(net3755),
    .X(net3754));
 sky130_fd_sc_hd__clkbuf_1 wire3755 (.A(net3756),
    .X(net3755));
 sky130_fd_sc_hd__clkbuf_1 max_length3756 (.A(_02925_),
    .X(net3756));
 sky130_fd_sc_hd__buf_1 wire3757 (.A(_02866_),
    .X(net3757));
 sky130_fd_sc_hd__buf_1 max_length3758 (.A(_02866_),
    .X(net3758));
 sky130_fd_sc_hd__buf_1 wire3759 (.A(net3760),
    .X(net3759));
 sky130_fd_sc_hd__clkbuf_1 wire3760 (.A(net3761),
    .X(net3760));
 sky130_fd_sc_hd__buf_1 wire3761 (.A(net3762),
    .X(net3761));
 sky130_fd_sc_hd__buf_1 wire3762 (.A(_02716_),
    .X(net3762));
 sky130_fd_sc_hd__clkbuf_1 wire3763 (.A(_02712_),
    .X(net3763));
 sky130_fd_sc_hd__buf_1 wire3764 (.A(net3765),
    .X(net3764));
 sky130_fd_sc_hd__clkbuf_1 wire3765 (.A(net3766),
    .X(net3765));
 sky130_fd_sc_hd__clkbuf_1 wire3766 (.A(_02659_),
    .X(net3766));
 sky130_fd_sc_hd__buf_1 wire3767 (.A(_02560_),
    .X(net3767));
 sky130_fd_sc_hd__buf_1 max_length3768 (.A(net3769),
    .X(net3768));
 sky130_fd_sc_hd__buf_1 wire3769 (.A(net3770),
    .X(net3769));
 sky130_fd_sc_hd__buf_1 wire3770 (.A(net3771),
    .X(net3770));
 sky130_fd_sc_hd__clkbuf_1 wire3771 (.A(net3772),
    .X(net3771));
 sky130_fd_sc_hd__clkbuf_1 wire3772 (.A(net3773),
    .X(net3772));
 sky130_fd_sc_hd__clkbuf_1 wire3773 (.A(_02545_),
    .X(net3773));
 sky130_fd_sc_hd__buf_1 wire3774 (.A(_02541_),
    .X(net3774));
 sky130_fd_sc_hd__buf_1 max_length3775 (.A(_02541_),
    .X(net3775));
 sky130_fd_sc_hd__buf_1 wire3776 (.A(_01873_),
    .X(net3776));
 sky130_fd_sc_hd__clkbuf_1 wire3777 (.A(net3779),
    .X(net3777));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3778 (.A(net3779),
    .X(net3778));
 sky130_fd_sc_hd__buf_1 max_length3779 (.A(_01873_),
    .X(net3779));
 sky130_fd_sc_hd__buf_1 wire3780 (.A(net3781),
    .X(net3780));
 sky130_fd_sc_hd__clkbuf_1 wire3781 (.A(net3782),
    .X(net3781));
 sky130_fd_sc_hd__clkbuf_1 wire3782 (.A(net3783),
    .X(net3782));
 sky130_fd_sc_hd__clkbuf_1 wire3783 (.A(net3784),
    .X(net3783));
 sky130_fd_sc_hd__clkbuf_1 wire3784 (.A(_01863_),
    .X(net3784));
 sky130_fd_sc_hd__clkbuf_1 wire3785 (.A(net3787),
    .X(net3785));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3786 (.A(net3788),
    .X(net3786));
 sky130_fd_sc_hd__buf_1 max_length3787 (.A(net3788),
    .X(net3787));
 sky130_fd_sc_hd__buf_1 wire3788 (.A(_01709_),
    .X(net3788));
 sky130_fd_sc_hd__buf_1 wire3789 (.A(net3790),
    .X(net3789));
 sky130_fd_sc_hd__clkbuf_1 wire3790 (.A(net3791),
    .X(net3790));
 sky130_fd_sc_hd__clkbuf_1 wire3791 (.A(net3792),
    .X(net3791));
 sky130_fd_sc_hd__clkbuf_1 wire3792 (.A(net3793),
    .X(net3792));
 sky130_fd_sc_hd__clkbuf_1 wire3793 (.A(net3794),
    .X(net3793));
 sky130_fd_sc_hd__clkbuf_1 wire3794 (.A(net3795),
    .X(net3794));
 sky130_fd_sc_hd__clkbuf_1 max_length3795 (.A(_01405_),
    .X(net3795));
 sky130_fd_sc_hd__buf_1 wire3796 (.A(net3797),
    .X(net3796));
 sky130_fd_sc_hd__clkbuf_1 wire3797 (.A(net3798),
    .X(net3797));
 sky130_fd_sc_hd__clkbuf_1 wire3798 (.A(net3799),
    .X(net3798));
 sky130_fd_sc_hd__clkbuf_1 wire3799 (.A(net3800),
    .X(net3799));
 sky130_fd_sc_hd__clkbuf_1 wire3800 (.A(net3801),
    .X(net3800));
 sky130_fd_sc_hd__clkbuf_1 wire3801 (.A(net3802),
    .X(net3801));
 sky130_fd_sc_hd__clkbuf_1 wire3802 (.A(_01317_),
    .X(net3802));
 sky130_fd_sc_hd__clkbuf_1 wire3803 (.A(net3804),
    .X(net3803));
 sky130_fd_sc_hd__clkbuf_1 wire3804 (.A(_01174_),
    .X(net3804));
 sky130_fd_sc_hd__buf_1 wire3805 (.A(_01066_),
    .X(net3805));
 sky130_fd_sc_hd__buf_1 wire3806 (.A(_01054_),
    .X(net3806));
 sky130_fd_sc_hd__buf_1 wire3807 (.A(_01049_),
    .X(net3807));
 sky130_fd_sc_hd__clkbuf_1 wire3808 (.A(net3809),
    .X(net3808));
 sky130_fd_sc_hd__clkbuf_1 wire3809 (.A(net3810),
    .X(net3809));
 sky130_fd_sc_hd__clkbuf_1 wire3810 (.A(net3811),
    .X(net3810));
 sky130_fd_sc_hd__buf_1 wire3811 (.A(net3812),
    .X(net3811));
 sky130_fd_sc_hd__buf_1 wire3812 (.A(net3813),
    .X(net3812));
 sky130_fd_sc_hd__clkbuf_1 wire3813 (.A(net3814),
    .X(net3813));
 sky130_fd_sc_hd__clkbuf_1 wire3814 (.A(net3815),
    .X(net3814));
 sky130_fd_sc_hd__clkbuf_1 wire3815 (.A(_00978_),
    .X(net3815));
 sky130_fd_sc_hd__buf_1 wire3816 (.A(net3817),
    .X(net3816));
 sky130_fd_sc_hd__clkbuf_1 wire3817 (.A(net3818),
    .X(net3817));
 sky130_fd_sc_hd__buf_1 wire3818 (.A(net3819),
    .X(net3818));
 sky130_fd_sc_hd__clkbuf_1 wire3819 (.A(net3820),
    .X(net3819));
 sky130_fd_sc_hd__clkbuf_1 wire3820 (.A(net3821),
    .X(net3820));
 sky130_fd_sc_hd__buf_1 wire3821 (.A(net3822),
    .X(net3821));
 sky130_fd_sc_hd__clkbuf_1 wire3822 (.A(_00978_),
    .X(net3822));
 sky130_fd_sc_hd__clkbuf_2 wire3823 (.A(net3824),
    .X(net3823));
 sky130_fd_sc_hd__clkbuf_1 wire3824 (.A(_00977_),
    .X(net3824));
 sky130_fd_sc_hd__clkbuf_1 wire3825 (.A(net3826),
    .X(net3825));
 sky130_fd_sc_hd__clkbuf_1 wire3826 (.A(net3827),
    .X(net3826));
 sky130_fd_sc_hd__clkbuf_1 wire3827 (.A(net3828),
    .X(net3827));
 sky130_fd_sc_hd__clkbuf_1 wire3828 (.A(_00960_),
    .X(net3828));
 sky130_fd_sc_hd__buf_1 max_length3829 (.A(_00960_),
    .X(net3829));
 sky130_fd_sc_hd__buf_1 wire3830 (.A(net3831),
    .X(net3830));
 sky130_fd_sc_hd__clkbuf_1 wire3831 (.A(net3832),
    .X(net3831));
 sky130_fd_sc_hd__clkbuf_1 wire3832 (.A(net3833),
    .X(net3832));
 sky130_fd_sc_hd__clkbuf_1 wire3833 (.A(net3834),
    .X(net3833));
 sky130_fd_sc_hd__clkbuf_1 wire3834 (.A(net3835),
    .X(net3834));
 sky130_fd_sc_hd__clkbuf_1 wire3835 (.A(_00917_),
    .X(net3835));
 sky130_fd_sc_hd__clkbuf_2 wire3836 (.A(net3837),
    .X(net3836));
 sky130_fd_sc_hd__clkbuf_1 wire3837 (.A(net3838),
    .X(net3837));
 sky130_fd_sc_hd__clkbuf_1 wire3838 (.A(_00882_),
    .X(net3838));
 sky130_fd_sc_hd__buf_1 wire3839 (.A(_00881_),
    .X(net3839));
 sky130_fd_sc_hd__buf_1 wire3840 (.A(net3841),
    .X(net3840));
 sky130_fd_sc_hd__buf_1 wire3841 (.A(_00871_),
    .X(net3841));
 sky130_fd_sc_hd__buf_1 wire3842 (.A(_00851_),
    .X(net3842));
 sky130_fd_sc_hd__buf_1 wire3843 (.A(net3844),
    .X(net3843));
 sky130_fd_sc_hd__buf_1 max_length3844 (.A(_12499_),
    .X(net3844));
 sky130_fd_sc_hd__clkbuf_1 wire3845 (.A(_12298_),
    .X(net3845));
 sky130_fd_sc_hd__buf_1 wire3846 (.A(_12296_),
    .X(net3846));
 sky130_fd_sc_hd__buf_1 wire3847 (.A(_12276_),
    .X(net3847));
 sky130_fd_sc_hd__buf_1 wire3848 (.A(_12274_),
    .X(net3848));
 sky130_fd_sc_hd__buf_1 wire3849 (.A(net3850),
    .X(net3849));
 sky130_fd_sc_hd__buf_1 max_length3850 (.A(_12269_),
    .X(net3850));
 sky130_fd_sc_hd__clkbuf_1 wire3851 (.A(_12267_),
    .X(net3851));
 sky130_fd_sc_hd__buf_1 wire3852 (.A(_12266_),
    .X(net3852));
 sky130_fd_sc_hd__buf_1 wire3853 (.A(_12265_),
    .X(net3853));
 sky130_fd_sc_hd__buf_1 wire3854 (.A(_12264_),
    .X(net3854));
 sky130_fd_sc_hd__clkbuf_1 wire3855 (.A(_11559_),
    .X(net3855));
 sky130_fd_sc_hd__buf_2 wire3856 (.A(_11559_),
    .X(net3856));
 sky130_fd_sc_hd__buf_1 wire3857 (.A(net3858),
    .X(net3857));
 sky130_fd_sc_hd__buf_1 max_length3858 (.A(net3859),
    .X(net3858));
 sky130_fd_sc_hd__buf_1 wire3859 (.A(net3860),
    .X(net3859));
 sky130_fd_sc_hd__buf_1 max_length3860 (.A(net3861),
    .X(net3860));
 sky130_fd_sc_hd__buf_1 wire3861 (.A(_11549_),
    .X(net3861));
 sky130_fd_sc_hd__buf_1 wire3862 (.A(net3863),
    .X(net3862));
 sky130_fd_sc_hd__buf_1 wire3863 (.A(_11490_),
    .X(net3863));
 sky130_fd_sc_hd__buf_1 wire3864 (.A(net3865),
    .X(net3864));
 sky130_fd_sc_hd__clkbuf_1 max_length3865 (.A(_11436_),
    .X(net3865));
 sky130_fd_sc_hd__buf_1 wire3866 (.A(_11289_),
    .X(net3866));
 sky130_fd_sc_hd__clkbuf_1 wire3867 (.A(net3868),
    .X(net3867));
 sky130_fd_sc_hd__buf_1 max_length3868 (.A(_11274_),
    .X(net3868));
 sky130_fd_sc_hd__buf_1 wire3869 (.A(_11271_),
    .X(net3869));
 sky130_fd_sc_hd__clkbuf_1 max_length3870 (.A(_11271_),
    .X(net3870));
 sky130_fd_sc_hd__clkbuf_1 wire3871 (.A(net3872),
    .X(net3871));
 sky130_fd_sc_hd__clkbuf_1 wire3872 (.A(net3873),
    .X(net3872));
 sky130_fd_sc_hd__clkbuf_1 max_length3873 (.A(_11164_),
    .X(net3873));
 sky130_fd_sc_hd__clkbuf_1 wire3874 (.A(net3875),
    .X(net3874));
 sky130_fd_sc_hd__clkbuf_1 wire3875 (.A(_11054_),
    .X(net3875));
 sky130_fd_sc_hd__clkbuf_1 wire3876 (.A(_11035_),
    .X(net3876));
 sky130_fd_sc_hd__buf_1 wire3877 (.A(_11025_),
    .X(net3877));
 sky130_fd_sc_hd__buf_1 wire3878 (.A(net3879),
    .X(net3878));
 sky130_fd_sc_hd__buf_1 max_length3879 (.A(_10996_),
    .X(net3879));
 sky130_fd_sc_hd__buf_1 wire3880 (.A(net3881),
    .X(net3880));
 sky130_fd_sc_hd__buf_1 wire3881 (.A(_10995_),
    .X(net3881));
 sky130_fd_sc_hd__clkbuf_1 wire3882 (.A(_10983_),
    .X(net3882));
 sky130_fd_sc_hd__buf_1 wire3883 (.A(_10946_),
    .X(net3883));
 sky130_fd_sc_hd__clkbuf_1 wire3884 (.A(_10943_),
    .X(net3884));
 sky130_fd_sc_hd__clkbuf_1 wire3885 (.A(_10930_),
    .X(net3885));
 sky130_fd_sc_hd__buf_1 wire3886 (.A(net3887),
    .X(net3886));
 sky130_fd_sc_hd__buf_1 max_length3887 (.A(net3888),
    .X(net3887));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3888 (.A(_10898_),
    .X(net3888));
 sky130_fd_sc_hd__clkbuf_1 wire3889 (.A(_10882_),
    .X(net3889));
 sky130_fd_sc_hd__buf_1 wire3890 (.A(_10879_),
    .X(net3890));
 sky130_fd_sc_hd__clkbuf_1 wire3891 (.A(net3892),
    .X(net3891));
 sky130_fd_sc_hd__buf_1 max_length3892 (.A(net3893),
    .X(net3892));
 sky130_fd_sc_hd__buf_1 wire3893 (.A(net3894),
    .X(net3893));
 sky130_fd_sc_hd__buf_1 wire3894 (.A(_10879_),
    .X(net3894));
 sky130_fd_sc_hd__buf_1 wire3895 (.A(_10878_),
    .X(net3895));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3896 (.A(_10878_),
    .X(net3896));
 sky130_fd_sc_hd__buf_1 wire3897 (.A(_10839_),
    .X(net3897));
 sky130_fd_sc_hd__buf_1 wire3898 (.A(_10837_),
    .X(net3898));
 sky130_fd_sc_hd__clkbuf_1 max_length3899 (.A(net3900),
    .X(net3899));
 sky130_fd_sc_hd__clkbuf_1 max_length3900 (.A(net3901),
    .X(net3900));
 sky130_fd_sc_hd__buf_1 wire3901 (.A(_10822_),
    .X(net3901));
 sky130_fd_sc_hd__buf_1 wire3902 (.A(_10813_),
    .X(net3902));
 sky130_fd_sc_hd__clkbuf_1 wire3903 (.A(_10812_),
    .X(net3903));
 sky130_fd_sc_hd__clkbuf_1 wire3904 (.A(net3905),
    .X(net3904));
 sky130_fd_sc_hd__buf_1 wire3905 (.A(_10803_),
    .X(net3905));
 sky130_fd_sc_hd__buf_1 wire3906 (.A(_10801_),
    .X(net3906));
 sky130_fd_sc_hd__buf_1 max_length3907 (.A(_10801_),
    .X(net3907));
 sky130_fd_sc_hd__buf_1 wire3908 (.A(net3909),
    .X(net3908));
 sky130_fd_sc_hd__buf_1 wire3909 (.A(_10794_),
    .X(net3909));
 sky130_fd_sc_hd__buf_1 wire3910 (.A(net3911),
    .X(net3910));
 sky130_fd_sc_hd__clkbuf_1 wire3911 (.A(net3912),
    .X(net3911));
 sky130_fd_sc_hd__clkbuf_1 wire3912 (.A(net3913),
    .X(net3912));
 sky130_fd_sc_hd__buf_1 wire3913 (.A(_10790_),
    .X(net3913));
 sky130_fd_sc_hd__clkbuf_1 wire3914 (.A(net3917),
    .X(net3914));
 sky130_fd_sc_hd__buf_1 wire3915 (.A(net3916),
    .X(net3915));
 sky130_fd_sc_hd__buf_1 wire3916 (.A(net3917),
    .X(net3916));
 sky130_fd_sc_hd__buf_1 wire3917 (.A(_10787_),
    .X(net3917));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3918 (.A(net3919),
    .X(net3918));
 sky130_fd_sc_hd__buf_1 max_length3919 (.A(_10787_),
    .X(net3919));
 sky130_fd_sc_hd__clkbuf_2 wire3920 (.A(net3921),
    .X(net3920));
 sky130_fd_sc_hd__clkbuf_1 max_length3921 (.A(_10597_),
    .X(net3921));
 sky130_fd_sc_hd__buf_1 wire3922 (.A(_10479_),
    .X(net3922));
 sky130_fd_sc_hd__buf_1 wire3923 (.A(_10335_),
    .X(net3923));
 sky130_fd_sc_hd__clkbuf_1 wire3924 (.A(_10218_),
    .X(net3924));
 sky130_fd_sc_hd__buf_1 wire3925 (.A(_10211_),
    .X(net3925));
 sky130_fd_sc_hd__buf_1 wire3926 (.A(_10123_),
    .X(net3926));
 sky130_fd_sc_hd__buf_1 wire3927 (.A(net3931),
    .X(net3927));
 sky130_fd_sc_hd__buf_1 wire3928 (.A(net3929),
    .X(net3928));
 sky130_fd_sc_hd__buf_1 wire3929 (.A(net3930),
    .X(net3929));
 sky130_fd_sc_hd__buf_1 wire3930 (.A(net3931),
    .X(net3930));
 sky130_fd_sc_hd__buf_1 wire3931 (.A(_10122_),
    .X(net3931));
 sky130_fd_sc_hd__buf_1 wire3932 (.A(_10103_),
    .X(net3932));
 sky130_fd_sc_hd__clkbuf_1 wire3933 (.A(_10094_),
    .X(net3933));
 sky130_fd_sc_hd__buf_1 wire3934 (.A(net3935),
    .X(net3934));
 sky130_fd_sc_hd__clkbuf_1 wire3935 (.A(_10064_),
    .X(net3935));
 sky130_fd_sc_hd__buf_1 wire3936 (.A(net3937),
    .X(net3936));
 sky130_fd_sc_hd__clkbuf_1 wire3937 (.A(net3939),
    .X(net3937));
 sky130_fd_sc_hd__clkbuf_1 wire3938 (.A(_10045_),
    .X(net3938));
 sky130_fd_sc_hd__clkbuf_1 max_length3939 (.A(_10045_),
    .X(net3939));
 sky130_fd_sc_hd__clkbuf_1 wire3940 (.A(_09934_),
    .X(net3940));
 sky130_fd_sc_hd__buf_1 wire3941 (.A(_09934_),
    .X(net3941));
 sky130_fd_sc_hd__buf_1 wire3942 (.A(_09910_),
    .X(net3942));
 sky130_fd_sc_hd__clkbuf_1 wire3943 (.A(net3944),
    .X(net3943));
 sky130_fd_sc_hd__clkbuf_1 wire3944 (.A(net3946),
    .X(net3944));
 sky130_fd_sc_hd__clkbuf_1 wire3945 (.A(_09879_),
    .X(net3945));
 sky130_fd_sc_hd__clkbuf_1 max_length3946 (.A(_09879_),
    .X(net3946));
 sky130_fd_sc_hd__buf_1 wire3947 (.A(net3948),
    .X(net3947));
 sky130_fd_sc_hd__buf_1 wire3948 (.A(net3951),
    .X(net3948));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3949 (.A(net3950),
    .X(net3949));
 sky130_fd_sc_hd__clkbuf_1 wire3950 (.A(_09876_),
    .X(net3950));
 sky130_fd_sc_hd__clkbuf_1 max_length3951 (.A(_09876_),
    .X(net3951));
 sky130_fd_sc_hd__clkbuf_2 wire3952 (.A(_09808_),
    .X(net3952));
 sky130_fd_sc_hd__clkbuf_1 wire3953 (.A(net3954),
    .X(net3953));
 sky130_fd_sc_hd__clkbuf_1 wire3954 (.A(net3955),
    .X(net3954));
 sky130_fd_sc_hd__buf_1 max_length3955 (.A(_09798_),
    .X(net3955));
 sky130_fd_sc_hd__buf_1 wire3956 (.A(net3961),
    .X(net3956));
 sky130_fd_sc_hd__clkbuf_1 wire3957 (.A(net3958),
    .X(net3957));
 sky130_fd_sc_hd__clkbuf_1 wire3958 (.A(net3959),
    .X(net3958));
 sky130_fd_sc_hd__buf_1 wire3959 (.A(net3960),
    .X(net3959));
 sky130_fd_sc_hd__buf_1 wire3960 (.A(net3961),
    .X(net3960));
 sky130_fd_sc_hd__buf_1 wire3961 (.A(net3962),
    .X(net3961));
 sky130_fd_sc_hd__clkbuf_1 wire3962 (.A(_09795_),
    .X(net3962));
 sky130_fd_sc_hd__buf_1 max_length3963 (.A(_09795_),
    .X(net3963));
 sky130_fd_sc_hd__buf_1 wire3964 (.A(net3965),
    .X(net3964));
 sky130_fd_sc_hd__clkbuf_1 wire3965 (.A(_09735_),
    .X(net3965));
 sky130_fd_sc_hd__buf_1 wire3966 (.A(net3967),
    .X(net3966));
 sky130_fd_sc_hd__buf_1 wire3967 (.A(net3968),
    .X(net3967));
 sky130_fd_sc_hd__clkbuf_1 wire3968 (.A(_09735_),
    .X(net3968));
 sky130_fd_sc_hd__buf_1 wire3969 (.A(_09703_),
    .X(net3969));
 sky130_fd_sc_hd__buf_1 wire3970 (.A(net3971),
    .X(net3970));
 sky130_fd_sc_hd__clkbuf_1 max_length3971 (.A(_09696_),
    .X(net3971));
 sky130_fd_sc_hd__clkbuf_1 wire3972 (.A(_09689_),
    .X(net3972));
 sky130_fd_sc_hd__clkbuf_1 wire3973 (.A(_09685_),
    .X(net3973));
 sky130_fd_sc_hd__clkbuf_1 wire3974 (.A(net3975),
    .X(net3974));
 sky130_fd_sc_hd__clkbuf_1 wire3975 (.A(_09682_),
    .X(net3975));
 sky130_fd_sc_hd__buf_1 wire3976 (.A(_09679_),
    .X(net3976));
 sky130_fd_sc_hd__clkbuf_2 wire3977 (.A(net3978),
    .X(net3977));
 sky130_fd_sc_hd__clkbuf_1 wire3978 (.A(net3979),
    .X(net3978));
 sky130_fd_sc_hd__clkbuf_1 wire3979 (.A(net3980),
    .X(net3979));
 sky130_fd_sc_hd__clkbuf_1 wire3980 (.A(net3984),
    .X(net3980));
 sky130_fd_sc_hd__buf_1 wire3981 (.A(net3982),
    .X(net3981));
 sky130_fd_sc_hd__buf_1 wire3982 (.A(net3983),
    .X(net3982));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire3983 (.A(net3984),
    .X(net3983));
 sky130_fd_sc_hd__clkbuf_1 wire3984 (.A(_09663_),
    .X(net3984));
 sky130_fd_sc_hd__clkbuf_1 wire3985 (.A(_09661_),
    .X(net3985));
 sky130_fd_sc_hd__buf_1 wire3986 (.A(net3987),
    .X(net3986));
 sky130_fd_sc_hd__buf_1 wire3987 (.A(_09660_),
    .X(net3987));
 sky130_fd_sc_hd__buf_1 wire3988 (.A(net3989),
    .X(net3988));
 sky130_fd_sc_hd__buf_1 wire3989 (.A(_09660_),
    .X(net3989));
 sky130_fd_sc_hd__buf_1 wire3990 (.A(net3991),
    .X(net3990));
 sky130_fd_sc_hd__clkbuf_1 max_length3991 (.A(_09641_),
    .X(net3991));
 sky130_fd_sc_hd__clkbuf_1 wire3992 (.A(_09636_),
    .X(net3992));
 sky130_fd_sc_hd__buf_1 wire3993 (.A(_09634_),
    .X(net3993));
 sky130_fd_sc_hd__buf_1 wire3994 (.A(net3995),
    .X(net3994));
 sky130_fd_sc_hd__buf_1 wire3995 (.A(_09624_),
    .X(net3995));
 sky130_fd_sc_hd__buf_1 wire3996 (.A(_09617_),
    .X(net3996));
 sky130_fd_sc_hd__buf_2 wire3997 (.A(_09606_),
    .X(net3997));
 sky130_fd_sc_hd__buf_1 wire3998 (.A(_09604_),
    .X(net3998));
 sky130_fd_sc_hd__clkbuf_1 wire3999 (.A(net4000),
    .X(net3999));
 sky130_fd_sc_hd__buf_1 wire4000 (.A(_09581_),
    .X(net4000));
 sky130_fd_sc_hd__buf_1 max_length4001 (.A(_09581_),
    .X(net4001));
 sky130_fd_sc_hd__buf_1 wire4002 (.A(net4003),
    .X(net4002));
 sky130_fd_sc_hd__buf_1 max_length4003 (.A(_09451_),
    .X(net4003));
 sky130_fd_sc_hd__buf_1 wire4004 (.A(_09426_),
    .X(net4004));
 sky130_fd_sc_hd__clkbuf_1 wire4005 (.A(_09376_),
    .X(net4005));
 sky130_fd_sc_hd__clkbuf_2 wire4006 (.A(net4007),
    .X(net4006));
 sky130_fd_sc_hd__buf_1 wire4007 (.A(_09376_),
    .X(net4007));
 sky130_fd_sc_hd__clkbuf_1 wire4008 (.A(_09358_),
    .X(net4008));
 sky130_fd_sc_hd__buf_1 wire4009 (.A(net4010),
    .X(net4009));
 sky130_fd_sc_hd__clkbuf_1 wire4010 (.A(net4011),
    .X(net4010));
 sky130_fd_sc_hd__buf_1 max_length4011 (.A(_09358_),
    .X(net4011));
 sky130_fd_sc_hd__buf_1 wire4012 (.A(net4013),
    .X(net4012));
 sky130_fd_sc_hd__buf_1 wire4013 (.A(_09339_),
    .X(net4013));
 sky130_fd_sc_hd__buf_1 wire4014 (.A(_09291_),
    .X(net4014));
 sky130_fd_sc_hd__buf_1 wire4015 (.A(_09257_),
    .X(net4015));
 sky130_fd_sc_hd__buf_1 max_length4016 (.A(_09257_),
    .X(net4016));
 sky130_fd_sc_hd__buf_1 wire4017 (.A(net4018),
    .X(net4017));
 sky130_fd_sc_hd__buf_1 max_length4018 (.A(net4019),
    .X(net4018));
 sky130_fd_sc_hd__buf_1 wire4019 (.A(_09243_),
    .X(net4019));
 sky130_fd_sc_hd__buf_1 wire4020 (.A(net4021),
    .X(net4020));
 sky130_fd_sc_hd__buf_1 wire4021 (.A(_09230_),
    .X(net4021));
 sky130_fd_sc_hd__buf_1 wire4022 (.A(net4023),
    .X(net4022));
 sky130_fd_sc_hd__buf_1 wire4023 (.A(_09230_),
    .X(net4023));
 sky130_fd_sc_hd__clkbuf_1 wire4024 (.A(net4025),
    .X(net4024));
 sky130_fd_sc_hd__buf_1 wire4025 (.A(net4026),
    .X(net4025));
 sky130_fd_sc_hd__buf_1 wire4026 (.A(_09223_),
    .X(net4026));
 sky130_fd_sc_hd__buf_1 wire4027 (.A(_09223_),
    .X(net4027));
 sky130_fd_sc_hd__clkbuf_1 wire4028 (.A(net4029),
    .X(net4028));
 sky130_fd_sc_hd__clkbuf_1 wire4029 (.A(net4030),
    .X(net4029));
 sky130_fd_sc_hd__clkbuf_2 wire4030 (.A(_09215_),
    .X(net4030));
 sky130_fd_sc_hd__buf_1 wire4031 (.A(_09215_),
    .X(net4031));
 sky130_fd_sc_hd__buf_1 wire4032 (.A(net4033),
    .X(net4032));
 sky130_fd_sc_hd__buf_1 wire4033 (.A(net4034),
    .X(net4033));
 sky130_fd_sc_hd__clkbuf_1 wire4034 (.A(_09196_),
    .X(net4034));
 sky130_fd_sc_hd__buf_1 max_length4035 (.A(_09196_),
    .X(net4035));
 sky130_fd_sc_hd__buf_1 wire4036 (.A(_09156_),
    .X(net4036));
 sky130_fd_sc_hd__buf_1 wire4037 (.A(_09054_),
    .X(net4037));
 sky130_fd_sc_hd__buf_1 wire4038 (.A(_09054_),
    .X(net4038));
 sky130_fd_sc_hd__buf_1 wire4039 (.A(net4042),
    .X(net4039));
 sky130_fd_sc_hd__buf_1 max_length4040 (.A(net4042),
    .X(net4040));
 sky130_fd_sc_hd__buf_1 max_length4041 (.A(_09032_),
    .X(net4041));
 sky130_fd_sc_hd__buf_1 max_length4042 (.A(_09032_),
    .X(net4042));
 sky130_fd_sc_hd__buf_1 wire4043 (.A(net4044),
    .X(net4043));
 sky130_fd_sc_hd__buf_1 wire4044 (.A(_08966_),
    .X(net4044));
 sky130_fd_sc_hd__buf_1 max_length4045 (.A(net4046),
    .X(net4045));
 sky130_fd_sc_hd__clkbuf_2 wire4046 (.A(_08954_),
    .X(net4046));
 sky130_fd_sc_hd__clkbuf_1 max_length4047 (.A(net4048),
    .X(net4047));
 sky130_fd_sc_hd__buf_1 wire4048 (.A(_08954_),
    .X(net4048));
 sky130_fd_sc_hd__clkbuf_1 wire4049 (.A(_08949_),
    .X(net4049));
 sky130_fd_sc_hd__clkbuf_1 wire4050 (.A(net4051),
    .X(net4050));
 sky130_fd_sc_hd__clkbuf_1 max_length4051 (.A(_08945_),
    .X(net4051));
 sky130_fd_sc_hd__clkbuf_1 max_length4052 (.A(_08943_),
    .X(net4052));
 sky130_fd_sc_hd__clkbuf_1 wire4053 (.A(_08932_),
    .X(net4053));
 sky130_fd_sc_hd__buf_1 wire4054 (.A(_08900_),
    .X(net4054));
 sky130_fd_sc_hd__buf_1 wire4055 (.A(_08896_),
    .X(net4055));
 sky130_fd_sc_hd__clkbuf_1 wire4056 (.A(_08848_),
    .X(net4056));
 sky130_fd_sc_hd__buf_1 wire4057 (.A(net4058),
    .X(net4057));
 sky130_fd_sc_hd__buf_1 max_length4058 (.A(_08834_),
    .X(net4058));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4059 (.A(_08832_),
    .X(net4059));
 sky130_fd_sc_hd__buf_1 wire4060 (.A(_08832_),
    .X(net4060));
 sky130_fd_sc_hd__clkbuf_1 wire4061 (.A(_08830_),
    .X(net4061));
 sky130_fd_sc_hd__clkbuf_2 wire4062 (.A(_08824_),
    .X(net4062));
 sky130_fd_sc_hd__buf_1 wire4063 (.A(net4064),
    .X(net4063));
 sky130_fd_sc_hd__clkbuf_1 wire4064 (.A(net4065),
    .X(net4064));
 sky130_fd_sc_hd__clkbuf_1 wire4065 (.A(net4066),
    .X(net4065));
 sky130_fd_sc_hd__clkbuf_1 wire4066 (.A(_08659_),
    .X(net4066));
 sky130_fd_sc_hd__buf_1 wire4067 (.A(_08644_),
    .X(net4067));
 sky130_fd_sc_hd__buf_1 max_length4068 (.A(net4069),
    .X(net4068));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4069 (.A(net4070),
    .X(net4069));
 sky130_fd_sc_hd__clkbuf_1 wire4070 (.A(_07683_),
    .X(net4070));
 sky130_fd_sc_hd__buf_1 wire4071 (.A(net4072),
    .X(net4071));
 sky130_fd_sc_hd__buf_1 wire4072 (.A(net4073),
    .X(net4072));
 sky130_fd_sc_hd__clkbuf_1 wire4073 (.A(_07682_),
    .X(net4073));
 sky130_fd_sc_hd__buf_1 wire4074 (.A(_07602_),
    .X(net4074));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4075 (.A(net4076),
    .X(net4075));
 sky130_fd_sc_hd__buf_1 wire4076 (.A(_07601_),
    .X(net4076));
 sky130_fd_sc_hd__buf_1 wire4077 (.A(net4078),
    .X(net4077));
 sky130_fd_sc_hd__clkbuf_1 wire4078 (.A(_07573_),
    .X(net4078));
 sky130_fd_sc_hd__buf_1 wire4079 (.A(net4080),
    .X(net4079));
 sky130_fd_sc_hd__clkbuf_1 wire4080 (.A(_07572_),
    .X(net4080));
 sky130_fd_sc_hd__buf_1 wire4081 (.A(net4082),
    .X(net4081));
 sky130_fd_sc_hd__clkbuf_1 wire4082 (.A(_07515_),
    .X(net4082));
 sky130_fd_sc_hd__buf_1 wire4083 (.A(net4084),
    .X(net4083));
 sky130_fd_sc_hd__clkbuf_1 wire4084 (.A(net4085),
    .X(net4084));
 sky130_fd_sc_hd__clkbuf_1 wire4085 (.A(_07514_),
    .X(net4085));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4086 (.A(_07484_),
    .X(net4086));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4087 (.A(net4088),
    .X(net4087));
 sky130_fd_sc_hd__clkbuf_1 wire4088 (.A(_07483_),
    .X(net4088));
 sky130_fd_sc_hd__buf_1 wire4089 (.A(net4090),
    .X(net4089));
 sky130_fd_sc_hd__clkbuf_1 wire4090 (.A(net4091),
    .X(net4090));
 sky130_fd_sc_hd__clkbuf_1 wire4091 (.A(_07370_),
    .X(net4091));
 sky130_fd_sc_hd__buf_1 wire4092 (.A(net4093),
    .X(net4092));
 sky130_fd_sc_hd__clkbuf_1 wire4093 (.A(_07369_),
    .X(net4093));
 sky130_fd_sc_hd__buf_1 wire4094 (.A(_07352_),
    .X(net4094));
 sky130_fd_sc_hd__buf_1 wire4095 (.A(_07351_),
    .X(net4095));
 sky130_fd_sc_hd__clkbuf_2 wire4096 (.A(net4097),
    .X(net4096));
 sky130_fd_sc_hd__clkbuf_1 wire4097 (.A(_07144_),
    .X(net4097));
 sky130_fd_sc_hd__buf_1 wire4098 (.A(net4099),
    .X(net4098));
 sky130_fd_sc_hd__buf_1 wire4099 (.A(net4100),
    .X(net4099));
 sky130_fd_sc_hd__clkbuf_1 wire4100 (.A(_07143_),
    .X(net4100));
 sky130_fd_sc_hd__clkbuf_2 wire4101 (.A(net4102),
    .X(net4101));
 sky130_fd_sc_hd__clkbuf_1 wire4102 (.A(net4103),
    .X(net4102));
 sky130_fd_sc_hd__clkbuf_1 wire4103 (.A(net4104),
    .X(net4103));
 sky130_fd_sc_hd__clkbuf_1 wire4104 (.A(_07132_),
    .X(net4104));
 sky130_fd_sc_hd__buf_1 wire4105 (.A(net4106),
    .X(net4105));
 sky130_fd_sc_hd__clkbuf_1 wire4106 (.A(net4107),
    .X(net4106));
 sky130_fd_sc_hd__clkbuf_1 wire4107 (.A(_07131_),
    .X(net4107));
 sky130_fd_sc_hd__buf_1 wire4108 (.A(net4109),
    .X(net4108));
 sky130_fd_sc_hd__clkbuf_1 wire4109 (.A(net4110),
    .X(net4109));
 sky130_fd_sc_hd__clkbuf_1 wire4110 (.A(_07127_),
    .X(net4110));
 sky130_fd_sc_hd__buf_1 wire4111 (.A(net4112),
    .X(net4111));
 sky130_fd_sc_hd__clkbuf_1 wire4112 (.A(net4113),
    .X(net4112));
 sky130_fd_sc_hd__clkbuf_1 wire4113 (.A(_07126_),
    .X(net4113));
 sky130_fd_sc_hd__clkbuf_1 max_length4114 (.A(net4115),
    .X(net4114));
 sky130_fd_sc_hd__buf_1 wire4115 (.A(net4117),
    .X(net4115));
 sky130_fd_sc_hd__buf_1 wire4116 (.A(net4117),
    .X(net4116));
 sky130_fd_sc_hd__buf_1 wire4117 (.A(net4118),
    .X(net4117));
 sky130_fd_sc_hd__buf_1 wire4118 (.A(_07089_),
    .X(net4118));
 sky130_fd_sc_hd__clkbuf_1 max_length4119 (.A(net4120),
    .X(net4119));
 sky130_fd_sc_hd__buf_1 wire4120 (.A(net4122),
    .X(net4120));
 sky130_fd_sc_hd__buf_1 wire4121 (.A(net4122),
    .X(net4121));
 sky130_fd_sc_hd__buf_1 wire4122 (.A(net4123),
    .X(net4122));
 sky130_fd_sc_hd__buf_1 wire4123 (.A(_07088_),
    .X(net4123));
 sky130_fd_sc_hd__buf_1 wire4124 (.A(net4125),
    .X(net4124));
 sky130_fd_sc_hd__buf_1 wire4125 (.A(_07037_),
    .X(net4125));
 sky130_fd_sc_hd__buf_1 wire4126 (.A(net4127),
    .X(net4126));
 sky130_fd_sc_hd__buf_1 wire4127 (.A(_07036_),
    .X(net4127));
 sky130_fd_sc_hd__clkbuf_1 wire4128 (.A(net4129),
    .X(net4128));
 sky130_fd_sc_hd__buf_1 wire4129 (.A(net4130),
    .X(net4129));
 sky130_fd_sc_hd__buf_1 wire4130 (.A(net4131),
    .X(net4130));
 sky130_fd_sc_hd__buf_1 wire4131 (.A(net4132),
    .X(net4131));
 sky130_fd_sc_hd__buf_1 wire4132 (.A(net4133),
    .X(net4132));
 sky130_fd_sc_hd__clkbuf_1 wire4133 (.A(net4134),
    .X(net4133));
 sky130_fd_sc_hd__clkbuf_1 wire4134 (.A(_07030_),
    .X(net4134));
 sky130_fd_sc_hd__clkbuf_1 wire4135 (.A(net4136),
    .X(net4135));
 sky130_fd_sc_hd__buf_1 wire4136 (.A(net4137),
    .X(net4136));
 sky130_fd_sc_hd__buf_1 wire4137 (.A(net4138),
    .X(net4137));
 sky130_fd_sc_hd__buf_1 wire4138 (.A(_07029_),
    .X(net4138));
 sky130_fd_sc_hd__buf_1 wire4139 (.A(_07025_),
    .X(net4139));
 sky130_fd_sc_hd__clkbuf_2 wire4140 (.A(net4141),
    .X(net4140));
 sky130_fd_sc_hd__clkbuf_1 wire4141 (.A(net4142),
    .X(net4141));
 sky130_fd_sc_hd__buf_1 wire4142 (.A(_07023_),
    .X(net4142));
 sky130_fd_sc_hd__clkbuf_2 wire4143 (.A(net4144),
    .X(net4143));
 sky130_fd_sc_hd__clkbuf_1 wire4144 (.A(net4145),
    .X(net4144));
 sky130_fd_sc_hd__clkbuf_1 wire4145 (.A(_07022_),
    .X(net4145));
 sky130_fd_sc_hd__buf_1 wire4146 (.A(net4147),
    .X(net4146));
 sky130_fd_sc_hd__clkbuf_1 wire4147 (.A(_07020_),
    .X(net4147));
 sky130_fd_sc_hd__buf_1 wire4148 (.A(net4149),
    .X(net4148));
 sky130_fd_sc_hd__buf_1 wire4149 (.A(net4150),
    .X(net4149));
 sky130_fd_sc_hd__clkbuf_1 wire4150 (.A(net4151),
    .X(net4150));
 sky130_fd_sc_hd__buf_1 wire4151 (.A(net4152),
    .X(net4151));
 sky130_fd_sc_hd__clkbuf_1 wire4152 (.A(_07014_),
    .X(net4152));
 sky130_fd_sc_hd__buf_1 wire4153 (.A(net4154),
    .X(net4153));
 sky130_fd_sc_hd__buf_1 wire4154 (.A(net4155),
    .X(net4154));
 sky130_fd_sc_hd__clkbuf_1 wire4155 (.A(_07013_),
    .X(net4155));
 sky130_fd_sc_hd__buf_1 wire4156 (.A(net4157),
    .X(net4156));
 sky130_fd_sc_hd__buf_1 wire4157 (.A(net4158),
    .X(net4157));
 sky130_fd_sc_hd__buf_1 wire4158 (.A(net4159),
    .X(net4158));
 sky130_fd_sc_hd__buf_1 wire4159 (.A(_07010_),
    .X(net4159));
 sky130_fd_sc_hd__buf_1 wire4160 (.A(net4161),
    .X(net4160));
 sky130_fd_sc_hd__buf_1 wire4161 (.A(net4162),
    .X(net4161));
 sky130_fd_sc_hd__buf_1 wire4162 (.A(net4163),
    .X(net4162));
 sky130_fd_sc_hd__buf_1 wire4163 (.A(_07009_),
    .X(net4163));
 sky130_fd_sc_hd__buf_1 wire4164 (.A(net4165),
    .X(net4164));
 sky130_fd_sc_hd__buf_1 wire4165 (.A(net4166),
    .X(net4165));
 sky130_fd_sc_hd__buf_1 wire4166 (.A(net4167),
    .X(net4166));
 sky130_fd_sc_hd__buf_1 wire4167 (.A(net4168),
    .X(net4167));
 sky130_fd_sc_hd__clkbuf_1 wire4168 (.A(_07003_),
    .X(net4168));
 sky130_fd_sc_hd__buf_1 wire4169 (.A(net4170),
    .X(net4169));
 sky130_fd_sc_hd__buf_1 wire4170 (.A(net4172),
    .X(net4170));
 sky130_fd_sc_hd__buf_1 max_length4171 (.A(net4172),
    .X(net4171));
 sky130_fd_sc_hd__buf_1 wire4172 (.A(_07002_),
    .X(net4172));
 sky130_fd_sc_hd__buf_1 wire4173 (.A(net4174),
    .X(net4173));
 sky130_fd_sc_hd__buf_1 wire4174 (.A(_07000_),
    .X(net4174));
 sky130_fd_sc_hd__buf_1 wire4175 (.A(net4176),
    .X(net4175));
 sky130_fd_sc_hd__buf_1 wire4176 (.A(net4177),
    .X(net4176));
 sky130_fd_sc_hd__clkbuf_1 wire4177 (.A(_06999_),
    .X(net4177));
 sky130_fd_sc_hd__buf_1 wire4178 (.A(_06997_),
    .X(net4178));
 sky130_fd_sc_hd__buf_1 wire4179 (.A(net4180),
    .X(net4179));
 sky130_fd_sc_hd__buf_1 wire4180 (.A(_06995_),
    .X(net4180));
 sky130_fd_sc_hd__buf_1 wire4181 (.A(net4182),
    .X(net4181));
 sky130_fd_sc_hd__buf_1 wire4182 (.A(net4183),
    .X(net4182));
 sky130_fd_sc_hd__clkbuf_1 wire4183 (.A(_06994_),
    .X(net4183));
 sky130_fd_sc_hd__buf_1 max_length4184 (.A(net4185),
    .X(net4184));
 sky130_fd_sc_hd__buf_1 wire4185 (.A(net4187),
    .X(net4185));
 sky130_fd_sc_hd__buf_1 wire4186 (.A(net4187),
    .X(net4186));
 sky130_fd_sc_hd__buf_1 wire4187 (.A(net4188),
    .X(net4187));
 sky130_fd_sc_hd__clkbuf_1 wire4188 (.A(net4189),
    .X(net4188));
 sky130_fd_sc_hd__clkbuf_1 wire4189 (.A(_06993_),
    .X(net4189));
 sky130_fd_sc_hd__buf_1 max_length4190 (.A(net4191),
    .X(net4190));
 sky130_fd_sc_hd__buf_1 wire4191 (.A(net4192),
    .X(net4191));
 sky130_fd_sc_hd__buf_1 wire4192 (.A(_06992_),
    .X(net4192));
 sky130_fd_sc_hd__buf_1 max_length4193 (.A(net4194),
    .X(net4193));
 sky130_fd_sc_hd__buf_1 wire4194 (.A(_06983_),
    .X(net4194));
 sky130_fd_sc_hd__buf_1 max_length4195 (.A(net4196),
    .X(net4195));
 sky130_fd_sc_hd__buf_1 wire4196 (.A(_06982_),
    .X(net4196));
 sky130_fd_sc_hd__buf_1 wire4197 (.A(_06977_),
    .X(net4197));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4198 (.A(net4199),
    .X(net4198));
 sky130_fd_sc_hd__buf_1 wire4199 (.A(net4200),
    .X(net4199));
 sky130_fd_sc_hd__clkbuf_1 wire4200 (.A(_06976_),
    .X(net4200));
 sky130_fd_sc_hd__buf_1 wire4201 (.A(net4203),
    .X(net4201));
 sky130_fd_sc_hd__buf_1 max_length4202 (.A(net4203),
    .X(net4202));
 sky130_fd_sc_hd__buf_1 wire4203 (.A(net4204),
    .X(net4203));
 sky130_fd_sc_hd__buf_1 wire4204 (.A(_06975_),
    .X(net4204));
 sky130_fd_sc_hd__buf_1 max_length4205 (.A(net4206),
    .X(net4205));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4206 (.A(net4207),
    .X(net4206));
 sky130_fd_sc_hd__buf_1 wire4207 (.A(_06974_),
    .X(net4207));
 sky130_fd_sc_hd__clkbuf_2 wire4208 (.A(net4209),
    .X(net4208));
 sky130_fd_sc_hd__clkbuf_1 wire4209 (.A(_06972_),
    .X(net4209));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4210 (.A(_06971_),
    .X(net4210));
 sky130_fd_sc_hd__buf_1 wire4211 (.A(net4212),
    .X(net4211));
 sky130_fd_sc_hd__buf_1 wire4212 (.A(_06970_),
    .X(net4212));
 sky130_fd_sc_hd__buf_1 wire4213 (.A(_06969_),
    .X(net4213));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4214 (.A(net4215),
    .X(net4214));
 sky130_fd_sc_hd__clkbuf_1 wire4215 (.A(_06966_),
    .X(net4215));
 sky130_fd_sc_hd__clkbuf_2 wire4216 (.A(net4217),
    .X(net4216));
 sky130_fd_sc_hd__clkbuf_1 wire4217 (.A(net4218),
    .X(net4217));
 sky130_fd_sc_hd__clkbuf_1 wire4218 (.A(_06965_),
    .X(net4218));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4219 (.A(net4220),
    .X(net4219));
 sky130_fd_sc_hd__buf_1 wire4220 (.A(_06963_),
    .X(net4220));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4221 (.A(net4222),
    .X(net4221));
 sky130_fd_sc_hd__buf_1 wire4222 (.A(_06962_),
    .X(net4222));
 sky130_fd_sc_hd__clkbuf_1 wire4223 (.A(_06826_),
    .X(net4223));
 sky130_fd_sc_hd__clkbuf_1 max_length4224 (.A(_06826_),
    .X(net4224));
 sky130_fd_sc_hd__clkbuf_1 wire4225 (.A(_06708_),
    .X(net4225));
 sky130_fd_sc_hd__buf_1 wire4226 (.A(net4227),
    .X(net4226));
 sky130_fd_sc_hd__clkbuf_1 wire4227 (.A(net4228),
    .X(net4227));
 sky130_fd_sc_hd__clkbuf_1 wire4228 (.A(net4229),
    .X(net4228));
 sky130_fd_sc_hd__clkbuf_1 wire4229 (.A(net4230),
    .X(net4229));
 sky130_fd_sc_hd__clkbuf_1 wire4230 (.A(net4231),
    .X(net4230));
 sky130_fd_sc_hd__clkbuf_1 max_length4231 (.A(_06708_),
    .X(net4231));
 sky130_fd_sc_hd__buf_1 wire4232 (.A(_06532_),
    .X(net4232));
 sky130_fd_sc_hd__buf_1 wire4233 (.A(net4234),
    .X(net4233));
 sky130_fd_sc_hd__clkbuf_1 wire4234 (.A(_06526_),
    .X(net4234));
 sky130_fd_sc_hd__buf_1 max_length4235 (.A(_06512_),
    .X(net4235));
 sky130_fd_sc_hd__clkbuf_1 wire4236 (.A(_06512_),
    .X(net4236));
 sky130_fd_sc_hd__clkbuf_1 max_length4237 (.A(_06503_),
    .X(net4237));
 sky130_fd_sc_hd__clkbuf_1 max_length4238 (.A(_06503_),
    .X(net4238));
 sky130_fd_sc_hd__clkbuf_1 wire4239 (.A(net4240),
    .X(net4239));
 sky130_fd_sc_hd__clkbuf_1 max_length4240 (.A(net4241),
    .X(net4240));
 sky130_fd_sc_hd__buf_1 wire4241 (.A(net4242),
    .X(net4241));
 sky130_fd_sc_hd__clkbuf_1 wire4242 (.A(net4243),
    .X(net4242));
 sky130_fd_sc_hd__clkbuf_1 wire4243 (.A(net4244),
    .X(net4243));
 sky130_fd_sc_hd__clkbuf_1 wire4244 (.A(net4246),
    .X(net4244));
 sky130_fd_sc_hd__buf_1 wire4245 (.A(net4246),
    .X(net4245));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4246 (.A(net4247),
    .X(net4246));
 sky130_fd_sc_hd__clkbuf_1 max_length4247 (.A(_06499_),
    .X(net4247));
 sky130_fd_sc_hd__buf_1 wire4248 (.A(net4249),
    .X(net4248));
 sky130_fd_sc_hd__buf_1 wire4249 (.A(net4250),
    .X(net4249));
 sky130_fd_sc_hd__buf_1 max_length4250 (.A(_05972_),
    .X(net4250));
 sky130_fd_sc_hd__clkbuf_1 wire4251 (.A(net4252),
    .X(net4251));
 sky130_fd_sc_hd__clkbuf_1 wire4252 (.A(net4253),
    .X(net4252));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4253 (.A(_05776_),
    .X(net4253));
 sky130_fd_sc_hd__buf_1 wire4254 (.A(net4255),
    .X(net4254));
 sky130_fd_sc_hd__buf_1 wire4255 (.A(_05347_),
    .X(net4255));
 sky130_fd_sc_hd__buf_1 wire4256 (.A(net4257),
    .X(net4256));
 sky130_fd_sc_hd__clkbuf_1 wire4257 (.A(net4258),
    .X(net4257));
 sky130_fd_sc_hd__clkbuf_1 max_length4258 (.A(_05127_),
    .X(net4258));
 sky130_fd_sc_hd__buf_1 wire4259 (.A(net4261),
    .X(net4259));
 sky130_fd_sc_hd__buf_1 wire4260 (.A(net4261),
    .X(net4260));
 sky130_fd_sc_hd__buf_1 wire4261 (.A(net4262),
    .X(net4261));
 sky130_fd_sc_hd__clkbuf_1 wire4262 (.A(net4263),
    .X(net4262));
 sky130_fd_sc_hd__clkbuf_1 wire4263 (.A(net4264),
    .X(net4263));
 sky130_fd_sc_hd__clkbuf_1 max_length4264 (.A(_04973_),
    .X(net4264));
 sky130_fd_sc_hd__buf_1 wire4265 (.A(_04928_),
    .X(net4265));
 sky130_fd_sc_hd__clkbuf_1 wire4266 (.A(net4267),
    .X(net4266));
 sky130_fd_sc_hd__clkbuf_1 max_length4267 (.A(_04928_),
    .X(net4267));
 sky130_fd_sc_hd__clkbuf_1 wire4268 (.A(_04911_),
    .X(net4268));
 sky130_fd_sc_hd__clkbuf_1 wire4269 (.A(net4270),
    .X(net4269));
 sky130_fd_sc_hd__clkbuf_1 wire4270 (.A(net4271),
    .X(net4270));
 sky130_fd_sc_hd__clkbuf_1 wire4271 (.A(_04911_),
    .X(net4271));
 sky130_fd_sc_hd__buf_1 wire4272 (.A(net4273),
    .X(net4272));
 sky130_fd_sc_hd__clkbuf_1 wire4273 (.A(net4274),
    .X(net4273));
 sky130_fd_sc_hd__clkbuf_1 wire4274 (.A(net4276),
    .X(net4274));
 sky130_fd_sc_hd__clkbuf_1 wire4275 (.A(_04898_),
    .X(net4275));
 sky130_fd_sc_hd__clkbuf_1 max_length4276 (.A(_04898_),
    .X(net4276));
 sky130_fd_sc_hd__buf_1 max_cap4277 (.A(_04896_),
    .X(net4277));
 sky130_fd_sc_hd__buf_1 wire4278 (.A(_04893_),
    .X(net4278));
 sky130_fd_sc_hd__clkbuf_1 wire4279 (.A(net4280),
    .X(net4279));
 sky130_fd_sc_hd__clkbuf_1 wire4280 (.A(net4281),
    .X(net4280));
 sky130_fd_sc_hd__buf_1 wire4281 (.A(net4286),
    .X(net4281));
 sky130_fd_sc_hd__clkbuf_1 wire4282 (.A(net4283),
    .X(net4282));
 sky130_fd_sc_hd__buf_1 wire4283 (.A(net4284),
    .X(net4283));
 sky130_fd_sc_hd__buf_1 wire4284 (.A(net4285),
    .X(net4284));
 sky130_fd_sc_hd__buf_1 wire4285 (.A(net4286),
    .X(net4285));
 sky130_fd_sc_hd__buf_1 wire4286 (.A(_04883_),
    .X(net4286));
 sky130_fd_sc_hd__clkbuf_2 wire4287 (.A(net4288),
    .X(net4287));
 sky130_fd_sc_hd__clkbuf_1 wire4288 (.A(net4289),
    .X(net4288));
 sky130_fd_sc_hd__buf_1 wire4289 (.A(net4290),
    .X(net4289));
 sky130_fd_sc_hd__clkbuf_1 max_length4290 (.A(net4291),
    .X(net4290));
 sky130_fd_sc_hd__buf_1 wire4291 (.A(net4292),
    .X(net4291));
 sky130_fd_sc_hd__buf_1 wire4292 (.A(_04876_),
    .X(net4292));
 sky130_fd_sc_hd__clkbuf_1 wire4293 (.A(net4294),
    .X(net4293));
 sky130_fd_sc_hd__clkbuf_1 wire4294 (.A(net4295),
    .X(net4294));
 sky130_fd_sc_hd__clkbuf_1 wire4295 (.A(net4296),
    .X(net4295));
 sky130_fd_sc_hd__clkbuf_1 wire4296 (.A(_04875_),
    .X(net4296));
 sky130_fd_sc_hd__buf_1 wire4297 (.A(_04872_),
    .X(net4297));
 sky130_fd_sc_hd__buf_1 wire4298 (.A(net4299),
    .X(net4298));
 sky130_fd_sc_hd__buf_1 wire4299 (.A(net4300),
    .X(net4299));
 sky130_fd_sc_hd__buf_1 wire4300 (.A(net4301),
    .X(net4300));
 sky130_fd_sc_hd__buf_1 wire4301 (.A(_04872_),
    .X(net4301));
 sky130_fd_sc_hd__buf_1 wire4302 (.A(net4303),
    .X(net4302));
 sky130_fd_sc_hd__buf_1 wire4303 (.A(net4304),
    .X(net4303));
 sky130_fd_sc_hd__clkbuf_1 wire4304 (.A(net4305),
    .X(net4304));
 sky130_fd_sc_hd__clkbuf_1 wire4305 (.A(net4306),
    .X(net4305));
 sky130_fd_sc_hd__clkbuf_1 wire4306 (.A(net4307),
    .X(net4306));
 sky130_fd_sc_hd__clkbuf_1 wire4307 (.A(net4309),
    .X(net4307));
 sky130_fd_sc_hd__clkbuf_1 wire4308 (.A(_04866_),
    .X(net4308));
 sky130_fd_sc_hd__clkbuf_1 max_length4309 (.A(_04866_),
    .X(net4309));
 sky130_fd_sc_hd__buf_1 wire4310 (.A(_04862_),
    .X(net4310));
 sky130_fd_sc_hd__clkbuf_1 wire4311 (.A(net4312),
    .X(net4311));
 sky130_fd_sc_hd__clkbuf_1 wire4312 (.A(_04861_),
    .X(net4312));
 sky130_fd_sc_hd__clkbuf_1 wire4313 (.A(_04861_),
    .X(net4313));
 sky130_fd_sc_hd__clkbuf_1 fanout4314 (.A(net4322),
    .X(net4314));
 sky130_fd_sc_hd__buf_1 wire4315 (.A(net4316),
    .X(net4315));
 sky130_fd_sc_hd__buf_1 wire4316 (.A(net4317),
    .X(net4316));
 sky130_fd_sc_hd__buf_1 max_length4317 (.A(net4314),
    .X(net4317));
 sky130_fd_sc_hd__buf_1 fanout4318 (.A(net4323),
    .X(net4318));
 sky130_fd_sc_hd__buf_1 wire4319 (.A(net4318),
    .X(net4319));
 sky130_fd_sc_hd__buf_1 wire4320 (.A(net4318),
    .X(net4320));
 sky130_fd_sc_hd__clkbuf_1 wire4321 (.A(net4322),
    .X(net4321));
 sky130_fd_sc_hd__buf_1 wire4322 (.A(net4323),
    .X(net4322));
 sky130_fd_sc_hd__buf_1 wire4323 (.A(\pid_d.state[5] ),
    .X(net4323));
 sky130_fd_sc_hd__buf_1 fanout4324 (.A(\pid_d.state[4] ),
    .X(net4324));
 sky130_fd_sc_hd__buf_1 wire4325 (.A(net4326),
    .X(net4325));
 sky130_fd_sc_hd__buf_1 max_length4326 (.A(net4327),
    .X(net4326));
 sky130_fd_sc_hd__buf_1 wire4327 (.A(net4324),
    .X(net4327));
 sky130_fd_sc_hd__buf_1 wire4328 (.A(net4329),
    .X(net4328));
 sky130_fd_sc_hd__clkbuf_1 wire4329 (.A(net4330),
    .X(net4329));
 sky130_fd_sc_hd__clkbuf_1 wire4330 (.A(net4324),
    .X(net4330));
 sky130_fd_sc_hd__clkbuf_2 fanout4331 (.A(net4334),
    .X(net4331));
 sky130_fd_sc_hd__clkbuf_1 wire4332 (.A(net4333),
    .X(net4332));
 sky130_fd_sc_hd__buf_1 wire4333 (.A(net4331),
    .X(net4333));
 sky130_fd_sc_hd__clkbuf_1 fanout4334 (.A(net4340),
    .X(net4334));
 sky130_fd_sc_hd__buf_1 max_length4335 (.A(net4336),
    .X(net4335));
 sky130_fd_sc_hd__buf_1 wire4336 (.A(net4337),
    .X(net4336));
 sky130_fd_sc_hd__buf_1 wire4337 (.A(net4338),
    .X(net4337));
 sky130_fd_sc_hd__buf_1 wire4338 (.A(net4339),
    .X(net4338));
 sky130_fd_sc_hd__clkbuf_1 wire4339 (.A(net4334),
    .X(net4339));
 sky130_fd_sc_hd__clkbuf_1 wire4340 (.A(\pid_d.state[4] ),
    .X(net4340));
 sky130_fd_sc_hd__clkbuf_1 wire4341 (.A(net4342),
    .X(net4341));
 sky130_fd_sc_hd__clkbuf_1 wire4342 (.A(net4343),
    .X(net4342));
 sky130_fd_sc_hd__clkbuf_1 wire4343 (.A(net4344),
    .X(net4343));
 sky130_fd_sc_hd__clkbuf_1 wire4344 (.A(net4345),
    .X(net4344));
 sky130_fd_sc_hd__clkbuf_1 wire4345 (.A(net4346),
    .X(net4345));
 sky130_fd_sc_hd__buf_1 wire4346 (.A(net4351),
    .X(net4346));
 sky130_fd_sc_hd__clkbuf_1 wire4347 (.A(net4348),
    .X(net4347));
 sky130_fd_sc_hd__clkbuf_1 wire4348 (.A(net4349),
    .X(net4348));
 sky130_fd_sc_hd__clkbuf_1 wire4349 (.A(net4350),
    .X(net4349));
 sky130_fd_sc_hd__clkbuf_1 wire4350 (.A(net4351),
    .X(net4350));
 sky130_fd_sc_hd__buf_1 wire4351 (.A(\pid_d.state[3] ),
    .X(net4351));
 sky130_fd_sc_hd__buf_1 fanout4352 (.A(net4369),
    .X(net4352));
 sky130_fd_sc_hd__clkbuf_1 wire4353 (.A(net4352),
    .X(net4353));
 sky130_fd_sc_hd__buf_1 wire4354 (.A(net4355),
    .X(net4354));
 sky130_fd_sc_hd__clkbuf_1 wire4355 (.A(net4356),
    .X(net4355));
 sky130_fd_sc_hd__buf_1 wire4356 (.A(net4357),
    .X(net4356));
 sky130_fd_sc_hd__buf_1 wire4357 (.A(net4358),
    .X(net4357));
 sky130_fd_sc_hd__buf_1 wire4358 (.A(net4352),
    .X(net4358));
 sky130_fd_sc_hd__buf_1 fanout4359 (.A(net4371),
    .X(net4359));
 sky130_fd_sc_hd__buf_1 wire4360 (.A(net4359),
    .X(net4360));
 sky130_fd_sc_hd__clkbuf_1 fanout4361 (.A(net4368),
    .X(net4361));
 sky130_fd_sc_hd__buf_1 wire4362 (.A(net4363),
    .X(net4362));
 sky130_fd_sc_hd__buf_1 max_length4363 (.A(net4365),
    .X(net4363));
 sky130_fd_sc_hd__buf_1 max_length4364 (.A(net4365),
    .X(net4364));
 sky130_fd_sc_hd__buf_1 wire4365 (.A(net4366),
    .X(net4365));
 sky130_fd_sc_hd__buf_1 wire4366 (.A(net4361),
    .X(net4366));
 sky130_fd_sc_hd__buf_1 wire4367 (.A(net4361),
    .X(net4367));
 sky130_fd_sc_hd__buf_1 fanout4368 (.A(net4376),
    .X(net4368));
 sky130_fd_sc_hd__clkbuf_1 wire4369 (.A(net4375),
    .X(net4369));
 sky130_fd_sc_hd__buf_1 wire4370 (.A(net4372),
    .X(net4370));
 sky130_fd_sc_hd__clkbuf_1 wire4371 (.A(net4372),
    .X(net4371));
 sky130_fd_sc_hd__buf_1 wire4372 (.A(net4373),
    .X(net4372));
 sky130_fd_sc_hd__clkbuf_1 wire4373 (.A(net4374),
    .X(net4373));
 sky130_fd_sc_hd__clkbuf_1 wire4374 (.A(net4375),
    .X(net4374));
 sky130_fd_sc_hd__buf_1 wire4375 (.A(net4368),
    .X(net4375));
 sky130_fd_sc_hd__clkbuf_1 wire4376 (.A(net4377),
    .X(net4376));
 sky130_fd_sc_hd__clkbuf_1 wire4377 (.A(net4378),
    .X(net4377));
 sky130_fd_sc_hd__clkbuf_1 wire4378 (.A(\pid_d.state[2] ),
    .X(net4378));
 sky130_fd_sc_hd__buf_1 fanout4379 (.A(net4388),
    .X(net4379));
 sky130_fd_sc_hd__buf_1 wire4380 (.A(net4379),
    .X(net4380));
 sky130_fd_sc_hd__buf_1 wire4381 (.A(net4382),
    .X(net4381));
 sky130_fd_sc_hd__buf_1 wire4382 (.A(net4379),
    .X(net4382));
 sky130_fd_sc_hd__buf_1 fanout4383 (.A(net4386),
    .X(net4383));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4384 (.A(net4385),
    .X(net4384));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4385 (.A(net4383),
    .X(net4385));
 sky130_fd_sc_hd__clkbuf_1 wire4386 (.A(net4387),
    .X(net4386));
 sky130_fd_sc_hd__clkbuf_1 wire4387 (.A(net4388),
    .X(net4387));
 sky130_fd_sc_hd__buf_1 max_length4388 (.A(\pid_d.state[1] ),
    .X(net4388));
 sky130_fd_sc_hd__buf_1 wire4389 (.A(net4390),
    .X(net4389));
 sky130_fd_sc_hd__buf_1 wire4390 (.A(\pid_d.state[0] ),
    .X(net4390));
 sky130_fd_sc_hd__buf_1 wire4391 (.A(\pid_d.prev_int[12] ),
    .X(net4391));
 sky130_fd_sc_hd__buf_1 wire4392 (.A(\pid_d.prev_int[0] ),
    .X(net4392));
 sky130_fd_sc_hd__buf_1 wire4393 (.A(\pid_q.out[15] ),
    .X(net4393));
 sky130_fd_sc_hd__clkbuf_1 wire4394 (.A(net4395),
    .X(net4394));
 sky130_fd_sc_hd__clkbuf_1 wire4395 (.A(net4396),
    .X(net4395));
 sky130_fd_sc_hd__clkbuf_1 wire4396 (.A(\pid_q.out[15] ),
    .X(net4396));
 sky130_fd_sc_hd__clkbuf_1 wire4397 (.A(net4398),
    .X(net4397));
 sky130_fd_sc_hd__clkbuf_1 wire4398 (.A(net4399),
    .X(net4398));
 sky130_fd_sc_hd__clkbuf_1 wire4399 (.A(\pid_q.out[14] ),
    .X(net4399));
 sky130_fd_sc_hd__buf_1 max_length4400 (.A(\pid_q.out[14] ),
    .X(net4400));
 sky130_fd_sc_hd__clkbuf_2 wire4401 (.A(\pid_q.out[13] ),
    .X(net4401));
 sky130_fd_sc_hd__clkbuf_1 wire4402 (.A(net4403),
    .X(net4402));
 sky130_fd_sc_hd__clkbuf_1 wire4403 (.A(net4404),
    .X(net4403));
 sky130_fd_sc_hd__clkbuf_1 wire4404 (.A(net4405),
    .X(net4404));
 sky130_fd_sc_hd__clkbuf_1 wire4405 (.A(\pid_q.out[13] ),
    .X(net4405));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4406 (.A(\pid_q.out[12] ),
    .X(net4406));
 sky130_fd_sc_hd__clkbuf_1 wire4407 (.A(net4408),
    .X(net4407));
 sky130_fd_sc_hd__clkbuf_1 wire4408 (.A(net4409),
    .X(net4408));
 sky130_fd_sc_hd__clkbuf_1 wire4409 (.A(net4410),
    .X(net4409));
 sky130_fd_sc_hd__clkbuf_1 wire4410 (.A(net4411),
    .X(net4410));
 sky130_fd_sc_hd__clkbuf_1 wire4411 (.A(net4412),
    .X(net4411));
 sky130_fd_sc_hd__clkbuf_1 wire4412 (.A(\pid_q.out[12] ),
    .X(net4412));
 sky130_fd_sc_hd__clkbuf_1 wire4413 (.A(net4414),
    .X(net4413));
 sky130_fd_sc_hd__clkbuf_1 wire4414 (.A(net4415),
    .X(net4414));
 sky130_fd_sc_hd__clkbuf_1 wire4415 (.A(net4416),
    .X(net4415));
 sky130_fd_sc_hd__clkbuf_1 wire4416 (.A(net4417),
    .X(net4416));
 sky130_fd_sc_hd__clkbuf_1 wire4417 (.A(\pid_q.out[11] ),
    .X(net4417));
 sky130_fd_sc_hd__buf_1 max_length4418 (.A(\pid_q.out[11] ),
    .X(net4418));
 sky130_fd_sc_hd__clkbuf_1 wire4419 (.A(net4420),
    .X(net4419));
 sky130_fd_sc_hd__clkbuf_1 wire4420 (.A(net4421),
    .X(net4420));
 sky130_fd_sc_hd__clkbuf_1 wire4421 (.A(net4422),
    .X(net4421));
 sky130_fd_sc_hd__clkbuf_1 wire4422 (.A(net4423),
    .X(net4422));
 sky130_fd_sc_hd__clkbuf_1 wire4423 (.A(\pid_q.out[10] ),
    .X(net4423));
 sky130_fd_sc_hd__buf_1 max_length4424 (.A(\pid_q.out[10] ),
    .X(net4424));
 sky130_fd_sc_hd__clkbuf_1 wire4425 (.A(net4426),
    .X(net4425));
 sky130_fd_sc_hd__clkbuf_1 wire4426 (.A(net4427),
    .X(net4426));
 sky130_fd_sc_hd__clkbuf_1 wire4427 (.A(net4428),
    .X(net4427));
 sky130_fd_sc_hd__clkbuf_1 wire4428 (.A(net4429),
    .X(net4428));
 sky130_fd_sc_hd__clkbuf_1 wire4429 (.A(\pid_q.out[9] ),
    .X(net4429));
 sky130_fd_sc_hd__buf_1 max_length4430 (.A(\pid_q.out[9] ),
    .X(net4430));
 sky130_fd_sc_hd__clkbuf_1 wire4431 (.A(net4432),
    .X(net4431));
 sky130_fd_sc_hd__clkbuf_1 wire4432 (.A(net4433),
    .X(net4432));
 sky130_fd_sc_hd__clkbuf_1 wire4433 (.A(net4434),
    .X(net4433));
 sky130_fd_sc_hd__clkbuf_1 wire4434 (.A(net4435),
    .X(net4434));
 sky130_fd_sc_hd__clkbuf_1 max_length4435 (.A(\pid_q.out[8] ),
    .X(net4435));
 sky130_fd_sc_hd__clkbuf_1 wire4436 (.A(net4437),
    .X(net4436));
 sky130_fd_sc_hd__clkbuf_1 wire4437 (.A(net4438),
    .X(net4437));
 sky130_fd_sc_hd__clkbuf_1 wire4438 (.A(net4439),
    .X(net4438));
 sky130_fd_sc_hd__clkbuf_1 wire4439 (.A(net4440),
    .X(net4439));
 sky130_fd_sc_hd__clkbuf_1 wire4440 (.A(net4441),
    .X(net4440));
 sky130_fd_sc_hd__clkbuf_1 wire4441 (.A(net4442),
    .X(net4441));
 sky130_fd_sc_hd__clkbuf_1 wire4442 (.A(\pid_q.out[7] ),
    .X(net4442));
 sky130_fd_sc_hd__clkbuf_1 wire4443 (.A(net4444),
    .X(net4443));
 sky130_fd_sc_hd__clkbuf_1 wire4444 (.A(net4445),
    .X(net4444));
 sky130_fd_sc_hd__clkbuf_1 wire4445 (.A(net4446),
    .X(net4445));
 sky130_fd_sc_hd__clkbuf_1 wire4446 (.A(net4447),
    .X(net4446));
 sky130_fd_sc_hd__clkbuf_1 max_length4447 (.A(\pid_q.out[6] ),
    .X(net4447));
 sky130_fd_sc_hd__clkbuf_1 wire4448 (.A(net4449),
    .X(net4448));
 sky130_fd_sc_hd__clkbuf_1 wire4449 (.A(net4450),
    .X(net4449));
 sky130_fd_sc_hd__clkbuf_1 wire4450 (.A(net4451),
    .X(net4450));
 sky130_fd_sc_hd__clkbuf_1 max_length4451 (.A(\pid_q.out[5] ),
    .X(net4451));
 sky130_fd_sc_hd__clkbuf_1 wire4452 (.A(net4453),
    .X(net4452));
 sky130_fd_sc_hd__clkbuf_1 wire4453 (.A(net4454),
    .X(net4453));
 sky130_fd_sc_hd__clkbuf_1 wire4454 (.A(net4455),
    .X(net4454));
 sky130_fd_sc_hd__clkbuf_1 wire4455 (.A(net4456),
    .X(net4455));
 sky130_fd_sc_hd__clkbuf_1 wire4456 (.A(\pid_q.out[4] ),
    .X(net4456));
 sky130_fd_sc_hd__buf_1 max_length4457 (.A(\pid_q.out[4] ),
    .X(net4457));
 sky130_fd_sc_hd__clkbuf_1 wire4458 (.A(net4459),
    .X(net4458));
 sky130_fd_sc_hd__clkbuf_1 wire4459 (.A(net4460),
    .X(net4459));
 sky130_fd_sc_hd__clkbuf_1 wire4460 (.A(net4461),
    .X(net4460));
 sky130_fd_sc_hd__clkbuf_1 wire4461 (.A(\pid_q.out[3] ),
    .X(net4461));
 sky130_fd_sc_hd__buf_1 max_length4462 (.A(\pid_q.out[3] ),
    .X(net4462));
 sky130_fd_sc_hd__clkbuf_1 wire4463 (.A(net4464),
    .X(net4463));
 sky130_fd_sc_hd__clkbuf_1 wire4464 (.A(net4465),
    .X(net4464));
 sky130_fd_sc_hd__clkbuf_1 wire4465 (.A(\pid_q.out[2] ),
    .X(net4465));
 sky130_fd_sc_hd__buf_1 max_length4466 (.A(\pid_q.out[2] ),
    .X(net4466));
 sky130_fd_sc_hd__clkbuf_1 wire4467 (.A(net4468),
    .X(net4467));
 sky130_fd_sc_hd__clkbuf_1 wire4468 (.A(net4469),
    .X(net4468));
 sky130_fd_sc_hd__clkbuf_1 wire4469 (.A(net4470),
    .X(net4469));
 sky130_fd_sc_hd__clkbuf_1 max_length4470 (.A(\pid_q.out[1] ),
    .X(net4470));
 sky130_fd_sc_hd__clkbuf_1 wire4471 (.A(net4472),
    .X(net4471));
 sky130_fd_sc_hd__clkbuf_1 wire4472 (.A(net4473),
    .X(net4472));
 sky130_fd_sc_hd__clkbuf_1 wire4473 (.A(net4474),
    .X(net4473));
 sky130_fd_sc_hd__clkbuf_2 max_length4474 (.A(\pid_q.out[0] ),
    .X(net4474));
 sky130_fd_sc_hd__clkbuf_1 wire4475 (.A(\pid_q.kp[15] ),
    .X(net4475));
 sky130_fd_sc_hd__clkbuf_1 wire4476 (.A(net4477),
    .X(net4476));
 sky130_fd_sc_hd__clkbuf_1 max_length4477 (.A(\pid_q.kp[9] ),
    .X(net4477));
 sky130_fd_sc_hd__clkbuf_1 wire4478 (.A(\pid_q.kp[5] ),
    .X(net4478));
 sky130_fd_sc_hd__clkbuf_1 wire4479 (.A(net4480),
    .X(net4479));
 sky130_fd_sc_hd__clkbuf_1 wire4480 (.A(\pid_q.ki[9] ),
    .X(net4480));
 sky130_fd_sc_hd__clkbuf_1 wire4481 (.A(\pid_q.ki[5] ),
    .X(net4481));
 sky130_fd_sc_hd__buf_1 fanout4482 (.A(net4489),
    .X(net4482));
 sky130_fd_sc_hd__buf_1 wire4483 (.A(net4486),
    .X(net4483));
 sky130_fd_sc_hd__buf_1 wire4484 (.A(net4485),
    .X(net4484));
 sky130_fd_sc_hd__buf_1 wire4485 (.A(net4482),
    .X(net4485));
 sky130_fd_sc_hd__buf_1 max_length4486 (.A(net4482),
    .X(net4486));
 sky130_fd_sc_hd__buf_1 fanout4487 (.A(net4493),
    .X(net4487));
 sky130_fd_sc_hd__buf_1 wire4488 (.A(net4489),
    .X(net4488));
 sky130_fd_sc_hd__buf_1 wire4489 (.A(net4490),
    .X(net4489));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4490 (.A(net4487),
    .X(net4490));
 sky130_fd_sc_hd__buf_1 wire4491 (.A(net4487),
    .X(net4491));
 sky130_fd_sc_hd__clkbuf_1 fanout4492 (.A(\pid_q.mult0.a[15] ),
    .X(net4492));
 sky130_fd_sc_hd__buf_1 wire4493 (.A(net4494),
    .X(net4493));
 sky130_fd_sc_hd__clkbuf_1 max_length4494 (.A(net4495),
    .X(net4494));
 sky130_fd_sc_hd__buf_1 wire4495 (.A(net4496),
    .X(net4495));
 sky130_fd_sc_hd__buf_1 wire4496 (.A(net4497),
    .X(net4496));
 sky130_fd_sc_hd__clkbuf_1 wire4497 (.A(net4492),
    .X(net4497));
 sky130_fd_sc_hd__buf_1 fanout4498 (.A(net4509),
    .X(net4498));
 sky130_fd_sc_hd__buf_1 wire4499 (.A(net4500),
    .X(net4499));
 sky130_fd_sc_hd__buf_1 wire4500 (.A(net4501),
    .X(net4500));
 sky130_fd_sc_hd__buf_1 max_length4501 (.A(net4502),
    .X(net4501));
 sky130_fd_sc_hd__buf_1 wire4502 (.A(net4498),
    .X(net4502));
 sky130_fd_sc_hd__buf_1 fanout4503 (.A(net4509),
    .X(net4503));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4504 (.A(net4503),
    .X(net4504));
 sky130_fd_sc_hd__clkbuf_1 max_length4505 (.A(net4506),
    .X(net4505));
 sky130_fd_sc_hd__buf_1 max_length4506 (.A(net4503),
    .X(net4506));
 sky130_fd_sc_hd__clkbuf_1 fanout4507 (.A(\pid_q.mult0.a[14] ),
    .X(net4507));
 sky130_fd_sc_hd__clkbuf_1 wire4508 (.A(net4511),
    .X(net4508));
 sky130_fd_sc_hd__buf_1 wire4509 (.A(net4510),
    .X(net4509));
 sky130_fd_sc_hd__clkbuf_1 wire4510 (.A(net4511),
    .X(net4510));
 sky130_fd_sc_hd__buf_1 wire4511 (.A(net4512),
    .X(net4511));
 sky130_fd_sc_hd__buf_1 wire4512 (.A(net4513),
    .X(net4512));
 sky130_fd_sc_hd__buf_1 wire4513 (.A(net4507),
    .X(net4513));
 sky130_fd_sc_hd__clkbuf_2 fanout4514 (.A(net4524),
    .X(net4514));
 sky130_fd_sc_hd__clkbuf_2 max_length4515 (.A(net4516),
    .X(net4515));
 sky130_fd_sc_hd__buf_1 wire4516 (.A(net4514),
    .X(net4516));
 sky130_fd_sc_hd__clkbuf_1 fanout4517 (.A(net4528),
    .X(net4517));
 sky130_fd_sc_hd__clkbuf_1 wire4518 (.A(net4519),
    .X(net4518));
 sky130_fd_sc_hd__buf_1 wire4519 (.A(net4521),
    .X(net4519));
 sky130_fd_sc_hd__clkbuf_1 max_length4520 (.A(net4521),
    .X(net4520));
 sky130_fd_sc_hd__buf_1 wire4521 (.A(net4522),
    .X(net4521));
 sky130_fd_sc_hd__buf_1 wire4522 (.A(net4524),
    .X(net4522));
 sky130_fd_sc_hd__buf_1 wire4523 (.A(net4524),
    .X(net4523));
 sky130_fd_sc_hd__buf_1 wire4524 (.A(net4517),
    .X(net4524));
 sky130_fd_sc_hd__buf_1 fanout4525 (.A(\pid_q.mult0.a[13] ),
    .X(net4525));
 sky130_fd_sc_hd__clkbuf_1 wire4526 (.A(net4527),
    .X(net4526));
 sky130_fd_sc_hd__buf_1 wire4527 (.A(net4530),
    .X(net4527));
 sky130_fd_sc_hd__clkbuf_1 wire4528 (.A(net4529),
    .X(net4528));
 sky130_fd_sc_hd__clkbuf_1 wire4529 (.A(net4531),
    .X(net4529));
 sky130_fd_sc_hd__clkbuf_1 max_length4530 (.A(net4531),
    .X(net4530));
 sky130_fd_sc_hd__buf_1 wire4531 (.A(net4532),
    .X(net4531));
 sky130_fd_sc_hd__buf_1 wire4532 (.A(net4525),
    .X(net4532));
 sky130_fd_sc_hd__clkbuf_1 fanout4533 (.A(net4546),
    .X(net4533));
 sky130_fd_sc_hd__buf_1 wire4534 (.A(net4535),
    .X(net4534));
 sky130_fd_sc_hd__buf_1 wire4535 (.A(net4536),
    .X(net4535));
 sky130_fd_sc_hd__buf_1 wire4536 (.A(net4537),
    .X(net4536));
 sky130_fd_sc_hd__buf_1 wire4537 (.A(net4539),
    .X(net4537));
 sky130_fd_sc_hd__clkbuf_1 wire4538 (.A(net4539),
    .X(net4538));
 sky130_fd_sc_hd__buf_1 wire4539 (.A(net4533),
    .X(net4539));
 sky130_fd_sc_hd__buf_1 fanout4540 (.A(net4550),
    .X(net4540));
 sky130_fd_sc_hd__clkbuf_1 wire4541 (.A(net4542),
    .X(net4541));
 sky130_fd_sc_hd__buf_1 wire4542 (.A(net4543),
    .X(net4542));
 sky130_fd_sc_hd__buf_1 wire4543 (.A(net4548),
    .X(net4543));
 sky130_fd_sc_hd__clkbuf_1 max_length4544 (.A(net4545),
    .X(net4544));
 sky130_fd_sc_hd__buf_1 wire4545 (.A(net4546),
    .X(net4545));
 sky130_fd_sc_hd__buf_1 wire4546 (.A(net4547),
    .X(net4546));
 sky130_fd_sc_hd__clkbuf_1 wire4547 (.A(net4549),
    .X(net4547));
 sky130_fd_sc_hd__buf_1 max_length4548 (.A(net4549),
    .X(net4548));
 sky130_fd_sc_hd__buf_1 wire4549 (.A(net4540),
    .X(net4549));
 sky130_fd_sc_hd__buf_1 wire4550 (.A(\pid_q.mult0.a[12] ),
    .X(net4550));
 sky130_fd_sc_hd__clkbuf_1 fanout4551 (.A(net4565),
    .X(net4551));
 sky130_fd_sc_hd__clkbuf_1 wire4552 (.A(net4553),
    .X(net4552));
 sky130_fd_sc_hd__buf_1 wire4553 (.A(net4554),
    .X(net4553));
 sky130_fd_sc_hd__buf_1 wire4554 (.A(net4555),
    .X(net4554));
 sky130_fd_sc_hd__clkbuf_2 wire4555 (.A(net4551),
    .X(net4555));
 sky130_fd_sc_hd__buf_1 fanout4556 (.A(\pid_q.mult0.a[11] ),
    .X(net4556));
 sky130_fd_sc_hd__clkbuf_1 wire4557 (.A(net4558),
    .X(net4557));
 sky130_fd_sc_hd__buf_1 max_length4558 (.A(net4562),
    .X(net4558));
 sky130_fd_sc_hd__clkbuf_1 wire4559 (.A(net4560),
    .X(net4559));
 sky130_fd_sc_hd__buf_1 wire4560 (.A(net4561),
    .X(net4560));
 sky130_fd_sc_hd__buf_1 wire4561 (.A(net4562),
    .X(net4561));
 sky130_fd_sc_hd__buf_1 wire4562 (.A(net4556),
    .X(net4562));
 sky130_fd_sc_hd__buf_1 wire4563 (.A(net4564),
    .X(net4563));
 sky130_fd_sc_hd__clkbuf_1 wire4564 (.A(net4556),
    .X(net4564));
 sky130_fd_sc_hd__buf_1 wire4565 (.A(net4566),
    .X(net4565));
 sky130_fd_sc_hd__clkbuf_1 wire4566 (.A(net4567),
    .X(net4566));
 sky130_fd_sc_hd__clkbuf_1 wire4567 (.A(net4569),
    .X(net4567));
 sky130_fd_sc_hd__clkbuf_1 max_length4568 (.A(net4569),
    .X(net4568));
 sky130_fd_sc_hd__buf_1 max_length4569 (.A(\pid_q.mult0.a[11] ),
    .X(net4569));
 sky130_fd_sc_hd__buf_1 fanout4570 (.A(net4577),
    .X(net4570));
 sky130_fd_sc_hd__clkbuf_1 wire4571 (.A(net4574),
    .X(net4571));
 sky130_fd_sc_hd__clkbuf_1 wire4572 (.A(net4573),
    .X(net4572));
 sky130_fd_sc_hd__buf_1 wire4573 (.A(net4574),
    .X(net4573));
 sky130_fd_sc_hd__buf_1 wire4574 (.A(net4570),
    .X(net4574));
 sky130_fd_sc_hd__buf_1 wire4575 (.A(net4576),
    .X(net4575));
 sky130_fd_sc_hd__buf_1 wire4576 (.A(net4570),
    .X(net4576));
 sky130_fd_sc_hd__clkbuf_1 fanout4577 (.A(\pid_q.mult0.a[10] ),
    .X(net4577));
 sky130_fd_sc_hd__clkbuf_1 wire4578 (.A(net4579),
    .X(net4578));
 sky130_fd_sc_hd__buf_1 wire4579 (.A(net4580),
    .X(net4579));
 sky130_fd_sc_hd__buf_1 wire4580 (.A(net4581),
    .X(net4580));
 sky130_fd_sc_hd__buf_1 wire4581 (.A(net4582),
    .X(net4581));
 sky130_fd_sc_hd__clkbuf_1 wire4582 (.A(net4583),
    .X(net4582));
 sky130_fd_sc_hd__clkbuf_1 wire4583 (.A(net4584),
    .X(net4583));
 sky130_fd_sc_hd__clkbuf_1 wire4584 (.A(net4585),
    .X(net4584));
 sky130_fd_sc_hd__clkbuf_1 wire4585 (.A(net4586),
    .X(net4585));
 sky130_fd_sc_hd__clkbuf_1 max_length4586 (.A(net4577),
    .X(net4586));
 sky130_fd_sc_hd__clkbuf_1 wire4587 (.A(\pid_q.mult0.a[10] ),
    .X(net4587));
 sky130_fd_sc_hd__buf_1 fanout4588 (.A(net4594),
    .X(net4588));
 sky130_fd_sc_hd__buf_1 wire4589 (.A(net4590),
    .X(net4589));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4590 (.A(net4591),
    .X(net4590));
 sky130_fd_sc_hd__buf_1 wire4591 (.A(net4592),
    .X(net4591));
 sky130_fd_sc_hd__buf_1 wire4592 (.A(net4593),
    .X(net4592));
 sky130_fd_sc_hd__clkbuf_1 wire4593 (.A(net4588),
    .X(net4593));
 sky130_fd_sc_hd__buf_1 fanout4594 (.A(\pid_q.mult0.a[9] ),
    .X(net4594));
 sky130_fd_sc_hd__buf_1 wire4595 (.A(net4594),
    .X(net4595));
 sky130_fd_sc_hd__clkbuf_1 wire4596 (.A(net4599),
    .X(net4596));
 sky130_fd_sc_hd__buf_1 wire4597 (.A(net4598),
    .X(net4597));
 sky130_fd_sc_hd__buf_1 wire4598 (.A(net4599),
    .X(net4598));
 sky130_fd_sc_hd__buf_1 wire4599 (.A(net4594),
    .X(net4599));
 sky130_fd_sc_hd__clkbuf_1 wire4600 (.A(net4601),
    .X(net4600));
 sky130_fd_sc_hd__clkbuf_1 wire4601 (.A(\pid_q.mult0.a[9] ),
    .X(net4601));
 sky130_fd_sc_hd__clkbuf_1 fanout4602 (.A(net4609),
    .X(net4602));
 sky130_fd_sc_hd__buf_1 wire4603 (.A(net4604),
    .X(net4603));
 sky130_fd_sc_hd__buf_1 wire4604 (.A(net4605),
    .X(net4604));
 sky130_fd_sc_hd__buf_1 wire4605 (.A(net4606),
    .X(net4605));
 sky130_fd_sc_hd__buf_1 wire4606 (.A(net4607),
    .X(net4606));
 sky130_fd_sc_hd__clkbuf_1 wire4607 (.A(net4608),
    .X(net4607));
 sky130_fd_sc_hd__buf_1 wire4608 (.A(net4602),
    .X(net4608));
 sky130_fd_sc_hd__buf_1 fanout4609 (.A(\pid_q.mult0.a[8] ),
    .X(net4609));
 sky130_fd_sc_hd__buf_1 wire4610 (.A(net4613),
    .X(net4610));
 sky130_fd_sc_hd__clkbuf_1 wire4611 (.A(net4612),
    .X(net4611));
 sky130_fd_sc_hd__clkbuf_1 max_length4612 (.A(net4613),
    .X(net4612));
 sky130_fd_sc_hd__buf_1 wire4613 (.A(net4609),
    .X(net4613));
 sky130_fd_sc_hd__clkbuf_1 wire4614 (.A(net4615),
    .X(net4614));
 sky130_fd_sc_hd__buf_1 wire4615 (.A(net4616),
    .X(net4615));
 sky130_fd_sc_hd__buf_1 wire4616 (.A(net4617),
    .X(net4616));
 sky130_fd_sc_hd__buf_1 wire4617 (.A(net4618),
    .X(net4617));
 sky130_fd_sc_hd__buf_1 wire4618 (.A(net4609),
    .X(net4618));
 sky130_fd_sc_hd__buf_1 wire4619 (.A(net4620),
    .X(net4619));
 sky130_fd_sc_hd__clkbuf_1 wire4620 (.A(net4621),
    .X(net4620));
 sky130_fd_sc_hd__clkbuf_1 wire4621 (.A(net4622),
    .X(net4621));
 sky130_fd_sc_hd__clkbuf_1 max_length4622 (.A(\pid_q.mult0.a[8] ),
    .X(net4622));
 sky130_fd_sc_hd__buf_1 fanout4623 (.A(net4633),
    .X(net4623));
 sky130_fd_sc_hd__buf_1 wire4624 (.A(net4625),
    .X(net4624));
 sky130_fd_sc_hd__buf_1 wire4625 (.A(net4626),
    .X(net4625));
 sky130_fd_sc_hd__buf_1 wire4626 (.A(net4627),
    .X(net4626));
 sky130_fd_sc_hd__clkbuf_1 wire4627 (.A(net4628),
    .X(net4627));
 sky130_fd_sc_hd__clkbuf_1 wire4628 (.A(net4629),
    .X(net4628));
 sky130_fd_sc_hd__buf_1 max_length4629 (.A(net4623),
    .X(net4629));
 sky130_fd_sc_hd__buf_1 fanout4630 (.A(\pid_q.mult0.a[7] ),
    .X(net4630));
 sky130_fd_sc_hd__buf_1 wire4631 (.A(net4632),
    .X(net4631));
 sky130_fd_sc_hd__clkbuf_1 wire4632 (.A(net4633),
    .X(net4632));
 sky130_fd_sc_hd__buf_1 wire4633 (.A(net4634),
    .X(net4633));
 sky130_fd_sc_hd__buf_1 wire4634 (.A(net4630),
    .X(net4634));
 sky130_fd_sc_hd__clkbuf_1 wire4635 (.A(net4638),
    .X(net4635));
 sky130_fd_sc_hd__buf_1 wire4636 (.A(net4637),
    .X(net4636));
 sky130_fd_sc_hd__buf_1 wire4637 (.A(net4638),
    .X(net4637));
 sky130_fd_sc_hd__buf_1 wire4638 (.A(net4630),
    .X(net4638));
 sky130_fd_sc_hd__buf_1 fanout4639 (.A(net4643),
    .X(net4639));
 sky130_fd_sc_hd__clkbuf_1 wire4640 (.A(net4639),
    .X(net4640));
 sky130_fd_sc_hd__buf_1 wire4641 (.A(net4642),
    .X(net4641));
 sky130_fd_sc_hd__clkbuf_1 wire4642 (.A(net4639),
    .X(net4642));
 sky130_fd_sc_hd__clkbuf_1 wire4643 (.A(net4644),
    .X(net4643));
 sky130_fd_sc_hd__clkbuf_1 wire4644 (.A(net4645),
    .X(net4644));
 sky130_fd_sc_hd__clkbuf_1 max_length4645 (.A(\pid_q.mult0.a[7] ),
    .X(net4645));
 sky130_fd_sc_hd__clkbuf_1 fanout4646 (.A(net4668),
    .X(net4646));
 sky130_fd_sc_hd__buf_1 wire4647 (.A(net4654),
    .X(net4647));
 sky130_fd_sc_hd__clkbuf_1 wire4648 (.A(net4649),
    .X(net4648));
 sky130_fd_sc_hd__clkbuf_1 wire4649 (.A(net4650),
    .X(net4649));
 sky130_fd_sc_hd__clkbuf_1 wire4650 (.A(net4652),
    .X(net4650));
 sky130_fd_sc_hd__buf_1 wire4651 (.A(net4652),
    .X(net4651));
 sky130_fd_sc_hd__buf_1 wire4652 (.A(net4653),
    .X(net4652));
 sky130_fd_sc_hd__clkbuf_1 wire4653 (.A(net4655),
    .X(net4653));
 sky130_fd_sc_hd__buf_1 max_length4654 (.A(net4655),
    .X(net4654));
 sky130_fd_sc_hd__buf_1 wire4655 (.A(net4646),
    .X(net4655));
 sky130_fd_sc_hd__clkbuf_1 fanout4656 (.A(\pid_q.mult0.a[6] ),
    .X(net4656));
 sky130_fd_sc_hd__clkbuf_1 wire4657 (.A(net4658),
    .X(net4657));
 sky130_fd_sc_hd__clkbuf_1 wire4658 (.A(net4659),
    .X(net4658));
 sky130_fd_sc_hd__clkbuf_1 wire4659 (.A(net4660),
    .X(net4659));
 sky130_fd_sc_hd__clkbuf_1 wire4660 (.A(net4668),
    .X(net4660));
 sky130_fd_sc_hd__clkbuf_1 wire4661 (.A(net4667),
    .X(net4661));
 sky130_fd_sc_hd__buf_1 wire4662 (.A(net4666),
    .X(net4662));
 sky130_fd_sc_hd__clkbuf_1 wire4663 (.A(net4665),
    .X(net4663));
 sky130_fd_sc_hd__buf_1 wire4664 (.A(net4665),
    .X(net4664));
 sky130_fd_sc_hd__buf_1 wire4665 (.A(net4666),
    .X(net4665));
 sky130_fd_sc_hd__buf_1 wire4666 (.A(net4667),
    .X(net4666));
 sky130_fd_sc_hd__buf_1 wire4667 (.A(net4668),
    .X(net4667));
 sky130_fd_sc_hd__buf_1 wire4668 (.A(net4656),
    .X(net4668));
 sky130_fd_sc_hd__buf_1 wire4669 (.A(net4670),
    .X(net4669));
 sky130_fd_sc_hd__clkbuf_1 wire4670 (.A(net4671),
    .X(net4670));
 sky130_fd_sc_hd__clkbuf_1 wire4671 (.A(net4672),
    .X(net4671));
 sky130_fd_sc_hd__clkbuf_1 wire4672 (.A(\pid_q.mult0.a[6] ),
    .X(net4672));
 sky130_fd_sc_hd__buf_1 fanout4673 (.A(net4686),
    .X(net4673));
 sky130_fd_sc_hd__buf_1 wire4674 (.A(net4675),
    .X(net4674));
 sky130_fd_sc_hd__buf_1 wire4675 (.A(net4676),
    .X(net4675));
 sky130_fd_sc_hd__buf_1 wire4676 (.A(net4673),
    .X(net4676));
 sky130_fd_sc_hd__buf_1 wire4677 (.A(net4678),
    .X(net4677));
 sky130_fd_sc_hd__clkbuf_1 wire4678 (.A(net4679),
    .X(net4678));
 sky130_fd_sc_hd__buf_1 max_length4679 (.A(net4673),
    .X(net4679));
 sky130_fd_sc_hd__buf_1 fanout4680 (.A(\pid_q.mult0.a[5] ),
    .X(net4680));
 sky130_fd_sc_hd__buf_1 wire4681 (.A(net4682),
    .X(net4681));
 sky130_fd_sc_hd__clkbuf_1 wire4682 (.A(net4683),
    .X(net4682));
 sky130_fd_sc_hd__buf_1 wire4683 (.A(net4684),
    .X(net4683));
 sky130_fd_sc_hd__buf_1 wire4684 (.A(net4685),
    .X(net4684));
 sky130_fd_sc_hd__buf_1 wire4685 (.A(net4687),
    .X(net4685));
 sky130_fd_sc_hd__clkbuf_1 wire4686 (.A(net4680),
    .X(net4686));
 sky130_fd_sc_hd__buf_1 max_length4687 (.A(net4680),
    .X(net4687));
 sky130_fd_sc_hd__buf_1 wire4688 (.A(net4689),
    .X(net4688));
 sky130_fd_sc_hd__clkbuf_1 wire4689 (.A(net4690),
    .X(net4689));
 sky130_fd_sc_hd__clkbuf_1 wire4690 (.A(net4691),
    .X(net4690));
 sky130_fd_sc_hd__clkbuf_1 wire4691 (.A(\pid_q.mult0.a[5] ),
    .X(net4691));
 sky130_fd_sc_hd__buf_1 fanout4692 (.A(net4714),
    .X(net4692));
 sky130_fd_sc_hd__buf_1 wire4693 (.A(net4694),
    .X(net4693));
 sky130_fd_sc_hd__buf_1 wire4694 (.A(net4695),
    .X(net4694));
 sky130_fd_sc_hd__clkbuf_1 wire4695 (.A(net4692),
    .X(net4695));
 sky130_fd_sc_hd__clkbuf_1 wire4696 (.A(net4697),
    .X(net4696));
 sky130_fd_sc_hd__buf_1 wire4697 (.A(net4698),
    .X(net4697));
 sky130_fd_sc_hd__buf_1 wire4698 (.A(net4699),
    .X(net4698));
 sky130_fd_sc_hd__clkbuf_1 wire4699 (.A(net4700),
    .X(net4699));
 sky130_fd_sc_hd__buf_1 max_length4700 (.A(net4692),
    .X(net4700));
 sky130_fd_sc_hd__clkbuf_1 fanout4701 (.A(\pid_q.mult0.a[4] ),
    .X(net4701));
 sky130_fd_sc_hd__buf_1 wire4702 (.A(net4703),
    .X(net4702));
 sky130_fd_sc_hd__buf_1 wire4703 (.A(net4704),
    .X(net4703));
 sky130_fd_sc_hd__clkbuf_2 wire4704 (.A(net4705),
    .X(net4704));
 sky130_fd_sc_hd__clkbuf_1 wire4705 (.A(net4706),
    .X(net4705));
 sky130_fd_sc_hd__clkbuf_1 max_length4706 (.A(net4707),
    .X(net4706));
 sky130_fd_sc_hd__buf_1 wire4707 (.A(net4701),
    .X(net4707));
 sky130_fd_sc_hd__clkbuf_1 wire4708 (.A(net4709),
    .X(net4708));
 sky130_fd_sc_hd__clkbuf_1 wire4709 (.A(net4710),
    .X(net4709));
 sky130_fd_sc_hd__clkbuf_1 wire4710 (.A(net4711),
    .X(net4710));
 sky130_fd_sc_hd__clkbuf_1 wire4711 (.A(\pid_q.mult0.a[4] ),
    .X(net4711));
 sky130_fd_sc_hd__clkbuf_1 wire4712 (.A(net4713),
    .X(net4712));
 sky130_fd_sc_hd__clkbuf_1 max_length4713 (.A(net4714),
    .X(net4713));
 sky130_fd_sc_hd__buf_1 wire4714 (.A(\pid_q.mult0.a[4] ),
    .X(net4714));
 sky130_fd_sc_hd__buf_1 fanout4715 (.A(net4725),
    .X(net4715));
 sky130_fd_sc_hd__buf_1 wire4716 (.A(net4717),
    .X(net4716));
 sky130_fd_sc_hd__buf_1 wire4717 (.A(net4718),
    .X(net4717));
 sky130_fd_sc_hd__buf_1 wire4718 (.A(net4715),
    .X(net4718));
 sky130_fd_sc_hd__buf_1 wire4719 (.A(net4720),
    .X(net4719));
 sky130_fd_sc_hd__clkbuf_1 wire4720 (.A(net4715),
    .X(net4720));
 sky130_fd_sc_hd__clkbuf_1 fanout4721 (.A(net4732),
    .X(net4721));
 sky130_fd_sc_hd__clkbuf_1 max_length4722 (.A(net4723),
    .X(net4722));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4723 (.A(net4721),
    .X(net4723));
 sky130_fd_sc_hd__clkbuf_1 fanout4724 (.A(\pid_q.mult0.a[3] ),
    .X(net4724));
 sky130_fd_sc_hd__clkbuf_1 wire4725 (.A(net4726),
    .X(net4725));
 sky130_fd_sc_hd__clkbuf_1 wire4726 (.A(net4733),
    .X(net4726));
 sky130_fd_sc_hd__buf_1 wire4727 (.A(net4728),
    .X(net4727));
 sky130_fd_sc_hd__clkbuf_1 max_length4728 (.A(net4729),
    .X(net4728));
 sky130_fd_sc_hd__clkbuf_2 wire4729 (.A(net4730),
    .X(net4729));
 sky130_fd_sc_hd__clkbuf_1 wire4730 (.A(net4731),
    .X(net4730));
 sky130_fd_sc_hd__clkbuf_1 wire4731 (.A(net4732),
    .X(net4731));
 sky130_fd_sc_hd__buf_1 wire4732 (.A(net4733),
    .X(net4732));
 sky130_fd_sc_hd__buf_1 wire4733 (.A(net4724),
    .X(net4733));
 sky130_fd_sc_hd__buf_1 fanout4734 (.A(net4745),
    .X(net4734));
 sky130_fd_sc_hd__clkbuf_1 wire4735 (.A(net4736),
    .X(net4735));
 sky130_fd_sc_hd__buf_1 wire4736 (.A(net4737),
    .X(net4736));
 sky130_fd_sc_hd__clkbuf_1 wire4737 (.A(net4734),
    .X(net4737));
 sky130_fd_sc_hd__buf_1 wire4738 (.A(net4739),
    .X(net4738));
 sky130_fd_sc_hd__buf_1 wire4739 (.A(net4740),
    .X(net4739));
 sky130_fd_sc_hd__buf_1 max_length4740 (.A(net4734),
    .X(net4740));
 sky130_fd_sc_hd__buf_1 fanout4741 (.A(net4747),
    .X(net4741));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4742 (.A(net4743),
    .X(net4742));
 sky130_fd_sc_hd__buf_1 wire4743 (.A(net4741),
    .X(net4743));
 sky130_fd_sc_hd__buf_1 fanout4744 (.A(\pid_q.mult0.a[2] ),
    .X(net4744));
 sky130_fd_sc_hd__clkbuf_1 wire4745 (.A(net4746),
    .X(net4745));
 sky130_fd_sc_hd__clkbuf_1 wire4746 (.A(net4747),
    .X(net4746));
 sky130_fd_sc_hd__buf_1 wire4747 (.A(net4744),
    .X(net4747));
 sky130_fd_sc_hd__buf_1 wire4748 (.A(net4749),
    .X(net4748));
 sky130_fd_sc_hd__buf_1 wire4749 (.A(net4750),
    .X(net4749));
 sky130_fd_sc_hd__clkbuf_1 wire4750 (.A(net4751),
    .X(net4750));
 sky130_fd_sc_hd__clkbuf_1 wire4751 (.A(net4752),
    .X(net4751));
 sky130_fd_sc_hd__clkbuf_1 wire4752 (.A(net4744),
    .X(net4752));
 sky130_fd_sc_hd__buf_1 fanout4753 (.A(net4762),
    .X(net4753));
 sky130_fd_sc_hd__buf_1 wire4754 (.A(net4755),
    .X(net4754));
 sky130_fd_sc_hd__buf_1 wire4755 (.A(net4753),
    .X(net4755));
 sky130_fd_sc_hd__clkbuf_1 wire4756 (.A(net4757),
    .X(net4756));
 sky130_fd_sc_hd__buf_1 wire4757 (.A(net4758),
    .X(net4757));
 sky130_fd_sc_hd__buf_1 wire4758 (.A(net4753),
    .X(net4758));
 sky130_fd_sc_hd__clkbuf_1 fanout4759 (.A(net4764),
    .X(net4759));
 sky130_fd_sc_hd__buf_1 wire4760 (.A(net4759),
    .X(net4760));
 sky130_fd_sc_hd__clkbuf_1 fanout4761 (.A(\pid_q.mult0.a[1] ),
    .X(net4761));
 sky130_fd_sc_hd__clkbuf_1 wire4762 (.A(net4763),
    .X(net4762));
 sky130_fd_sc_hd__clkbuf_1 wire4763 (.A(net4765),
    .X(net4763));
 sky130_fd_sc_hd__clkbuf_1 wire4764 (.A(net4765),
    .X(net4764));
 sky130_fd_sc_hd__buf_1 wire4765 (.A(net4766),
    .X(net4765));
 sky130_fd_sc_hd__clkbuf_1 wire4766 (.A(net4767),
    .X(net4766));
 sky130_fd_sc_hd__buf_1 wire4767 (.A(net4761),
    .X(net4767));
 sky130_fd_sc_hd__buf_1 wire4768 (.A(net4769),
    .X(net4768));
 sky130_fd_sc_hd__clkbuf_1 wire4769 (.A(net4770),
    .X(net4769));
 sky130_fd_sc_hd__clkbuf_1 wire4770 (.A(net4761),
    .X(net4770));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout4771 (.A(net4780),
    .X(net4771));
 sky130_fd_sc_hd__clkbuf_2 wire4772 (.A(net4771),
    .X(net4772));
 sky130_fd_sc_hd__buf_1 fanout4773 (.A(net4780),
    .X(net4773));
 sky130_fd_sc_hd__clkbuf_1 wire4774 (.A(net4775),
    .X(net4774));
 sky130_fd_sc_hd__buf_1 wire4775 (.A(net4777),
    .X(net4775));
 sky130_fd_sc_hd__buf_1 wire4776 (.A(net4777),
    .X(net4776));
 sky130_fd_sc_hd__buf_1 wire4777 (.A(net4778),
    .X(net4777));
 sky130_fd_sc_hd__buf_1 wire4778 (.A(net4773),
    .X(net4778));
 sky130_fd_sc_hd__buf_1 fanout4779 (.A(\pid_q.mult0.a[0] ),
    .X(net4779));
 sky130_fd_sc_hd__buf_1 wire4780 (.A(net4781),
    .X(net4780));
 sky130_fd_sc_hd__clkbuf_1 wire4781 (.A(net4782),
    .X(net4781));
 sky130_fd_sc_hd__clkbuf_1 wire4782 (.A(net4783),
    .X(net4782));
 sky130_fd_sc_hd__clkbuf_1 wire4783 (.A(net4779),
    .X(net4783));
 sky130_fd_sc_hd__buf_1 wire4784 (.A(net4785),
    .X(net4784));
 sky130_fd_sc_hd__clkbuf_1 wire4785 (.A(net4786),
    .X(net4785));
 sky130_fd_sc_hd__clkbuf_1 wire4786 (.A(net4779),
    .X(net4786));
 sky130_fd_sc_hd__buf_1 fanout4787 (.A(\pid_q.mult0.b[15] ),
    .X(net4787));
 sky130_fd_sc_hd__buf_1 wire4788 (.A(net4789),
    .X(net4788));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4789 (.A(net4791),
    .X(net4789));
 sky130_fd_sc_hd__clkbuf_1 wire4790 (.A(net4792),
    .X(net4790));
 sky130_fd_sc_hd__buf_1 max_length4791 (.A(net4792),
    .X(net4791));
 sky130_fd_sc_hd__buf_1 wire4792 (.A(net4793),
    .X(net4792));
 sky130_fd_sc_hd__buf_1 max_length4793 (.A(net4794),
    .X(net4793));
 sky130_fd_sc_hd__buf_1 max_length4794 (.A(net4787),
    .X(net4794));
 sky130_fd_sc_hd__buf_1 wire4795 (.A(net4796),
    .X(net4795));
 sky130_fd_sc_hd__buf_1 wire4796 (.A(net4797),
    .X(net4796));
 sky130_fd_sc_hd__clkbuf_1 wire4797 (.A(\pid_q.mult0.b[15] ),
    .X(net4797));
 sky130_fd_sc_hd__buf_1 fanout4798 (.A(net4817),
    .X(net4798));
 sky130_fd_sc_hd__clkbuf_1 wire4799 (.A(net4800),
    .X(net4799));
 sky130_fd_sc_hd__clkbuf_1 wire4800 (.A(net4805),
    .X(net4800));
 sky130_fd_sc_hd__clkbuf_1 wire4801 (.A(net4802),
    .X(net4801));
 sky130_fd_sc_hd__buf_1 wire4802 (.A(net4803),
    .X(net4802));
 sky130_fd_sc_hd__buf_1 wire4803 (.A(net4804),
    .X(net4803));
 sky130_fd_sc_hd__buf_1 max_length4804 (.A(net4805),
    .X(net4804));
 sky130_fd_sc_hd__buf_1 wire4805 (.A(net4798),
    .X(net4805));
 sky130_fd_sc_hd__clkbuf_1 fanout4806 (.A(net4814),
    .X(net4806));
 sky130_fd_sc_hd__buf_1 wire4807 (.A(net4808),
    .X(net4807));
 sky130_fd_sc_hd__buf_1 wire4808 (.A(net4809),
    .X(net4808));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4809 (.A(net4806),
    .X(net4809));
 sky130_fd_sc_hd__buf_1 fanout4810 (.A(net4819),
    .X(net4810));
 sky130_fd_sc_hd__buf_1 wire4811 (.A(net4812),
    .X(net4811));
 sky130_fd_sc_hd__buf_1 wire4812 (.A(net4810),
    .X(net4812));
 sky130_fd_sc_hd__buf_1 wire4813 (.A(net4810),
    .X(net4813));
 sky130_fd_sc_hd__buf_1 fanout4814 (.A(\pid_q.mult0.b[14] ),
    .X(net4814));
 sky130_fd_sc_hd__clkbuf_1 wire4815 (.A(net4816),
    .X(net4815));
 sky130_fd_sc_hd__buf_1 wire4816 (.A(net4817),
    .X(net4816));
 sky130_fd_sc_hd__buf_1 wire4817 (.A(net4818),
    .X(net4817));
 sky130_fd_sc_hd__clkbuf_1 wire4818 (.A(net4814),
    .X(net4818));
 sky130_fd_sc_hd__clkbuf_1 wire4819 (.A(net4820),
    .X(net4819));
 sky130_fd_sc_hd__clkbuf_1 wire4820 (.A(net4814),
    .X(net4820));
 sky130_fd_sc_hd__buf_1 fanout4821 (.A(net4829),
    .X(net4821));
 sky130_fd_sc_hd__clkbuf_1 wire4822 (.A(net4821),
    .X(net4822));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4823 (.A(net4824),
    .X(net4823));
 sky130_fd_sc_hd__buf_1 wire4824 (.A(net4825),
    .X(net4824));
 sky130_fd_sc_hd__buf_1 wire4825 (.A(net4821),
    .X(net4825));
 sky130_fd_sc_hd__buf_1 fanout4826 (.A(net4832),
    .X(net4826));
 sky130_fd_sc_hd__buf_1 wire4827 (.A(net4828),
    .X(net4827));
 sky130_fd_sc_hd__buf_1 wire4828 (.A(net4826),
    .X(net4828));
 sky130_fd_sc_hd__buf_1 fanout4829 (.A(\pid_q.mult0.b[13] ),
    .X(net4829));
 sky130_fd_sc_hd__clkbuf_1 wire4830 (.A(net4831),
    .X(net4830));
 sky130_fd_sc_hd__clkbuf_1 wire4831 (.A(net4832),
    .X(net4831));
 sky130_fd_sc_hd__buf_1 wire4832 (.A(net4840),
    .X(net4832));
 sky130_fd_sc_hd__clkbuf_1 wire4833 (.A(net4834),
    .X(net4833));
 sky130_fd_sc_hd__buf_1 wire4834 (.A(net4835),
    .X(net4834));
 sky130_fd_sc_hd__buf_1 max_length4835 (.A(net4836),
    .X(net4835));
 sky130_fd_sc_hd__buf_1 wire4836 (.A(net4837),
    .X(net4836));
 sky130_fd_sc_hd__buf_1 wire4837 (.A(net4838),
    .X(net4837));
 sky130_fd_sc_hd__clkbuf_1 wire4838 (.A(net4839),
    .X(net4838));
 sky130_fd_sc_hd__clkbuf_1 wire4839 (.A(net4829),
    .X(net4839));
 sky130_fd_sc_hd__clkbuf_1 max_length4840 (.A(net4829),
    .X(net4840));
 sky130_fd_sc_hd__clkbuf_1 fanout4841 (.A(net4849),
    .X(net4841));
 sky130_fd_sc_hd__buf_1 wire4842 (.A(net4843),
    .X(net4842));
 sky130_fd_sc_hd__buf_1 max_length4843 (.A(net4844),
    .X(net4843));
 sky130_fd_sc_hd__buf_1 wire4844 (.A(net4848),
    .X(net4844));
 sky130_fd_sc_hd__buf_1 wire4845 (.A(net4846),
    .X(net4845));
 sky130_fd_sc_hd__buf_1 wire4846 (.A(net4847),
    .X(net4846));
 sky130_fd_sc_hd__clkbuf_1 max_length4847 (.A(net4848),
    .X(net4847));
 sky130_fd_sc_hd__buf_1 max_length4848 (.A(net4841),
    .X(net4848));
 sky130_fd_sc_hd__clkbuf_1 fanout4849 (.A(net4861),
    .X(net4849));
 sky130_fd_sc_hd__buf_1 wire4850 (.A(net4851),
    .X(net4850));
 sky130_fd_sc_hd__buf_1 wire4851 (.A(net4852),
    .X(net4851));
 sky130_fd_sc_hd__buf_1 wire4852 (.A(net4853),
    .X(net4852));
 sky130_fd_sc_hd__buf_1 wire4853 (.A(net4857),
    .X(net4853));
 sky130_fd_sc_hd__clkbuf_1 wire4854 (.A(net4855),
    .X(net4854));
 sky130_fd_sc_hd__buf_1 wire4855 (.A(net4856),
    .X(net4855));
 sky130_fd_sc_hd__clkbuf_1 wire4856 (.A(net4857),
    .X(net4856));
 sky130_fd_sc_hd__buf_1 wire4857 (.A(net4858),
    .X(net4857));
 sky130_fd_sc_hd__clkbuf_1 wire4858 (.A(net4849),
    .X(net4858));
 sky130_fd_sc_hd__clkbuf_1 wire4859 (.A(net4860),
    .X(net4859));
 sky130_fd_sc_hd__clkbuf_1 wire4860 (.A(net4861),
    .X(net4860));
 sky130_fd_sc_hd__buf_1 wire4861 (.A(\pid_q.mult0.b[12] ),
    .X(net4861));
 sky130_fd_sc_hd__buf_1 fanout4862 (.A(net4883),
    .X(net4862));
 sky130_fd_sc_hd__clkbuf_1 wire4863 (.A(net4864),
    .X(net4863));
 sky130_fd_sc_hd__buf_1 max_length4864 (.A(net4865),
    .X(net4864));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4865 (.A(net4866),
    .X(net4865));
 sky130_fd_sc_hd__buf_1 wire4866 (.A(net4867),
    .X(net4866));
 sky130_fd_sc_hd__buf_1 wire4867 (.A(net4862),
    .X(net4867));
 sky130_fd_sc_hd__clkbuf_1 wire4868 (.A(net4869),
    .X(net4868));
 sky130_fd_sc_hd__clkbuf_1 wire4869 (.A(net4870),
    .X(net4869));
 sky130_fd_sc_hd__clkbuf_1 wire4870 (.A(net4862),
    .X(net4870));
 sky130_fd_sc_hd__clkbuf_2 fanout4871 (.A(net4878),
    .X(net4871));
 sky130_fd_sc_hd__buf_1 wire4872 (.A(net4871),
    .X(net4872));
 sky130_fd_sc_hd__buf_1 wire4873 (.A(net4871),
    .X(net4873));
 sky130_fd_sc_hd__buf_1 fanout4874 (.A(net4879),
    .X(net4874));
 sky130_fd_sc_hd__buf_1 wire4875 (.A(net4876),
    .X(net4875));
 sky130_fd_sc_hd__buf_1 wire4876 (.A(net4877),
    .X(net4876));
 sky130_fd_sc_hd__clkbuf_1 wire4877 (.A(net4874),
    .X(net4877));
 sky130_fd_sc_hd__clkbuf_1 max_length4878 (.A(net4874),
    .X(net4878));
 sky130_fd_sc_hd__buf_1 fanout4879 (.A(\pid_q.mult0.b[11] ),
    .X(net4879));
 sky130_fd_sc_hd__buf_1 wire4880 (.A(net4881),
    .X(net4880));
 sky130_fd_sc_hd__buf_1 wire4881 (.A(net4882),
    .X(net4881));
 sky130_fd_sc_hd__clkbuf_1 wire4882 (.A(net4883),
    .X(net4882));
 sky130_fd_sc_hd__buf_1 wire4883 (.A(net4884),
    .X(net4883));
 sky130_fd_sc_hd__clkbuf_1 wire4884 (.A(net4879),
    .X(net4884));
 sky130_fd_sc_hd__buf_1 fanout4885 (.A(net4908),
    .X(net4885));
 sky130_fd_sc_hd__clkbuf_1 wire4886 (.A(net4887),
    .X(net4886));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4887 (.A(net4888),
    .X(net4887));
 sky130_fd_sc_hd__buf_1 wire4888 (.A(net4889),
    .X(net4888));
 sky130_fd_sc_hd__buf_1 wire4889 (.A(net4890),
    .X(net4889));
 sky130_fd_sc_hd__buf_1 wire4890 (.A(net4885),
    .X(net4890));
 sky130_fd_sc_hd__clkbuf_1 wire4891 (.A(net4892),
    .X(net4891));
 sky130_fd_sc_hd__clkbuf_1 wire4892 (.A(net4893),
    .X(net4892));
 sky130_fd_sc_hd__clkbuf_1 wire4893 (.A(net4885),
    .X(net4893));
 sky130_fd_sc_hd__buf_1 fanout4894 (.A(net4898),
    .X(net4894));
 sky130_fd_sc_hd__clkbuf_1 max_length4895 (.A(net4896),
    .X(net4895));
 sky130_fd_sc_hd__clkbuf_2 wire4896 (.A(net4894),
    .X(net4896));
 sky130_fd_sc_hd__buf_1 fanout4897 (.A(net4903),
    .X(net4897));
 sky130_fd_sc_hd__clkbuf_1 wire4898 (.A(net4897),
    .X(net4898));
 sky130_fd_sc_hd__buf_1 wire4899 (.A(net4900),
    .X(net4899));
 sky130_fd_sc_hd__buf_1 wire4900 (.A(net4901),
    .X(net4900));
 sky130_fd_sc_hd__clkbuf_1 wire4901 (.A(net4902),
    .X(net4901));
 sky130_fd_sc_hd__clkbuf_1 max_length4902 (.A(net4897),
    .X(net4902));
 sky130_fd_sc_hd__buf_1 fanout4903 (.A(\pid_q.mult0.b[10] ),
    .X(net4903));
 sky130_fd_sc_hd__clkbuf_1 wire4904 (.A(net4905),
    .X(net4904));
 sky130_fd_sc_hd__buf_1 wire4905 (.A(net4906),
    .X(net4905));
 sky130_fd_sc_hd__buf_1 wire4906 (.A(net4907),
    .X(net4906));
 sky130_fd_sc_hd__clkbuf_1 wire4907 (.A(net4908),
    .X(net4907));
 sky130_fd_sc_hd__buf_1 wire4908 (.A(net4909),
    .X(net4908));
 sky130_fd_sc_hd__clkbuf_1 wire4909 (.A(net4910),
    .X(net4909));
 sky130_fd_sc_hd__clkbuf_1 wire4910 (.A(net4903),
    .X(net4910));
 sky130_fd_sc_hd__buf_1 fanout4911 (.A(net4927),
    .X(net4911));
 sky130_fd_sc_hd__buf_1 wire4912 (.A(net4913),
    .X(net4912));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4913 (.A(net4915),
    .X(net4913));
 sky130_fd_sc_hd__clkbuf_1 wire4914 (.A(net4915),
    .X(net4914));
 sky130_fd_sc_hd__buf_1 max_length4915 (.A(net4911),
    .X(net4915));
 sky130_fd_sc_hd__clkbuf_1 fanout4916 (.A(net4923),
    .X(net4916));
 sky130_fd_sc_hd__buf_1 wire4917 (.A(net4918),
    .X(net4917));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4918 (.A(net4919),
    .X(net4918));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire4919 (.A(net4916),
    .X(net4919));
 sky130_fd_sc_hd__buf_1 fanout4920 (.A(net4924),
    .X(net4920));
 sky130_fd_sc_hd__clkbuf_1 wire4921 (.A(net4922),
    .X(net4921));
 sky130_fd_sc_hd__buf_1 wire4922 (.A(net4920),
    .X(net4922));
 sky130_fd_sc_hd__buf_1 fanout4923 (.A(\pid_q.mult0.b[9] ),
    .X(net4923));
 sky130_fd_sc_hd__clkbuf_1 wire4924 (.A(net4925),
    .X(net4924));
 sky130_fd_sc_hd__clkbuf_1 wire4925 (.A(net4923),
    .X(net4925));
 sky130_fd_sc_hd__buf_1 wire4926 (.A(net4927),
    .X(net4926));
 sky130_fd_sc_hd__buf_1 wire4927 (.A(net4929),
    .X(net4927));
 sky130_fd_sc_hd__buf_1 max_length4928 (.A(net4929),
    .X(net4928));
 sky130_fd_sc_hd__buf_1 wire4929 (.A(net4930),
    .X(net4929));
 sky130_fd_sc_hd__clkbuf_1 wire4930 (.A(net4931),
    .X(net4930));
 sky130_fd_sc_hd__clkbuf_1 wire4931 (.A(net4932),
    .X(net4931));
 sky130_fd_sc_hd__clkbuf_1 wire4932 (.A(net4923),
    .X(net4932));
 sky130_fd_sc_hd__buf_1 fanout4933 (.A(net4945),
    .X(net4933));
 sky130_fd_sc_hd__buf_1 wire4934 (.A(net4935),
    .X(net4934));
 sky130_fd_sc_hd__clkbuf_1 wire4935 (.A(net4936),
    .X(net4935));
 sky130_fd_sc_hd__clkbuf_1 wire4936 (.A(net4939),
    .X(net4936));
 sky130_fd_sc_hd__clkbuf_2 wire4937 (.A(net4938),
    .X(net4937));
 sky130_fd_sc_hd__clkbuf_1 wire4938 (.A(net4933),
    .X(net4938));
 sky130_fd_sc_hd__clkbuf_1 max_length4939 (.A(net4933),
    .X(net4939));
 sky130_fd_sc_hd__clkbuf_1 fanout4940 (.A(net4946),
    .X(net4940));
 sky130_fd_sc_hd__buf_1 wire4941 (.A(net4942),
    .X(net4941));
 sky130_fd_sc_hd__buf_1 wire4942 (.A(net4943),
    .X(net4942));
 sky130_fd_sc_hd__clkbuf_1 max_length4943 (.A(net4944),
    .X(net4943));
 sky130_fd_sc_hd__buf_1 max_length4944 (.A(net4940),
    .X(net4944));
 sky130_fd_sc_hd__buf_1 fanout4945 (.A(\pid_q.mult0.b[8] ),
    .X(net4945));
 sky130_fd_sc_hd__clkbuf_1 wire4946 (.A(net4947),
    .X(net4946));
 sky130_fd_sc_hd__clkbuf_1 wire4947 (.A(net4945),
    .X(net4947));
 sky130_fd_sc_hd__buf_1 wire4948 (.A(net4949),
    .X(net4948));
 sky130_fd_sc_hd__buf_1 wire4949 (.A(net4950),
    .X(net4949));
 sky130_fd_sc_hd__clkbuf_1 wire4950 (.A(net4951),
    .X(net4950));
 sky130_fd_sc_hd__buf_1 wire4951 (.A(net4952),
    .X(net4951));
 sky130_fd_sc_hd__buf_1 max_length4952 (.A(net4953),
    .X(net4952));
 sky130_fd_sc_hd__buf_1 wire4953 (.A(net4954),
    .X(net4953));
 sky130_fd_sc_hd__clkbuf_1 wire4954 (.A(net4955),
    .X(net4954));
 sky130_fd_sc_hd__clkbuf_1 wire4955 (.A(net4945),
    .X(net4955));
 sky130_fd_sc_hd__clkbuf_1 fanout4956 (.A(\pid_q.mult0.b[7] ),
    .X(net4956));
 sky130_fd_sc_hd__buf_1 wire4957 (.A(net4958),
    .X(net4957));
 sky130_fd_sc_hd__clkbuf_1 wire4958 (.A(net4959),
    .X(net4958));
 sky130_fd_sc_hd__clkbuf_2 max_length4959 (.A(net4960),
    .X(net4959));
 sky130_fd_sc_hd__buf_1 wire4960 (.A(net4961),
    .X(net4960));
 sky130_fd_sc_hd__clkbuf_1 wire4961 (.A(net4956),
    .X(net4961));
 sky130_fd_sc_hd__buf_1 fanout4962 (.A(net4976),
    .X(net4962));
 sky130_fd_sc_hd__clkbuf_1 wire4963 (.A(net4964),
    .X(net4963));
 sky130_fd_sc_hd__buf_1 wire4964 (.A(net4962),
    .X(net4964));
 sky130_fd_sc_hd__clkbuf_1 fanout4965 (.A(net4977),
    .X(net4965));
 sky130_fd_sc_hd__clkbuf_1 wire4966 (.A(net4967),
    .X(net4966));
 sky130_fd_sc_hd__buf_1 wire4967 (.A(net4968),
    .X(net4967));
 sky130_fd_sc_hd__buf_1 wire4968 (.A(net4969),
    .X(net4968));
 sky130_fd_sc_hd__buf_1 wire4969 (.A(net4973),
    .X(net4969));
 sky130_fd_sc_hd__clkbuf_1 max_length4970 (.A(net4971),
    .X(net4970));
 sky130_fd_sc_hd__buf_1 wire4971 (.A(net4972),
    .X(net4971));
 sky130_fd_sc_hd__buf_1 wire4972 (.A(net4973),
    .X(net4972));
 sky130_fd_sc_hd__buf_1 wire4973 (.A(net4974),
    .X(net4973));
 sky130_fd_sc_hd__clkbuf_1 wire4974 (.A(net4975),
    .X(net4974));
 sky130_fd_sc_hd__clkbuf_1 wire4975 (.A(net4976),
    .X(net4975));
 sky130_fd_sc_hd__buf_1 wire4976 (.A(net4965),
    .X(net4976));
 sky130_fd_sc_hd__clkbuf_1 wire4977 (.A(net4978),
    .X(net4977));
 sky130_fd_sc_hd__clkbuf_1 wire4978 (.A(net4979),
    .X(net4978));
 sky130_fd_sc_hd__clkbuf_1 wire4979 (.A(\pid_q.mult0.b[7] ),
    .X(net4979));
 sky130_fd_sc_hd__buf_1 fanout4980 (.A(net5005),
    .X(net4980));
 sky130_fd_sc_hd__buf_1 max_length4981 (.A(net4982),
    .X(net4981));
 sky130_fd_sc_hd__buf_1 wire4982 (.A(net4984),
    .X(net4982));
 sky130_fd_sc_hd__buf_1 wire4983 (.A(net4984),
    .X(net4983));
 sky130_fd_sc_hd__buf_1 wire4984 (.A(net4985),
    .X(net4984));
 sky130_fd_sc_hd__clkbuf_1 wire4985 (.A(net4986),
    .X(net4985));
 sky130_fd_sc_hd__buf_1 wire4986 (.A(net4987),
    .X(net4986));
 sky130_fd_sc_hd__buf_1 wire4987 (.A(net4980),
    .X(net4987));
 sky130_fd_sc_hd__clkbuf_1 fanout4988 (.A(net4999),
    .X(net4988));
 sky130_fd_sc_hd__clkbuf_1 wire4989 (.A(net4990),
    .X(net4989));
 sky130_fd_sc_hd__buf_1 wire4990 (.A(net4991),
    .X(net4990));
 sky130_fd_sc_hd__buf_1 wire4991 (.A(net4992),
    .X(net4991));
 sky130_fd_sc_hd__clkbuf_1 wire4992 (.A(net4993),
    .X(net4992));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length4993 (.A(net4994),
    .X(net4993));
 sky130_fd_sc_hd__buf_1 wire4994 (.A(net4995),
    .X(net4994));
 sky130_fd_sc_hd__clkbuf_1 wire4995 (.A(net4988),
    .X(net4995));
 sky130_fd_sc_hd__buf_1 fanout4996 (.A(net5008),
    .X(net4996));
 sky130_fd_sc_hd__buf_1 wire4997 (.A(net4998),
    .X(net4997));
 sky130_fd_sc_hd__buf_1 wire4998 (.A(net4996),
    .X(net4998));
 sky130_fd_sc_hd__buf_1 fanout4999 (.A(\pid_q.mult0.b[6] ),
    .X(net4999));
 sky130_fd_sc_hd__buf_1 wire5000 (.A(net5001),
    .X(net5000));
 sky130_fd_sc_hd__buf_1 wire5001 (.A(net5002),
    .X(net5001));
 sky130_fd_sc_hd__clkbuf_1 wire5002 (.A(net5003),
    .X(net5002));
 sky130_fd_sc_hd__clkbuf_1 wire5003 (.A(net5004),
    .X(net5003));
 sky130_fd_sc_hd__clkbuf_1 wire5004 (.A(net5005),
    .X(net5004));
 sky130_fd_sc_hd__buf_1 wire5005 (.A(net5006),
    .X(net5005));
 sky130_fd_sc_hd__clkbuf_1 wire5006 (.A(net5007),
    .X(net5006));
 sky130_fd_sc_hd__clkbuf_1 wire5007 (.A(net4999),
    .X(net5007));
 sky130_fd_sc_hd__clkbuf_1 wire5008 (.A(net5009),
    .X(net5008));
 sky130_fd_sc_hd__clkbuf_1 wire5009 (.A(net5010),
    .X(net5009));
 sky130_fd_sc_hd__clkbuf_1 wire5010 (.A(net4999),
    .X(net5010));
 sky130_fd_sc_hd__buf_1 fanout5011 (.A(net5027),
    .X(net5011));
 sky130_fd_sc_hd__buf_1 wire5012 (.A(net5013),
    .X(net5012));
 sky130_fd_sc_hd__buf_1 wire5013 (.A(net5014),
    .X(net5013));
 sky130_fd_sc_hd__clkbuf_1 wire5014 (.A(net5019),
    .X(net5014));
 sky130_fd_sc_hd__buf_1 wire5015 (.A(net5016),
    .X(net5015));
 sky130_fd_sc_hd__buf_1 wire5016 (.A(net5017),
    .X(net5016));
 sky130_fd_sc_hd__buf_1 wire5017 (.A(net5018),
    .X(net5017));
 sky130_fd_sc_hd__clkbuf_1 wire5018 (.A(net5020),
    .X(net5018));
 sky130_fd_sc_hd__clkbuf_1 max_length5019 (.A(net5020),
    .X(net5019));
 sky130_fd_sc_hd__buf_1 max_length5020 (.A(net5011),
    .X(net5020));
 sky130_fd_sc_hd__buf_1 fanout5021 (.A(\pid_q.mult0.b[5] ),
    .X(net5021));
 sky130_fd_sc_hd__buf_1 wire5022 (.A(net5023),
    .X(net5022));
 sky130_fd_sc_hd__buf_1 wire5023 (.A(net5025),
    .X(net5023));
 sky130_fd_sc_hd__buf_1 wire5024 (.A(net5025),
    .X(net5024));
 sky130_fd_sc_hd__buf_1 wire5025 (.A(net5026),
    .X(net5025));
 sky130_fd_sc_hd__clkbuf_1 wire5026 (.A(net5030),
    .X(net5026));
 sky130_fd_sc_hd__buf_1 wire5027 (.A(net5028),
    .X(net5027));
 sky130_fd_sc_hd__buf_1 wire5028 (.A(net5029),
    .X(net5028));
 sky130_fd_sc_hd__clkbuf_1 wire5029 (.A(net5030),
    .X(net5029));
 sky130_fd_sc_hd__buf_1 wire5030 (.A(net5021),
    .X(net5030));
 sky130_fd_sc_hd__clkbuf_1 wire5031 (.A(net5032),
    .X(net5031));
 sky130_fd_sc_hd__clkbuf_1 wire5032 (.A(net5034),
    .X(net5032));
 sky130_fd_sc_hd__clkbuf_1 wire5033 (.A(net5034),
    .X(net5033));
 sky130_fd_sc_hd__buf_1 wire5034 (.A(net5035),
    .X(net5034));
 sky130_fd_sc_hd__clkbuf_1 wire5035 (.A(\pid_q.mult0.b[5] ),
    .X(net5035));
 sky130_fd_sc_hd__buf_1 fanout5036 (.A(net5047),
    .X(net5036));
 sky130_fd_sc_hd__buf_1 wire5037 (.A(net5038),
    .X(net5037));
 sky130_fd_sc_hd__buf_1 wire5038 (.A(net5039),
    .X(net5038));
 sky130_fd_sc_hd__buf_1 wire5039 (.A(net5040),
    .X(net5039));
 sky130_fd_sc_hd__buf_1 wire5040 (.A(net5042),
    .X(net5040));
 sky130_fd_sc_hd__clkbuf_1 wire5041 (.A(net5042),
    .X(net5041));
 sky130_fd_sc_hd__buf_1 wire5042 (.A(net5036),
    .X(net5042));
 sky130_fd_sc_hd__buf_1 fanout5043 (.A(\pid_q.mult0.b[4] ),
    .X(net5043));
 sky130_fd_sc_hd__clkbuf_1 wire5044 (.A(net5045),
    .X(net5044));
 sky130_fd_sc_hd__clkbuf_1 wire5045 (.A(net5046),
    .X(net5045));
 sky130_fd_sc_hd__clkbuf_1 wire5046 (.A(net5047),
    .X(net5046));
 sky130_fd_sc_hd__clkbuf_1 wire5047 (.A(net5048),
    .X(net5047));
 sky130_fd_sc_hd__buf_1 wire5048 (.A(net5049),
    .X(net5048));
 sky130_fd_sc_hd__clkbuf_1 wire5049 (.A(net5050),
    .X(net5049));
 sky130_fd_sc_hd__clkbuf_1 wire5050 (.A(net5056),
    .X(net5050));
 sky130_fd_sc_hd__clkbuf_1 wire5051 (.A(net5052),
    .X(net5051));
 sky130_fd_sc_hd__buf_1 wire5052 (.A(net5053),
    .X(net5052));
 sky130_fd_sc_hd__buf_1 wire5053 (.A(net5054),
    .X(net5053));
 sky130_fd_sc_hd__buf_1 wire5054 (.A(net5055),
    .X(net5054));
 sky130_fd_sc_hd__clkbuf_1 wire5055 (.A(net5043),
    .X(net5055));
 sky130_fd_sc_hd__clkbuf_1 max_length5056 (.A(net5043),
    .X(net5056));
 sky130_fd_sc_hd__buf_1 wire5057 (.A(net5058),
    .X(net5057));
 sky130_fd_sc_hd__clkbuf_1 wire5058 (.A(net5059),
    .X(net5058));
 sky130_fd_sc_hd__buf_1 wire5059 (.A(net5060),
    .X(net5059));
 sky130_fd_sc_hd__clkbuf_1 wire5060 (.A(\pid_q.mult0.b[4] ),
    .X(net5060));
 sky130_fd_sc_hd__clkbuf_1 fanout5061 (.A(net5073),
    .X(net5061));
 sky130_fd_sc_hd__buf_1 wire5062 (.A(net5063),
    .X(net5062));
 sky130_fd_sc_hd__buf_1 wire5063 (.A(net5064),
    .X(net5063));
 sky130_fd_sc_hd__buf_1 wire5064 (.A(net5065),
    .X(net5064));
 sky130_fd_sc_hd__buf_1 wire5065 (.A(net5066),
    .X(net5065));
 sky130_fd_sc_hd__buf_1 wire5066 (.A(net5061),
    .X(net5066));
 sky130_fd_sc_hd__clkbuf_1 fanout5067 (.A(net5074),
    .X(net5067));
 sky130_fd_sc_hd__clkbuf_1 max_length5068 (.A(net5069),
    .X(net5068));
 sky130_fd_sc_hd__buf_1 wire5069 (.A(net5070),
    .X(net5069));
 sky130_fd_sc_hd__buf_1 wire5070 (.A(net5071),
    .X(net5070));
 sky130_fd_sc_hd__buf_1 wire5071 (.A(net5067),
    .X(net5071));
 sky130_fd_sc_hd__buf_1 fanout5072 (.A(\pid_q.mult0.b[3] ),
    .X(net5072));
 sky130_fd_sc_hd__clkbuf_1 max_length5073 (.A(net5074),
    .X(net5073));
 sky130_fd_sc_hd__buf_1 wire5074 (.A(net5075),
    .X(net5074));
 sky130_fd_sc_hd__buf_1 wire5075 (.A(net5076),
    .X(net5075));
 sky130_fd_sc_hd__clkbuf_1 wire5076 (.A(net5072),
    .X(net5076));
 sky130_fd_sc_hd__buf_1 wire5077 (.A(net5078),
    .X(net5077));
 sky130_fd_sc_hd__buf_1 wire5078 (.A(net5079),
    .X(net5078));
 sky130_fd_sc_hd__buf_1 wire5079 (.A(net5080),
    .X(net5079));
 sky130_fd_sc_hd__buf_1 wire5080 (.A(net5081),
    .X(net5080));
 sky130_fd_sc_hd__clkbuf_1 wire5081 (.A(net5082),
    .X(net5081));
 sky130_fd_sc_hd__clkbuf_1 wire5082 (.A(net5072),
    .X(net5082));
 sky130_fd_sc_hd__clkbuf_1 fanout5083 (.A(net5104),
    .X(net5083));
 sky130_fd_sc_hd__buf_1 wire5084 (.A(net5090),
    .X(net5084));
 sky130_fd_sc_hd__clkbuf_1 wire5085 (.A(net5088),
    .X(net5085));
 sky130_fd_sc_hd__clkbuf_1 max_length5086 (.A(net5087),
    .X(net5086));
 sky130_fd_sc_hd__buf_1 wire5087 (.A(net5088),
    .X(net5087));
 sky130_fd_sc_hd__buf_1 wire5088 (.A(net5089),
    .X(net5088));
 sky130_fd_sc_hd__buf_1 wire5089 (.A(net5090),
    .X(net5089));
 sky130_fd_sc_hd__buf_1 wire5090 (.A(net5083),
    .X(net5090));
 sky130_fd_sc_hd__clkbuf_1 fanout5091 (.A(net5103),
    .X(net5091));
 sky130_fd_sc_hd__clkbuf_1 wire5092 (.A(net5093),
    .X(net5092));
 sky130_fd_sc_hd__clkbuf_1 wire5093 (.A(net5095),
    .X(net5093));
 sky130_fd_sc_hd__clkbuf_1 wire5094 (.A(net5096),
    .X(net5094));
 sky130_fd_sc_hd__buf_1 max_length5095 (.A(net5096),
    .X(net5095));
 sky130_fd_sc_hd__buf_1 wire5096 (.A(net5097),
    .X(net5096));
 sky130_fd_sc_hd__buf_1 wire5097 (.A(net5098),
    .X(net5097));
 sky130_fd_sc_hd__clkbuf_1 wire5098 (.A(net5102),
    .X(net5098));
 sky130_fd_sc_hd__buf_1 wire5099 (.A(net5100),
    .X(net5099));
 sky130_fd_sc_hd__clkbuf_1 wire5100 (.A(net5101),
    .X(net5100));
 sky130_fd_sc_hd__clkbuf_1 wire5101 (.A(net5102),
    .X(net5101));
 sky130_fd_sc_hd__buf_1 max_length5102 (.A(net5091),
    .X(net5102));
 sky130_fd_sc_hd__clkbuf_1 fanout5103 (.A(\pid_q.mult0.b[2] ),
    .X(net5103));
 sky130_fd_sc_hd__buf_1 wire5104 (.A(net5105),
    .X(net5104));
 sky130_fd_sc_hd__clkbuf_1 wire5105 (.A(net5106),
    .X(net5105));
 sky130_fd_sc_hd__clkbuf_1 wire5106 (.A(net5107),
    .X(net5106));
 sky130_fd_sc_hd__clkbuf_1 wire5107 (.A(net5110),
    .X(net5107));
 sky130_fd_sc_hd__buf_1 wire5108 (.A(net5109),
    .X(net5108));
 sky130_fd_sc_hd__clkbuf_1 wire5109 (.A(net5110),
    .X(net5109));
 sky130_fd_sc_hd__buf_1 wire5110 (.A(net5103),
    .X(net5110));
 sky130_fd_sc_hd__buf_1 fanout5111 (.A(net5135),
    .X(net5111));
 sky130_fd_sc_hd__buf_1 wire5112 (.A(net5116),
    .X(net5112));
 sky130_fd_sc_hd__clkbuf_1 wire5113 (.A(net5114),
    .X(net5113));
 sky130_fd_sc_hd__clkbuf_1 wire5114 (.A(net5115),
    .X(net5114));
 sky130_fd_sc_hd__buf_1 wire5115 (.A(net5116),
    .X(net5115));
 sky130_fd_sc_hd__clkbuf_2 wire5116 (.A(net5111),
    .X(net5116));
 sky130_fd_sc_hd__buf_1 fanout5117 (.A(net5127),
    .X(net5117));
 sky130_fd_sc_hd__clkbuf_1 wire5118 (.A(net5119),
    .X(net5118));
 sky130_fd_sc_hd__clkbuf_1 wire5119 (.A(net5121),
    .X(net5119));
 sky130_fd_sc_hd__buf_1 wire5120 (.A(net5121),
    .X(net5120));
 sky130_fd_sc_hd__buf_1 wire5121 (.A(net5122),
    .X(net5121));
 sky130_fd_sc_hd__buf_1 wire5122 (.A(net5123),
    .X(net5122));
 sky130_fd_sc_hd__clkbuf_1 wire5123 (.A(net5117),
    .X(net5123));
 sky130_fd_sc_hd__buf_1 wire5124 (.A(net5125),
    .X(net5124));
 sky130_fd_sc_hd__clkbuf_1 wire5125 (.A(net5126),
    .X(net5125));
 sky130_fd_sc_hd__clkbuf_1 max_length5126 (.A(net5117),
    .X(net5126));
 sky130_fd_sc_hd__clkbuf_1 fanout5127 (.A(\pid_q.mult0.b[1] ),
    .X(net5127));
 sky130_fd_sc_hd__clkbuf_1 wire5128 (.A(net5129),
    .X(net5128));
 sky130_fd_sc_hd__buf_1 wire5129 (.A(net5138),
    .X(net5129));
 sky130_fd_sc_hd__clkbuf_1 wire5130 (.A(net5131),
    .X(net5130));
 sky130_fd_sc_hd__clkbuf_1 wire5131 (.A(net5132),
    .X(net5131));
 sky130_fd_sc_hd__buf_1 wire5132 (.A(net5133),
    .X(net5132));
 sky130_fd_sc_hd__buf_1 wire5133 (.A(net5134),
    .X(net5133));
 sky130_fd_sc_hd__clkbuf_1 wire5134 (.A(net5135),
    .X(net5134));
 sky130_fd_sc_hd__buf_1 wire5135 (.A(net5136),
    .X(net5135));
 sky130_fd_sc_hd__clkbuf_1 wire5136 (.A(net5137),
    .X(net5136));
 sky130_fd_sc_hd__clkbuf_1 wire5137 (.A(net5138),
    .X(net5137));
 sky130_fd_sc_hd__buf_1 wire5138 (.A(net5127),
    .X(net5138));
 sky130_fd_sc_hd__buf_1 fanout5139 (.A(net5157),
    .X(net5139));
 sky130_fd_sc_hd__buf_1 wire5140 (.A(net5139),
    .X(net5140));
 sky130_fd_sc_hd__buf_1 max_length5141 (.A(net5142),
    .X(net5141));
 sky130_fd_sc_hd__buf_1 wire5142 (.A(net5145),
    .X(net5142));
 sky130_fd_sc_hd__buf_1 wire5143 (.A(net5144),
    .X(net5143));
 sky130_fd_sc_hd__clkbuf_1 max_length5144 (.A(net5145),
    .X(net5144));
 sky130_fd_sc_hd__buf_1 wire5145 (.A(net5139),
    .X(net5145));
 sky130_fd_sc_hd__clkbuf_1 fanout5146 (.A(net5161),
    .X(net5146));
 sky130_fd_sc_hd__clkbuf_1 wire5147 (.A(net5148),
    .X(net5147));
 sky130_fd_sc_hd__clkbuf_1 wire5148 (.A(net5149),
    .X(net5148));
 sky130_fd_sc_hd__clkbuf_2 wire5149 (.A(net5155),
    .X(net5149));
 sky130_fd_sc_hd__clkbuf_1 wire5150 (.A(net5151),
    .X(net5150));
 sky130_fd_sc_hd__clkbuf_1 wire5151 (.A(net5152),
    .X(net5151));
 sky130_fd_sc_hd__clkbuf_1 wire5152 (.A(net5153),
    .X(net5152));
 sky130_fd_sc_hd__clkbuf_1 wire5153 (.A(net5154),
    .X(net5153));
 sky130_fd_sc_hd__buf_1 wire5154 (.A(net5155),
    .X(net5154));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5155 (.A(net5146),
    .X(net5155));
 sky130_fd_sc_hd__buf_1 fanout5156 (.A(\pid_q.mult0.b[0] ),
    .X(net5156));
 sky130_fd_sc_hd__buf_1 wire5157 (.A(net5158),
    .X(net5157));
 sky130_fd_sc_hd__buf_1 wire5158 (.A(net5159),
    .X(net5158));
 sky130_fd_sc_hd__clkbuf_1 wire5159 (.A(net5160),
    .X(net5159));
 sky130_fd_sc_hd__clkbuf_1 wire5160 (.A(net5161),
    .X(net5160));
 sky130_fd_sc_hd__buf_1 wire5161 (.A(net5165),
    .X(net5161));
 sky130_fd_sc_hd__buf_1 wire5162 (.A(net5163),
    .X(net5162));
 sky130_fd_sc_hd__buf_1 wire5163 (.A(net5164),
    .X(net5163));
 sky130_fd_sc_hd__clkbuf_1 max_length5164 (.A(net5165),
    .X(net5164));
 sky130_fd_sc_hd__buf_1 wire5165 (.A(net5156),
    .X(net5165));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length5166 (.A(\pid_q.curr_error[13] ),
    .X(net5166));
 sky130_fd_sc_hd__buf_1 wire5167 (.A(\pid_q.curr_error[12] ),
    .X(net5167));
 sky130_fd_sc_hd__clkbuf_2 wire5168 (.A(\pid_q.curr_error[1] ),
    .X(net5168));
 sky130_fd_sc_hd__clkbuf_2 wire5169 (.A(\pid_q.curr_int[15] ),
    .X(net5169));
 sky130_fd_sc_hd__clkbuf_2 wire5170 (.A(net5171),
    .X(net5170));
 sky130_fd_sc_hd__buf_1 wire5171 (.A(\pid_q.curr_int[14] ),
    .X(net5171));
 sky130_fd_sc_hd__clkbuf_2 wire5172 (.A(net5173),
    .X(net5172));
 sky130_fd_sc_hd__buf_1 wire5173 (.A(\pid_q.curr_int[13] ),
    .X(net5173));
 sky130_fd_sc_hd__clkbuf_2 wire5174 (.A(net5175),
    .X(net5174));
 sky130_fd_sc_hd__clkbuf_2 wire5175 (.A(\pid_q.curr_int[12] ),
    .X(net5175));
 sky130_fd_sc_hd__buf_1 wire5176 (.A(net5177),
    .X(net5176));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5177 (.A(\pid_q.curr_int[11] ),
    .X(net5177));
 sky130_fd_sc_hd__clkbuf_2 wire5178 (.A(\pid_q.curr_int[7] ),
    .X(net5178));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5179 (.A(net5180),
    .X(net5179));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length5180 (.A(\pid_q.curr_int[2] ),
    .X(net5180));
 sky130_fd_sc_hd__buf_1 wire5181 (.A(net5182),
    .X(net5181));
 sky130_fd_sc_hd__buf_1 max_length5182 (.A(\pid_q.curr_int[1] ),
    .X(net5182));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5183 (.A(net5184),
    .X(net5183));
 sky130_fd_sc_hd__buf_1 wire5184 (.A(\pid_q.curr_int[0] ),
    .X(net5184));
 sky130_fd_sc_hd__buf_1 wire5185 (.A(net5186),
    .X(net5185));
 sky130_fd_sc_hd__clkbuf_1 wire5186 (.A(net5187),
    .X(net5186));
 sky130_fd_sc_hd__clkbuf_1 wire5187 (.A(net5188),
    .X(net5187));
 sky130_fd_sc_hd__clkbuf_1 wire5188 (.A(\svm0.in_valid ),
    .X(net5188));
 sky130_fd_sc_hd__clkbuf_2 max_length5189 (.A(net5190),
    .X(net5189));
 sky130_fd_sc_hd__buf_1 wire5190 (.A(net5191),
    .X(net5190));
 sky130_fd_sc_hd__clkbuf_1 wire5191 (.A(net5192),
    .X(net5191));
 sky130_fd_sc_hd__buf_1 wire5192 (.A(\matmul0.beta_pass[15] ),
    .X(net5192));
 sky130_fd_sc_hd__clkbuf_1 wire5193 (.A(net5194),
    .X(net5193));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5194 (.A(net5195),
    .X(net5194));
 sky130_fd_sc_hd__buf_1 wire5195 (.A(net5196),
    .X(net5195));
 sky130_fd_sc_hd__clkbuf_1 wire5196 (.A(net5197),
    .X(net5196));
 sky130_fd_sc_hd__buf_1 max_length5197 (.A(\matmul0.beta_pass[14] ),
    .X(net5197));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5198 (.A(net5200),
    .X(net5198));
 sky130_fd_sc_hd__clkbuf_1 wire5199 (.A(net5200),
    .X(net5199));
 sky130_fd_sc_hd__buf_1 wire5200 (.A(net5201),
    .X(net5200));
 sky130_fd_sc_hd__clkbuf_1 wire5201 (.A(net5203),
    .X(net5201));
 sky130_fd_sc_hd__clkbuf_1 max_length5202 (.A(net5203),
    .X(net5202));
 sky130_fd_sc_hd__buf_1 max_length5203 (.A(\matmul0.beta_pass[13] ),
    .X(net5203));
 sky130_fd_sc_hd__clkbuf_1 wire5204 (.A(net5205),
    .X(net5204));
 sky130_fd_sc_hd__clkbuf_1 wire5205 (.A(net5207),
    .X(net5205));
 sky130_fd_sc_hd__buf_1 max_length5206 (.A(net5207),
    .X(net5206));
 sky130_fd_sc_hd__clkbuf_2 wire5207 (.A(net5208),
    .X(net5207));
 sky130_fd_sc_hd__clkbuf_1 wire5208 (.A(net5209),
    .X(net5208));
 sky130_fd_sc_hd__clkbuf_1 wire5209 (.A(\matmul0.beta_pass[12] ),
    .X(net5209));
 sky130_fd_sc_hd__clkbuf_1 wire5210 (.A(net5211),
    .X(net5210));
 sky130_fd_sc_hd__clkbuf_1 wire5211 (.A(net5212),
    .X(net5211));
 sky130_fd_sc_hd__clkbuf_1 max_length5212 (.A(\matmul0.beta_pass[12] ),
    .X(net5212));
 sky130_fd_sc_hd__buf_1 wire5213 (.A(net5214),
    .X(net5213));
 sky130_fd_sc_hd__buf_1 wire5214 (.A(net5215),
    .X(net5214));
 sky130_fd_sc_hd__clkbuf_2 wire5215 (.A(net5216),
    .X(net5215));
 sky130_fd_sc_hd__clkbuf_1 wire5216 (.A(net5217),
    .X(net5216));
 sky130_fd_sc_hd__clkbuf_1 wire5217 (.A(net5218),
    .X(net5217));
 sky130_fd_sc_hd__clkbuf_1 max_length5218 (.A(\matmul0.beta_pass[11] ),
    .X(net5218));
 sky130_fd_sc_hd__buf_1 fanout5219 (.A(\matmul0.beta_pass[10] ),
    .X(net5219));
 sky130_fd_sc_hd__buf_1 wire5220 (.A(net5221),
    .X(net5220));
 sky130_fd_sc_hd__clkbuf_1 wire5221 (.A(net5222),
    .X(net5221));
 sky130_fd_sc_hd__buf_1 max_length5222 (.A(net5223),
    .X(net5222));
 sky130_fd_sc_hd__clkbuf_2 wire5223 (.A(net5224),
    .X(net5223));
 sky130_fd_sc_hd__clkbuf_1 wire5224 (.A(net5225),
    .X(net5224));
 sky130_fd_sc_hd__clkbuf_1 wire5225 (.A(net5226),
    .X(net5225));
 sky130_fd_sc_hd__clkbuf_1 wire5226 (.A(net5227),
    .X(net5226));
 sky130_fd_sc_hd__clkbuf_1 max_length5227 (.A(net5219),
    .X(net5227));
 sky130_fd_sc_hd__clkbuf_1 wire5228 (.A(net5229),
    .X(net5228));
 sky130_fd_sc_hd__clkbuf_1 wire5229 (.A(net5230),
    .X(net5229));
 sky130_fd_sc_hd__clkbuf_1 wire5230 (.A(net5231),
    .X(net5230));
 sky130_fd_sc_hd__clkbuf_1 wire5231 (.A(net5232),
    .X(net5231));
 sky130_fd_sc_hd__buf_1 wire5232 (.A(net5233),
    .X(net5232));
 sky130_fd_sc_hd__clkbuf_1 wire5233 (.A(net5234),
    .X(net5233));
 sky130_fd_sc_hd__clkbuf_1 wire5234 (.A(\matmul0.beta_pass[10] ),
    .X(net5234));
 sky130_fd_sc_hd__clkbuf_1 wire5235 (.A(net5237),
    .X(net5235));
 sky130_fd_sc_hd__clkbuf_1 wire5236 (.A(net5237),
    .X(net5236));
 sky130_fd_sc_hd__buf_1 wire5237 (.A(net5238),
    .X(net5237));
 sky130_fd_sc_hd__buf_1 wire5238 (.A(net5239),
    .X(net5238));
 sky130_fd_sc_hd__clkbuf_2 wire5239 (.A(net5240),
    .X(net5239));
 sky130_fd_sc_hd__clkbuf_1 wire5240 (.A(net5241),
    .X(net5240));
 sky130_fd_sc_hd__clkbuf_1 wire5241 (.A(net5242),
    .X(net5241));
 sky130_fd_sc_hd__clkbuf_1 wire5242 (.A(\matmul0.beta_pass[9] ),
    .X(net5242));
 sky130_fd_sc_hd__buf_1 fanout5243 (.A(\matmul0.beta_pass[8] ),
    .X(net5243));
 sky130_fd_sc_hd__clkbuf_1 wire5244 (.A(net5245),
    .X(net5244));
 sky130_fd_sc_hd__buf_1 wire5245 (.A(net5246),
    .X(net5245));
 sky130_fd_sc_hd__buf_1 wire5246 (.A(net5247),
    .X(net5246));
 sky130_fd_sc_hd__clkbuf_2 wire5247 (.A(net5248),
    .X(net5247));
 sky130_fd_sc_hd__clkbuf_1 wire5248 (.A(net5249),
    .X(net5248));
 sky130_fd_sc_hd__clkbuf_1 wire5249 (.A(net5243),
    .X(net5249));
 sky130_fd_sc_hd__buf_1 wire5250 (.A(net5251),
    .X(net5250));
 sky130_fd_sc_hd__clkbuf_1 wire5251 (.A(net5252),
    .X(net5251));
 sky130_fd_sc_hd__clkbuf_1 wire5252 (.A(\matmul0.beta_pass[8] ),
    .X(net5252));
 sky130_fd_sc_hd__clkbuf_1 max_length5253 (.A(net5254),
    .X(net5253));
 sky130_fd_sc_hd__buf_1 wire5254 (.A(net5255),
    .X(net5254));
 sky130_fd_sc_hd__buf_1 wire5255 (.A(net5256),
    .X(net5255));
 sky130_fd_sc_hd__clkbuf_1 wire5256 (.A(net5257),
    .X(net5256));
 sky130_fd_sc_hd__clkbuf_1 wire5257 (.A(net5258),
    .X(net5257));
 sky130_fd_sc_hd__clkbuf_1 wire5258 (.A(\matmul0.beta_pass[7] ),
    .X(net5258));
 sky130_fd_sc_hd__buf_1 wire5259 (.A(net5260),
    .X(net5259));
 sky130_fd_sc_hd__clkbuf_1 wire5260 (.A(net5261),
    .X(net5260));
 sky130_fd_sc_hd__clkbuf_1 wire5261 (.A(net5262),
    .X(net5261));
 sky130_fd_sc_hd__clkbuf_2 wire5262 (.A(net5263),
    .X(net5262));
 sky130_fd_sc_hd__buf_1 wire5263 (.A(net5264),
    .X(net5263));
 sky130_fd_sc_hd__clkbuf_1 wire5264 (.A(\matmul0.beta_pass[6] ),
    .X(net5264));
 sky130_fd_sc_hd__buf_1 wire5265 (.A(net5266),
    .X(net5265));
 sky130_fd_sc_hd__clkbuf_1 wire5266 (.A(net5267),
    .X(net5266));
 sky130_fd_sc_hd__buf_1 wire5267 (.A(net5269),
    .X(net5267));
 sky130_fd_sc_hd__clkbuf_1 wire5268 (.A(net5269),
    .X(net5268));
 sky130_fd_sc_hd__buf_1 wire5269 (.A(net5270),
    .X(net5269));
 sky130_fd_sc_hd__buf_1 wire5270 (.A(net5271),
    .X(net5270));
 sky130_fd_sc_hd__clkbuf_1 wire5271 (.A(net5272),
    .X(net5271));
 sky130_fd_sc_hd__buf_1 wire5272 (.A(\matmul0.beta_pass[5] ),
    .X(net5272));
 sky130_fd_sc_hd__buf_1 wire5273 (.A(net5274),
    .X(net5273));
 sky130_fd_sc_hd__clkbuf_1 wire5274 (.A(net5275),
    .X(net5274));
 sky130_fd_sc_hd__clkbuf_1 wire5275 (.A(net5277),
    .X(net5275));
 sky130_fd_sc_hd__clkbuf_1 wire5276 (.A(net5278),
    .X(net5276));
 sky130_fd_sc_hd__clkbuf_1 max_length5277 (.A(net5278),
    .X(net5277));
 sky130_fd_sc_hd__buf_1 max_length5278 (.A(net5279),
    .X(net5278));
 sky130_fd_sc_hd__buf_1 wire5279 (.A(net5280),
    .X(net5279));
 sky130_fd_sc_hd__clkbuf_1 wire5280 (.A(net5281),
    .X(net5280));
 sky130_fd_sc_hd__clkbuf_1 wire5281 (.A(net5282),
    .X(net5281));
 sky130_fd_sc_hd__buf_1 wire5282 (.A(\matmul0.beta_pass[4] ),
    .X(net5282));
 sky130_fd_sc_hd__buf_1 wire5283 (.A(net5284),
    .X(net5283));
 sky130_fd_sc_hd__buf_1 wire5284 (.A(net5285),
    .X(net5284));
 sky130_fd_sc_hd__clkbuf_1 wire5285 (.A(net5286),
    .X(net5285));
 sky130_fd_sc_hd__buf_1 wire5286 (.A(net5287),
    .X(net5286));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5287 (.A(net5288),
    .X(net5287));
 sky130_fd_sc_hd__clkbuf_1 wire5288 (.A(net5289),
    .X(net5288));
 sky130_fd_sc_hd__buf_1 wire5289 (.A(\matmul0.beta_pass[3] ),
    .X(net5289));
 sky130_fd_sc_hd__buf_1 wire5290 (.A(net5291),
    .X(net5290));
 sky130_fd_sc_hd__clkbuf_1 wire5291 (.A(net5292),
    .X(net5291));
 sky130_fd_sc_hd__clkbuf_1 wire5292 (.A(net5293),
    .X(net5292));
 sky130_fd_sc_hd__clkbuf_1 wire5293 (.A(net5294),
    .X(net5293));
 sky130_fd_sc_hd__buf_1 wire5294 (.A(net5296),
    .X(net5294));
 sky130_fd_sc_hd__clkbuf_1 wire5295 (.A(net5296),
    .X(net5295));
 sky130_fd_sc_hd__buf_1 wire5296 (.A(net5297),
    .X(net5296));
 sky130_fd_sc_hd__buf_1 wire5297 (.A(net5298),
    .X(net5297));
 sky130_fd_sc_hd__clkbuf_1 wire5298 (.A(\matmul0.beta_pass[2] ),
    .X(net5298));
 sky130_fd_sc_hd__buf_1 wire5299 (.A(net5300),
    .X(net5299));
 sky130_fd_sc_hd__clkbuf_1 wire5300 (.A(net5301),
    .X(net5300));
 sky130_fd_sc_hd__clkbuf_1 wire5301 (.A(net5302),
    .X(net5301));
 sky130_fd_sc_hd__clkbuf_1 wire5302 (.A(net5303),
    .X(net5302));
 sky130_fd_sc_hd__clkbuf_1 wire5303 (.A(net5305),
    .X(net5303));
 sky130_fd_sc_hd__clkbuf_1 max_length5304 (.A(net5305),
    .X(net5304));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5305 (.A(net5306),
    .X(net5305));
 sky130_fd_sc_hd__buf_1 wire5306 (.A(\matmul0.beta_pass[1] ),
    .X(net5306));
 sky130_fd_sc_hd__clkbuf_1 wire5307 (.A(net5308),
    .X(net5307));
 sky130_fd_sc_hd__buf_1 wire5308 (.A(net5309),
    .X(net5308));
 sky130_fd_sc_hd__clkbuf_1 wire5309 (.A(net5310),
    .X(net5309));
 sky130_fd_sc_hd__clkbuf_1 wire5310 (.A(net5313),
    .X(net5310));
 sky130_fd_sc_hd__buf_1 wire5311 (.A(net5312),
    .X(net5311));
 sky130_fd_sc_hd__buf_1 wire5312 (.A(net5313),
    .X(net5312));
 sky130_fd_sc_hd__buf_1 wire5313 (.A(\matmul0.beta_pass[0] ),
    .X(net5313));
 sky130_fd_sc_hd__buf_1 wire5314 (.A(\pid_d.out[15] ),
    .X(net5314));
 sky130_fd_sc_hd__clkbuf_1 wire5315 (.A(net5316),
    .X(net5315));
 sky130_fd_sc_hd__clkbuf_1 wire5316 (.A(net5317),
    .X(net5316));
 sky130_fd_sc_hd__clkbuf_1 wire5317 (.A(net5318),
    .X(net5317));
 sky130_fd_sc_hd__clkbuf_1 wire5318 (.A(net5319),
    .X(net5318));
 sky130_fd_sc_hd__clkbuf_1 wire5319 (.A(\pid_d.out[15] ),
    .X(net5319));
 sky130_fd_sc_hd__clkbuf_1 wire5320 (.A(net5321),
    .X(net5320));
 sky130_fd_sc_hd__clkbuf_1 wire5321 (.A(net5322),
    .X(net5321));
 sky130_fd_sc_hd__clkbuf_1 wire5322 (.A(net5323),
    .X(net5322));
 sky130_fd_sc_hd__clkbuf_1 wire5323 (.A(net5324),
    .X(net5323));
 sky130_fd_sc_hd__clkbuf_1 wire5324 (.A(net5325),
    .X(net5324));
 sky130_fd_sc_hd__clkbuf_1 wire5325 (.A(net5326),
    .X(net5325));
 sky130_fd_sc_hd__clkbuf_1 wire5326 (.A(\pid_d.out[14] ),
    .X(net5326));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5327 (.A(\pid_d.out[13] ),
    .X(net5327));
 sky130_fd_sc_hd__clkbuf_1 wire5328 (.A(net5329),
    .X(net5328));
 sky130_fd_sc_hd__clkbuf_1 wire5329 (.A(net5330),
    .X(net5329));
 sky130_fd_sc_hd__clkbuf_1 wire5330 (.A(net5331),
    .X(net5330));
 sky130_fd_sc_hd__clkbuf_1 wire5331 (.A(net5332),
    .X(net5331));
 sky130_fd_sc_hd__clkbuf_1 wire5332 (.A(\pid_d.out[13] ),
    .X(net5332));
 sky130_fd_sc_hd__clkbuf_1 wire5333 (.A(net5334),
    .X(net5333));
 sky130_fd_sc_hd__clkbuf_1 wire5334 (.A(net5335),
    .X(net5334));
 sky130_fd_sc_hd__clkbuf_1 wire5335 (.A(net5336),
    .X(net5335));
 sky130_fd_sc_hd__clkbuf_1 wire5336 (.A(net5337),
    .X(net5336));
 sky130_fd_sc_hd__clkbuf_1 wire5337 (.A(net5338),
    .X(net5337));
 sky130_fd_sc_hd__clkbuf_1 wire5338 (.A(\pid_d.out[12] ),
    .X(net5338));
 sky130_fd_sc_hd__buf_1 max_length5339 (.A(\pid_d.out[12] ),
    .X(net5339));
 sky130_fd_sc_hd__buf_1 wire5340 (.A(\pid_d.out[11] ),
    .X(net5340));
 sky130_fd_sc_hd__clkbuf_1 wire5341 (.A(net5342),
    .X(net5341));
 sky130_fd_sc_hd__clkbuf_1 wire5342 (.A(net5343),
    .X(net5342));
 sky130_fd_sc_hd__clkbuf_1 wire5343 (.A(net5344),
    .X(net5343));
 sky130_fd_sc_hd__clkbuf_1 wire5344 (.A(net5345),
    .X(net5344));
 sky130_fd_sc_hd__clkbuf_1 wire5345 (.A(\pid_d.out[11] ),
    .X(net5345));
 sky130_fd_sc_hd__clkbuf_1 wire5346 (.A(net5347),
    .X(net5346));
 sky130_fd_sc_hd__clkbuf_1 wire5347 (.A(net5348),
    .X(net5347));
 sky130_fd_sc_hd__clkbuf_1 wire5348 (.A(net5349),
    .X(net5348));
 sky130_fd_sc_hd__clkbuf_1 wire5349 (.A(net5350),
    .X(net5349));
 sky130_fd_sc_hd__clkbuf_1 max_length5350 (.A(\pid_d.out[10] ),
    .X(net5350));
 sky130_fd_sc_hd__clkbuf_1 wire5351 (.A(net5352),
    .X(net5351));
 sky130_fd_sc_hd__clkbuf_1 wire5352 (.A(net5353),
    .X(net5352));
 sky130_fd_sc_hd__clkbuf_1 wire5353 (.A(\pid_d.out[9] ),
    .X(net5353));
 sky130_fd_sc_hd__buf_1 max_length5354 (.A(\pid_d.out[9] ),
    .X(net5354));
 sky130_fd_sc_hd__clkbuf_1 wire5355 (.A(net5356),
    .X(net5355));
 sky130_fd_sc_hd__clkbuf_1 wire5356 (.A(\pid_d.out[8] ),
    .X(net5356));
 sky130_fd_sc_hd__buf_1 max_length5357 (.A(\pid_d.out[8] ),
    .X(net5357));
 sky130_fd_sc_hd__clkbuf_1 wire5358 (.A(net5359),
    .X(net5358));
 sky130_fd_sc_hd__clkbuf_1 wire5359 (.A(\pid_d.out[7] ),
    .X(net5359));
 sky130_fd_sc_hd__buf_1 max_length5360 (.A(\pid_d.out[7] ),
    .X(net5360));
 sky130_fd_sc_hd__clkbuf_1 wire5361 (.A(net5362),
    .X(net5361));
 sky130_fd_sc_hd__clkbuf_1 wire5362 (.A(\pid_d.out[6] ),
    .X(net5362));
 sky130_fd_sc_hd__buf_1 max_length5363 (.A(\pid_d.out[6] ),
    .X(net5363));
 sky130_fd_sc_hd__buf_1 wire5364 (.A(\pid_d.out[5] ),
    .X(net5364));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5365 (.A(\pid_d.out[2] ),
    .X(net5365));
 sky130_fd_sc_hd__clkbuf_2 wire5366 (.A(\pid_d.out[1] ),
    .X(net5366));
 sky130_fd_sc_hd__clkbuf_1 wire5367 (.A(net5368),
    .X(net5367));
 sky130_fd_sc_hd__clkbuf_1 wire5368 (.A(net5369),
    .X(net5368));
 sky130_fd_sc_hd__clkbuf_1 wire5369 (.A(\pid_d.out[0] ),
    .X(net5369));
 sky130_fd_sc_hd__buf_1 wire5370 (.A(net5371),
    .X(net5370));
 sky130_fd_sc_hd__clkbuf_1 max_length5371 (.A(\pid_d.out_valid ),
    .X(net5371));
 sky130_fd_sc_hd__clkbuf_1 wire5372 (.A(\pid_d.kp[15] ),
    .X(net5372));
 sky130_fd_sc_hd__clkbuf_1 wire5373 (.A(\pid_d.ki[15] ),
    .X(net5373));
 sky130_fd_sc_hd__clkbuf_1 fanout5374 (.A(\pid_d.mult0.a[15] ),
    .X(net5374));
 sky130_fd_sc_hd__buf_1 wire5375 (.A(net5377),
    .X(net5375));
 sky130_fd_sc_hd__buf_1 wire5376 (.A(net5377),
    .X(net5376));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5377 (.A(net5378),
    .X(net5377));
 sky130_fd_sc_hd__buf_1 wire5378 (.A(net5379),
    .X(net5378));
 sky130_fd_sc_hd__clkbuf_1 wire5379 (.A(net5374),
    .X(net5379));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout5380 (.A(net5381),
    .X(net5380));
 sky130_fd_sc_hd__buf_1 fanout5381 (.A(net5387),
    .X(net5381));
 sky130_fd_sc_hd__clkbuf_1 max_length5382 (.A(net5383),
    .X(net5382));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5383 (.A(net5384),
    .X(net5383));
 sky130_fd_sc_hd__buf_1 max_length5384 (.A(net5385),
    .X(net5384));
 sky130_fd_sc_hd__buf_1 wire5385 (.A(net5386),
    .X(net5385));
 sky130_fd_sc_hd__clkbuf_1 wire5386 (.A(net5381),
    .X(net5386));
 sky130_fd_sc_hd__clkbuf_1 wire5387 (.A(\pid_d.mult0.a[15] ),
    .X(net5387));
 sky130_fd_sc_hd__buf_1 fanout5388 (.A(net5392),
    .X(net5388));
 sky130_fd_sc_hd__buf_1 wire5389 (.A(net5390),
    .X(net5389));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5390 (.A(net5388),
    .X(net5390));
 sky130_fd_sc_hd__clkbuf_1 fanout5391 (.A(net5398),
    .X(net5391));
 sky130_fd_sc_hd__clkbuf_1 wire5392 (.A(net5397),
    .X(net5392));
 sky130_fd_sc_hd__buf_1 wire5393 (.A(net5394),
    .X(net5393));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length5394 (.A(net5395),
    .X(net5394));
 sky130_fd_sc_hd__buf_1 wire5395 (.A(net5396),
    .X(net5395));
 sky130_fd_sc_hd__buf_1 wire5396 (.A(net5397),
    .X(net5396));
 sky130_fd_sc_hd__buf_1 wire5397 (.A(net5391),
    .X(net5397));
 sky130_fd_sc_hd__clkbuf_1 fanout5398 (.A(\pid_d.mult0.a[14] ),
    .X(net5398));
 sky130_fd_sc_hd__buf_1 wire5399 (.A(net5400),
    .X(net5399));
 sky130_fd_sc_hd__buf_1 wire5400 (.A(net5401),
    .X(net5400));
 sky130_fd_sc_hd__buf_1 wire5401 (.A(net5402),
    .X(net5401));
 sky130_fd_sc_hd__clkbuf_1 wire5402 (.A(net5403),
    .X(net5402));
 sky130_fd_sc_hd__clkbuf_1 wire5403 (.A(net5405),
    .X(net5403));
 sky130_fd_sc_hd__clkbuf_1 max_length5404 (.A(net5405),
    .X(net5404));
 sky130_fd_sc_hd__buf_1 wire5405 (.A(net5398),
    .X(net5405));
 sky130_fd_sc_hd__clkbuf_2 fanout5406 (.A(net5421),
    .X(net5406));
 sky130_fd_sc_hd__buf_1 wire5407 (.A(net5408),
    .X(net5407));
 sky130_fd_sc_hd__buf_1 wire5408 (.A(net5406),
    .X(net5408));
 sky130_fd_sc_hd__buf_1 fanout5409 (.A(net5422),
    .X(net5409));
 sky130_fd_sc_hd__clkbuf_1 max_length5410 (.A(net5411),
    .X(net5410));
 sky130_fd_sc_hd__buf_1 wire5411 (.A(net5412),
    .X(net5411));
 sky130_fd_sc_hd__buf_1 wire5412 (.A(net5409),
    .X(net5412));
 sky130_fd_sc_hd__clkbuf_1 fanout5413 (.A(net5419),
    .X(net5413));
 sky130_fd_sc_hd__clkbuf_1 wire5414 (.A(net5415),
    .X(net5414));
 sky130_fd_sc_hd__buf_1 wire5415 (.A(net5416),
    .X(net5415));
 sky130_fd_sc_hd__clkbuf_2 wire5416 (.A(net5417),
    .X(net5416));
 sky130_fd_sc_hd__clkbuf_1 wire5417 (.A(net5418),
    .X(net5417));
 sky130_fd_sc_hd__buf_1 wire5418 (.A(net5413),
    .X(net5418));
 sky130_fd_sc_hd__clkbuf_1 wire5419 (.A(net5420),
    .X(net5419));
 sky130_fd_sc_hd__buf_1 wire5420 (.A(net5421),
    .X(net5420));
 sky130_fd_sc_hd__clkbuf_1 wire5421 (.A(net5422),
    .X(net5421));
 sky130_fd_sc_hd__buf_1 wire5422 (.A(\pid_d.mult0.a[13] ),
    .X(net5422));
 sky130_fd_sc_hd__clkbuf_1 fanout5423 (.A(net5448),
    .X(net5423));
 sky130_fd_sc_hd__clkbuf_1 wire5424 (.A(net5425),
    .X(net5424));
 sky130_fd_sc_hd__buf_1 wire5425 (.A(net5426),
    .X(net5425));
 sky130_fd_sc_hd__buf_1 wire5426 (.A(net5427),
    .X(net5426));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5427 (.A(net5428),
    .X(net5427));
 sky130_fd_sc_hd__clkbuf_1 wire5428 (.A(net5429),
    .X(net5428));
 sky130_fd_sc_hd__buf_1 max_length5429 (.A(net5423),
    .X(net5429));
 sky130_fd_sc_hd__clkbuf_1 fanout5430 (.A(net5439),
    .X(net5430));
 sky130_fd_sc_hd__buf_1 wire5431 (.A(net5432),
    .X(net5431));
 sky130_fd_sc_hd__buf_1 max_length5432 (.A(net5433),
    .X(net5432));
 sky130_fd_sc_hd__buf_1 max_length5433 (.A(net5434),
    .X(net5433));
 sky130_fd_sc_hd__buf_1 wire5434 (.A(net5435),
    .X(net5434));
 sky130_fd_sc_hd__buf_1 wire5435 (.A(net5430),
    .X(net5435));
 sky130_fd_sc_hd__clkbuf_1 fanout5436 (.A(net5452),
    .X(net5436));
 sky130_fd_sc_hd__clkbuf_1 max_length5437 (.A(net5438),
    .X(net5437));
 sky130_fd_sc_hd__buf_1 wire5438 (.A(net5439),
    .X(net5438));
 sky130_fd_sc_hd__buf_1 wire5439 (.A(net5443),
    .X(net5439));
 sky130_fd_sc_hd__clkbuf_1 wire5440 (.A(net5441),
    .X(net5440));
 sky130_fd_sc_hd__clkbuf_1 wire5441 (.A(net5442),
    .X(net5441));
 sky130_fd_sc_hd__clkbuf_1 wire5442 (.A(net5443),
    .X(net5442));
 sky130_fd_sc_hd__buf_1 wire5443 (.A(net5436),
    .X(net5443));
 sky130_fd_sc_hd__clkbuf_1 wire5444 (.A(net5445),
    .X(net5444));
 sky130_fd_sc_hd__clkbuf_1 wire5445 (.A(net5446),
    .X(net5445));
 sky130_fd_sc_hd__clkbuf_1 wire5446 (.A(net5447),
    .X(net5446));
 sky130_fd_sc_hd__clkbuf_1 wire5447 (.A(net5448),
    .X(net5447));
 sky130_fd_sc_hd__buf_1 wire5448 (.A(net5449),
    .X(net5448));
 sky130_fd_sc_hd__clkbuf_1 wire5449 (.A(net5450),
    .X(net5449));
 sky130_fd_sc_hd__clkbuf_1 wire5450 (.A(net5451),
    .X(net5450));
 sky130_fd_sc_hd__clkbuf_1 wire5451 (.A(net5452),
    .X(net5451));
 sky130_fd_sc_hd__buf_1 wire5452 (.A(\pid_d.mult0.a[12] ),
    .X(net5452));
 sky130_fd_sc_hd__clkbuf_1 fanout5453 (.A(net5467),
    .X(net5453));
 sky130_fd_sc_hd__buf_1 wire5454 (.A(net5455),
    .X(net5454));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5455 (.A(net5456),
    .X(net5455));
 sky130_fd_sc_hd__buf_1 wire5456 (.A(net5457),
    .X(net5456));
 sky130_fd_sc_hd__buf_1 wire5457 (.A(net5458),
    .X(net5457));
 sky130_fd_sc_hd__buf_1 wire5458 (.A(net5453),
    .X(net5458));
 sky130_fd_sc_hd__clkbuf_1 fanout5459 (.A(\pid_d.mult0.a[11] ),
    .X(net5459));
 sky130_fd_sc_hd__clkbuf_1 max_length5460 (.A(net5461),
    .X(net5460));
 sky130_fd_sc_hd__buf_1 wire5461 (.A(net5462),
    .X(net5461));
 sky130_fd_sc_hd__buf_1 wire5462 (.A(net5466),
    .X(net5462));
 sky130_fd_sc_hd__clkbuf_1 wire5463 (.A(net5464),
    .X(net5463));
 sky130_fd_sc_hd__buf_1 wire5464 (.A(net5465),
    .X(net5464));
 sky130_fd_sc_hd__buf_1 wire5465 (.A(net5466),
    .X(net5465));
 sky130_fd_sc_hd__buf_1 wire5466 (.A(net5459),
    .X(net5466));
 sky130_fd_sc_hd__clkbuf_1 wire5467 (.A(net5468),
    .X(net5467));
 sky130_fd_sc_hd__clkbuf_1 wire5468 (.A(net5469),
    .X(net5468));
 sky130_fd_sc_hd__clkbuf_1 wire5469 (.A(net5470),
    .X(net5469));
 sky130_fd_sc_hd__clkbuf_1 wire5470 (.A(\pid_d.mult0.a[11] ),
    .X(net5470));
 sky130_fd_sc_hd__clkbuf_1 fanout5471 (.A(net5483),
    .X(net5471));
 sky130_fd_sc_hd__buf_1 wire5472 (.A(net5473),
    .X(net5472));
 sky130_fd_sc_hd__clkbuf_2 wire5473 (.A(net5474),
    .X(net5473));
 sky130_fd_sc_hd__clkbuf_1 wire5474 (.A(net5475),
    .X(net5474));
 sky130_fd_sc_hd__buf_1 max_length5475 (.A(net5476),
    .X(net5475));
 sky130_fd_sc_hd__buf_1 wire5476 (.A(net5477),
    .X(net5476));
 sky130_fd_sc_hd__clkbuf_1 wire5477 (.A(net5471),
    .X(net5477));
 sky130_fd_sc_hd__clkbuf_1 fanout5478 (.A(net5489),
    .X(net5478));
 sky130_fd_sc_hd__buf_1 wire5479 (.A(net5480),
    .X(net5479));
 sky130_fd_sc_hd__buf_1 max_length5480 (.A(net5481),
    .X(net5480));
 sky130_fd_sc_hd__buf_1 wire5481 (.A(net5487),
    .X(net5481));
 sky130_fd_sc_hd__clkbuf_1 wire5482 (.A(net5483),
    .X(net5482));
 sky130_fd_sc_hd__buf_1 wire5483 (.A(net5484),
    .X(net5483));
 sky130_fd_sc_hd__buf_1 wire5484 (.A(net5485),
    .X(net5484));
 sky130_fd_sc_hd__buf_1 wire5485 (.A(net5486),
    .X(net5485));
 sky130_fd_sc_hd__clkbuf_1 wire5486 (.A(net5488),
    .X(net5486));
 sky130_fd_sc_hd__buf_1 max_length5487 (.A(net5488),
    .X(net5487));
 sky130_fd_sc_hd__buf_1 wire5488 (.A(net5478),
    .X(net5488));
 sky130_fd_sc_hd__buf_1 wire5489 (.A(\pid_d.mult0.a[10] ),
    .X(net5489));
 sky130_fd_sc_hd__clkbuf_1 fanout5490 (.A(net5501),
    .X(net5490));
 sky130_fd_sc_hd__buf_1 wire5491 (.A(net5492),
    .X(net5491));
 sky130_fd_sc_hd__buf_1 wire5492 (.A(net5493),
    .X(net5492));
 sky130_fd_sc_hd__clkbuf_1 wire5493 (.A(net5494),
    .X(net5493));
 sky130_fd_sc_hd__buf_1 wire5494 (.A(net5495),
    .X(net5494));
 sky130_fd_sc_hd__buf_1 wire5495 (.A(net5490),
    .X(net5495));
 sky130_fd_sc_hd__clkbuf_1 fanout5496 (.A(\pid_d.mult0.a[9] ),
    .X(net5496));
 sky130_fd_sc_hd__clkbuf_1 max_length5497 (.A(net5498),
    .X(net5497));
 sky130_fd_sc_hd__buf_1 wire5498 (.A(net5499),
    .X(net5498));
 sky130_fd_sc_hd__buf_1 wire5499 (.A(net5500),
    .X(net5499));
 sky130_fd_sc_hd__buf_1 wire5500 (.A(net5502),
    .X(net5500));
 sky130_fd_sc_hd__buf_1 wire5501 (.A(net5502),
    .X(net5501));
 sky130_fd_sc_hd__clkbuf_2 wire5502 (.A(net5503),
    .X(net5502));
 sky130_fd_sc_hd__clkbuf_1 wire5503 (.A(net5504),
    .X(net5503));
 sky130_fd_sc_hd__clkbuf_1 wire5504 (.A(net5496),
    .X(net5504));
 sky130_fd_sc_hd__buf_1 fanout5505 (.A(net5519),
    .X(net5505));
 sky130_fd_sc_hd__clkbuf_1 wire5506 (.A(net5507),
    .X(net5506));
 sky130_fd_sc_hd__buf_1 wire5507 (.A(net5508),
    .X(net5507));
 sky130_fd_sc_hd__clkbuf_1 wire5508 (.A(net5509),
    .X(net5508));
 sky130_fd_sc_hd__buf_1 wire5509 (.A(net5510),
    .X(net5509));
 sky130_fd_sc_hd__buf_1 wire5510 (.A(net5511),
    .X(net5510));
 sky130_fd_sc_hd__buf_1 wire5511 (.A(net5505),
    .X(net5511));
 sky130_fd_sc_hd__clkbuf_1 fanout5512 (.A(\pid_d.mult0.a[8] ),
    .X(net5512));
 sky130_fd_sc_hd__buf_1 wire5513 (.A(net5514),
    .X(net5513));
 sky130_fd_sc_hd__buf_1 wire5514 (.A(net5515),
    .X(net5514));
 sky130_fd_sc_hd__buf_1 wire5515 (.A(net5516),
    .X(net5515));
 sky130_fd_sc_hd__buf_1 wire5516 (.A(net5517),
    .X(net5516));
 sky130_fd_sc_hd__clkbuf_1 wire5517 (.A(net5518),
    .X(net5517));
 sky130_fd_sc_hd__clkbuf_1 wire5518 (.A(net5512),
    .X(net5518));
 sky130_fd_sc_hd__clkbuf_1 wire5519 (.A(net5520),
    .X(net5519));
 sky130_fd_sc_hd__clkbuf_1 wire5520 (.A(net5521),
    .X(net5520));
 sky130_fd_sc_hd__clkbuf_1 wire5521 (.A(net5522),
    .X(net5521));
 sky130_fd_sc_hd__clkbuf_1 wire5522 (.A(\pid_d.mult0.a[8] ),
    .X(net5522));
 sky130_fd_sc_hd__clkbuf_1 fanout5523 (.A(net5533),
    .X(net5523));
 sky130_fd_sc_hd__buf_1 wire5524 (.A(net5525),
    .X(net5524));
 sky130_fd_sc_hd__buf_1 wire5525 (.A(net5526),
    .X(net5525));
 sky130_fd_sc_hd__clkbuf_1 max_length5526 (.A(net5527),
    .X(net5526));
 sky130_fd_sc_hd__buf_1 wire5527 (.A(net5528),
    .X(net5527));
 sky130_fd_sc_hd__buf_1 wire5528 (.A(net5523),
    .X(net5528));
 sky130_fd_sc_hd__clkbuf_1 wire5529 (.A(net5530),
    .X(net5529));
 sky130_fd_sc_hd__clkbuf_1 wire5530 (.A(net5531),
    .X(net5530));
 sky130_fd_sc_hd__clkbuf_1 wire5531 (.A(net5523),
    .X(net5531));
 sky130_fd_sc_hd__clkbuf_1 fanout5532 (.A(\pid_d.mult0.a[7] ),
    .X(net5532));
 sky130_fd_sc_hd__clkbuf_1 wire5533 (.A(net5534),
    .X(net5533));
 sky130_fd_sc_hd__clkbuf_1 wire5534 (.A(net5539),
    .X(net5534));
 sky130_fd_sc_hd__buf_1 wire5535 (.A(net5536),
    .X(net5535));
 sky130_fd_sc_hd__clkbuf_1 wire5536 (.A(net5537),
    .X(net5536));
 sky130_fd_sc_hd__buf_1 wire5537 (.A(net5538),
    .X(net5537));
 sky130_fd_sc_hd__buf_1 wire5538 (.A(net5539),
    .X(net5538));
 sky130_fd_sc_hd__buf_1 wire5539 (.A(net5540),
    .X(net5539));
 sky130_fd_sc_hd__buf_1 max_length5540 (.A(net5532),
    .X(net5540));
 sky130_fd_sc_hd__buf_1 fanout5541 (.A(net5554),
    .X(net5541));
 sky130_fd_sc_hd__buf_1 wire5542 (.A(net5543),
    .X(net5542));
 sky130_fd_sc_hd__buf_1 wire5543 (.A(net5544),
    .X(net5543));
 sky130_fd_sc_hd__buf_1 wire5544 (.A(net5545),
    .X(net5544));
 sky130_fd_sc_hd__buf_1 wire5545 (.A(net5546),
    .X(net5545));
 sky130_fd_sc_hd__buf_1 wire5546 (.A(net5547),
    .X(net5546));
 sky130_fd_sc_hd__clkbuf_1 wire5547 (.A(net5541),
    .X(net5547));
 sky130_fd_sc_hd__buf_1 fanout5548 (.A(\pid_d.mult0.a[6] ),
    .X(net5548));
 sky130_fd_sc_hd__buf_1 wire5549 (.A(net5550),
    .X(net5549));
 sky130_fd_sc_hd__buf_1 wire5550 (.A(net5551),
    .X(net5550));
 sky130_fd_sc_hd__buf_1 wire5551 (.A(net5548),
    .X(net5551));
 sky130_fd_sc_hd__buf_1 wire5552 (.A(net5553),
    .X(net5552));
 sky130_fd_sc_hd__buf_1 max_length5553 (.A(net5548),
    .X(net5553));
 sky130_fd_sc_hd__clkbuf_1 wire5554 (.A(net5555),
    .X(net5554));
 sky130_fd_sc_hd__clkbuf_1 wire5555 (.A(\pid_d.mult0.a[6] ),
    .X(net5555));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout5556 (.A(net5569),
    .X(net5556));
 sky130_fd_sc_hd__buf_1 wire5557 (.A(net5559),
    .X(net5557));
 sky130_fd_sc_hd__buf_1 max_length5558 (.A(net5559),
    .X(net5558));
 sky130_fd_sc_hd__buf_1 wire5559 (.A(net5562),
    .X(net5559));
 sky130_fd_sc_hd__clkbuf_1 wire5560 (.A(net5561),
    .X(net5560));
 sky130_fd_sc_hd__clkbuf_1 wire5561 (.A(net5562),
    .X(net5561));
 sky130_fd_sc_hd__buf_1 wire5562 (.A(net5556),
    .X(net5562));
 sky130_fd_sc_hd__clkbuf_1 fanout5563 (.A(net5568),
    .X(net5563));
 sky130_fd_sc_hd__buf_1 wire5564 (.A(net5567),
    .X(net5564));
 sky130_fd_sc_hd__buf_1 wire5565 (.A(net5566),
    .X(net5565));
 sky130_fd_sc_hd__buf_1 wire5566 (.A(net5567),
    .X(net5566));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5567 (.A(net5563),
    .X(net5567));
 sky130_fd_sc_hd__clkbuf_1 fanout5568 (.A(\pid_d.mult0.a[5] ),
    .X(net5568));
 sky130_fd_sc_hd__clkbuf_1 wire5569 (.A(net5574),
    .X(net5569));
 sky130_fd_sc_hd__buf_1 wire5570 (.A(net5571),
    .X(net5570));
 sky130_fd_sc_hd__clkbuf_1 wire5571 (.A(net5572),
    .X(net5571));
 sky130_fd_sc_hd__buf_1 wire5572 (.A(net5573),
    .X(net5572));
 sky130_fd_sc_hd__clkbuf_1 wire5573 (.A(net5574),
    .X(net5573));
 sky130_fd_sc_hd__buf_1 wire5574 (.A(net5568),
    .X(net5574));
 sky130_fd_sc_hd__buf_1 fanout5575 (.A(net5587),
    .X(net5575));
 sky130_fd_sc_hd__clkbuf_1 wire5576 (.A(net5577),
    .X(net5576));
 sky130_fd_sc_hd__buf_1 wire5577 (.A(net5578),
    .X(net5577));
 sky130_fd_sc_hd__buf_1 wire5578 (.A(net5579),
    .X(net5578));
 sky130_fd_sc_hd__buf_1 wire5579 (.A(net5575),
    .X(net5579));
 sky130_fd_sc_hd__clkbuf_1 fanout5580 (.A(net5586),
    .X(net5580));
 sky130_fd_sc_hd__buf_1 wire5581 (.A(net5584),
    .X(net5581));
 sky130_fd_sc_hd__clkbuf_1 wire5582 (.A(net5583),
    .X(net5582));
 sky130_fd_sc_hd__buf_1 wire5583 (.A(net5584),
    .X(net5583));
 sky130_fd_sc_hd__buf_1 wire5584 (.A(net5585),
    .X(net5584));
 sky130_fd_sc_hd__buf_1 max_length5585 (.A(net5580),
    .X(net5585));
 sky130_fd_sc_hd__buf_1 fanout5586 (.A(\pid_d.mult0.a[4] ),
    .X(net5586));
 sky130_fd_sc_hd__clkbuf_1 wire5587 (.A(net5588),
    .X(net5587));
 sky130_fd_sc_hd__clkbuf_1 wire5588 (.A(net5589),
    .X(net5588));
 sky130_fd_sc_hd__clkbuf_1 wire5589 (.A(net5586),
    .X(net5589));
 sky130_fd_sc_hd__clkbuf_1 wire5590 (.A(net5591),
    .X(net5590));
 sky130_fd_sc_hd__clkbuf_1 wire5591 (.A(net5592),
    .X(net5591));
 sky130_fd_sc_hd__buf_1 wire5592 (.A(net5593),
    .X(net5592));
 sky130_fd_sc_hd__buf_1 wire5593 (.A(net5594),
    .X(net5593));
 sky130_fd_sc_hd__clkbuf_1 wire5594 (.A(net5586),
    .X(net5594));
 sky130_fd_sc_hd__clkbuf_1 fanout5595 (.A(net5604),
    .X(net5595));
 sky130_fd_sc_hd__buf_1 max_length5596 (.A(net5597),
    .X(net5596));
 sky130_fd_sc_hd__buf_1 wire5597 (.A(net5598),
    .X(net5597));
 sky130_fd_sc_hd__buf_1 wire5598 (.A(net5599),
    .X(net5598));
 sky130_fd_sc_hd__buf_1 wire5599 (.A(net5595),
    .X(net5599));
 sky130_fd_sc_hd__clkbuf_1 fanout5600 (.A(\pid_d.mult0.a[3] ),
    .X(net5600));
 sky130_fd_sc_hd__buf_1 wire5601 (.A(net5602),
    .X(net5601));
 sky130_fd_sc_hd__buf_1 wire5602 (.A(net5606),
    .X(net5602));
 sky130_fd_sc_hd__buf_1 wire5603 (.A(net5605),
    .X(net5603));
 sky130_fd_sc_hd__clkbuf_1 wire5604 (.A(net5605),
    .X(net5604));
 sky130_fd_sc_hd__buf_1 wire5605 (.A(net5607),
    .X(net5605));
 sky130_fd_sc_hd__buf_1 max_length5606 (.A(net5607),
    .X(net5606));
 sky130_fd_sc_hd__buf_1 wire5607 (.A(net5600),
    .X(net5607));
 sky130_fd_sc_hd__clkbuf_1 wire5608 (.A(net5609),
    .X(net5608));
 sky130_fd_sc_hd__buf_1 wire5609 (.A(net5610),
    .X(net5609));
 sky130_fd_sc_hd__clkbuf_1 max_length5610 (.A(\pid_d.mult0.a[3] ),
    .X(net5610));
 sky130_fd_sc_hd__buf_1 fanout5611 (.A(net5616),
    .X(net5611));
 sky130_fd_sc_hd__buf_1 max_length5612 (.A(net5613),
    .X(net5612));
 sky130_fd_sc_hd__clkbuf_2 wire5613 (.A(net5611),
    .X(net5613));
 sky130_fd_sc_hd__clkbuf_1 fanout5614 (.A(net5619),
    .X(net5614));
 sky130_fd_sc_hd__buf_1 wire5615 (.A(net5616),
    .X(net5615));
 sky130_fd_sc_hd__buf_1 wire5616 (.A(net5614),
    .X(net5616));
 sky130_fd_sc_hd__buf_1 fanout5617 (.A(net5623),
    .X(net5617));
 sky130_fd_sc_hd__buf_1 wire5618 (.A(net5619),
    .X(net5618));
 sky130_fd_sc_hd__buf_1 max_length5619 (.A(net5617),
    .X(net5619));
 sky130_fd_sc_hd__buf_1 fanout5620 (.A(\pid_d.mult0.a[2] ),
    .X(net5620));
 sky130_fd_sc_hd__buf_1 wire5621 (.A(net5622),
    .X(net5621));
 sky130_fd_sc_hd__clkbuf_1 wire5622 (.A(net5620),
    .X(net5622));
 sky130_fd_sc_hd__clkbuf_1 wire5623 (.A(net5624),
    .X(net5623));
 sky130_fd_sc_hd__clkbuf_1 wire5624 (.A(net5620),
    .X(net5624));
 sky130_fd_sc_hd__buf_1 fanout5625 (.A(net5629),
    .X(net5625));
 sky130_fd_sc_hd__clkbuf_2 wire5626 (.A(net5625),
    .X(net5626));
 sky130_fd_sc_hd__buf_1 wire5627 (.A(net5625),
    .X(net5627));
 sky130_fd_sc_hd__buf_1 fanout5628 (.A(net5632),
    .X(net5628));
 sky130_fd_sc_hd__buf_1 wire5629 (.A(net5628),
    .X(net5629));
 sky130_fd_sc_hd__buf_1 fanout5630 (.A(\pid_d.mult0.a[1] ),
    .X(net5630));
 sky130_fd_sc_hd__buf_1 wire5631 (.A(net5630),
    .X(net5631));
 sky130_fd_sc_hd__clkbuf_1 wire5632 (.A(net5633),
    .X(net5632));
 sky130_fd_sc_hd__clkbuf_1 wire5633 (.A(net5630),
    .X(net5633));
 sky130_fd_sc_hd__buf_1 fanout5634 (.A(net5636),
    .X(net5634));
 sky130_fd_sc_hd__clkbuf_2 wire5635 (.A(net5634),
    .X(net5635));
 sky130_fd_sc_hd__buf_1 fanout5636 (.A(net5643),
    .X(net5636));
 sky130_fd_sc_hd__buf_1 wire5637 (.A(net5638),
    .X(net5637));
 sky130_fd_sc_hd__clkbuf_2 wire5638 (.A(net5636),
    .X(net5638));
 sky130_fd_sc_hd__buf_1 fanout5639 (.A(\pid_d.mult0.a[0] ),
    .X(net5639));
 sky130_fd_sc_hd__clkbuf_1 wire5640 (.A(net5644),
    .X(net5640));
 sky130_fd_sc_hd__buf_1 max_length5641 (.A(net5643),
    .X(net5641));
 sky130_fd_sc_hd__buf_1 wire5642 (.A(net5643),
    .X(net5642));
 sky130_fd_sc_hd__buf_1 wire5643 (.A(net5639),
    .X(net5643));
 sky130_fd_sc_hd__buf_1 max_length5644 (.A(net5639),
    .X(net5644));
 sky130_fd_sc_hd__buf_1 fanout5645 (.A(net5663),
    .X(net5645));
 sky130_fd_sc_hd__buf_1 wire5646 (.A(net5647),
    .X(net5646));
 sky130_fd_sc_hd__clkbuf_2 wire5647 (.A(net5648),
    .X(net5647));
 sky130_fd_sc_hd__clkbuf_1 wire5648 (.A(net5649),
    .X(net5648));
 sky130_fd_sc_hd__buf_1 wire5649 (.A(net5645),
    .X(net5649));
 sky130_fd_sc_hd__clkbuf_1 fanout5650 (.A(\pid_d.mult0.b[15] ),
    .X(net5650));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5651 (.A(net5652),
    .X(net5651));
 sky130_fd_sc_hd__clkbuf_1 wire5652 (.A(net5656),
    .X(net5652));
 sky130_fd_sc_hd__buf_1 wire5653 (.A(net5654),
    .X(net5653));
 sky130_fd_sc_hd__clkbuf_2 wire5654 (.A(net5655),
    .X(net5654));
 sky130_fd_sc_hd__clkbuf_1 wire5655 (.A(net5657),
    .X(net5655));
 sky130_fd_sc_hd__clkbuf_1 max_length5656 (.A(net5657),
    .X(net5656));
 sky130_fd_sc_hd__buf_1 wire5657 (.A(net5650),
    .X(net5657));
 sky130_fd_sc_hd__clkbuf_1 wire5658 (.A(net5659),
    .X(net5658));
 sky130_fd_sc_hd__clkbuf_1 wire5659 (.A(net5660),
    .X(net5659));
 sky130_fd_sc_hd__clkbuf_1 wire5660 (.A(net5661),
    .X(net5660));
 sky130_fd_sc_hd__buf_1 wire5661 (.A(net5662),
    .X(net5661));
 sky130_fd_sc_hd__clkbuf_1 wire5662 (.A(net5663),
    .X(net5662));
 sky130_fd_sc_hd__buf_1 wire5663 (.A(net5664),
    .X(net5663));
 sky130_fd_sc_hd__clkbuf_1 wire5664 (.A(net5665),
    .X(net5664));
 sky130_fd_sc_hd__clkbuf_1 wire5665 (.A(net5666),
    .X(net5665));
 sky130_fd_sc_hd__clkbuf_1 wire5666 (.A(net5667),
    .X(net5666));
 sky130_fd_sc_hd__clkbuf_1 wire5667 (.A(net5668),
    .X(net5667));
 sky130_fd_sc_hd__clkbuf_1 wire5668 (.A(\pid_d.mult0.b[15] ),
    .X(net5668));
 sky130_fd_sc_hd__buf_1 fanout5669 (.A(net5678),
    .X(net5669));
 sky130_fd_sc_hd__buf_1 wire5670 (.A(net5671),
    .X(net5670));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length5671 (.A(net5672),
    .X(net5671));
 sky130_fd_sc_hd__buf_1 wire5672 (.A(net5669),
    .X(net5672));
 sky130_fd_sc_hd__buf_1 fanout5673 (.A(net5681),
    .X(net5673));
 sky130_fd_sc_hd__buf_1 max_length5674 (.A(net5673),
    .X(net5674));
 sky130_fd_sc_hd__clkbuf_1 wire5675 (.A(net5676),
    .X(net5675));
 sky130_fd_sc_hd__buf_1 wire5676 (.A(net5677),
    .X(net5676));
 sky130_fd_sc_hd__clkbuf_1 wire5677 (.A(net5678),
    .X(net5677));
 sky130_fd_sc_hd__buf_1 wire5678 (.A(net5679),
    .X(net5678));
 sky130_fd_sc_hd__buf_1 wire5679 (.A(net5680),
    .X(net5679));
 sky130_fd_sc_hd__buf_1 wire5680 (.A(net5673),
    .X(net5680));
 sky130_fd_sc_hd__clkbuf_1 wire5681 (.A(net5682),
    .X(net5681));
 sky130_fd_sc_hd__clkbuf_1 wire5682 (.A(net5683),
    .X(net5682));
 sky130_fd_sc_hd__clkbuf_1 wire5683 (.A(net5684),
    .X(net5683));
 sky130_fd_sc_hd__clkbuf_1 wire5684 (.A(\pid_d.mult0.b[14] ),
    .X(net5684));
 sky130_fd_sc_hd__buf_1 fanout5685 (.A(net5697),
    .X(net5685));
 sky130_fd_sc_hd__buf_1 wire5686 (.A(net5688),
    .X(net5686));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5687 (.A(net5685),
    .X(net5687));
 sky130_fd_sc_hd__buf_1 max_length5688 (.A(net5685),
    .X(net5688));
 sky130_fd_sc_hd__buf_1 fanout5689 (.A(net5695),
    .X(net5689));
 sky130_fd_sc_hd__clkbuf_1 wire5690 (.A(net5691),
    .X(net5690));
 sky130_fd_sc_hd__buf_1 wire5691 (.A(net5692),
    .X(net5691));
 sky130_fd_sc_hd__buf_1 wire5692 (.A(net5694),
    .X(net5692));
 sky130_fd_sc_hd__buf_1 wire5693 (.A(net5689),
    .X(net5693));
 sky130_fd_sc_hd__buf_1 max_length5694 (.A(net5689),
    .X(net5694));
 sky130_fd_sc_hd__clkbuf_1 wire5695 (.A(net5696),
    .X(net5695));
 sky130_fd_sc_hd__clkbuf_1 wire5696 (.A(net5697),
    .X(net5696));
 sky130_fd_sc_hd__buf_1 wire5697 (.A(net5698),
    .X(net5697));
 sky130_fd_sc_hd__clkbuf_1 wire5698 (.A(net5699),
    .X(net5698));
 sky130_fd_sc_hd__clkbuf_1 wire5699 (.A(net5700),
    .X(net5699));
 sky130_fd_sc_hd__clkbuf_1 wire5700 (.A(\pid_d.mult0.b[13] ),
    .X(net5700));
 sky130_fd_sc_hd__buf_1 fanout5701 (.A(net5716),
    .X(net5701));
 sky130_fd_sc_hd__buf_1 wire5702 (.A(net5705),
    .X(net5702));
 sky130_fd_sc_hd__buf_1 wire5703 (.A(net5704),
    .X(net5703));
 sky130_fd_sc_hd__buf_1 wire5704 (.A(net5701),
    .X(net5704));
 sky130_fd_sc_hd__buf_1 max_length5705 (.A(net5701),
    .X(net5705));
 sky130_fd_sc_hd__clkbuf_1 fanout5706 (.A(net5715),
    .X(net5706));
 sky130_fd_sc_hd__buf_1 wire5707 (.A(net5708),
    .X(net5707));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5708 (.A(net5709),
    .X(net5708));
 sky130_fd_sc_hd__buf_1 wire5709 (.A(net5710),
    .X(net5709));
 sky130_fd_sc_hd__buf_1 wire5710 (.A(net5711),
    .X(net5710));
 sky130_fd_sc_hd__buf_1 wire5711 (.A(net5706),
    .X(net5711));
 sky130_fd_sc_hd__buf_1 fanout5712 (.A(\pid_d.mult0.b[12] ),
    .X(net5712));
 sky130_fd_sc_hd__clkbuf_1 wire5713 (.A(net5714),
    .X(net5713));
 sky130_fd_sc_hd__clkbuf_1 wire5714 (.A(net5715),
    .X(net5714));
 sky130_fd_sc_hd__buf_1 wire5715 (.A(net5716),
    .X(net5715));
 sky130_fd_sc_hd__buf_1 wire5716 (.A(net5717),
    .X(net5716));
 sky130_fd_sc_hd__clkbuf_1 wire5717 (.A(net5712),
    .X(net5717));
 sky130_fd_sc_hd__buf_1 fanout5718 (.A(net5734),
    .X(net5718));
 sky130_fd_sc_hd__buf_1 wire5719 (.A(net5718),
    .X(net5719));
 sky130_fd_sc_hd__buf_1 wire5720 (.A(net5721),
    .X(net5720));
 sky130_fd_sc_hd__buf_1 wire5721 (.A(net5723),
    .X(net5721));
 sky130_fd_sc_hd__clkbuf_1 wire5722 (.A(net5723),
    .X(net5722));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5723 (.A(net5718),
    .X(net5723));
 sky130_fd_sc_hd__buf_1 fanout5724 (.A(net5735),
    .X(net5724));
 sky130_fd_sc_hd__clkbuf_1 wire5725 (.A(net5729),
    .X(net5725));
 sky130_fd_sc_hd__clkbuf_1 wire5726 (.A(net5727),
    .X(net5726));
 sky130_fd_sc_hd__clkbuf_1 wire5727 (.A(net5728),
    .X(net5727));
 sky130_fd_sc_hd__clkbuf_1 wire5728 (.A(net5729),
    .X(net5728));
 sky130_fd_sc_hd__buf_1 wire5729 (.A(net5724),
    .X(net5729));
 sky130_fd_sc_hd__buf_1 wire5730 (.A(net5731),
    .X(net5730));
 sky130_fd_sc_hd__buf_1 wire5731 (.A(net5724),
    .X(net5731));
 sky130_fd_sc_hd__clkbuf_1 wire5732 (.A(net5733),
    .X(net5732));
 sky130_fd_sc_hd__clkbuf_1 wire5733 (.A(net5734),
    .X(net5733));
 sky130_fd_sc_hd__buf_1 wire5734 (.A(net5735),
    .X(net5734));
 sky130_fd_sc_hd__buf_1 wire5735 (.A(net5736),
    .X(net5735));
 sky130_fd_sc_hd__clkbuf_1 wire5736 (.A(net5737),
    .X(net5736));
 sky130_fd_sc_hd__clkbuf_1 wire5737 (.A(net5738),
    .X(net5737));
 sky130_fd_sc_hd__clkbuf_1 wire5738 (.A(\pid_d.mult0.b[11] ),
    .X(net5738));
 sky130_fd_sc_hd__buf_1 fanout5739 (.A(net5756),
    .X(net5739));
 sky130_fd_sc_hd__buf_1 wire5740 (.A(net5741),
    .X(net5740));
 sky130_fd_sc_hd__buf_1 wire5741 (.A(net5739),
    .X(net5741));
 sky130_fd_sc_hd__clkbuf_1 wire5742 (.A(net5743),
    .X(net5742));
 sky130_fd_sc_hd__buf_1 wire5743 (.A(net5739),
    .X(net5743));
 sky130_fd_sc_hd__buf_1 fanout5744 (.A(net5754),
    .X(net5744));
 sky130_fd_sc_hd__buf_1 wire5745 (.A(net5746),
    .X(net5745));
 sky130_fd_sc_hd__buf_1 wire5746 (.A(net5749),
    .X(net5746));
 sky130_fd_sc_hd__buf_1 wire5747 (.A(net5748),
    .X(net5747));
 sky130_fd_sc_hd__clkbuf_1 wire5748 (.A(net5749),
    .X(net5748));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5749 (.A(net5744),
    .X(net5749));
 sky130_fd_sc_hd__buf_1 wire5750 (.A(net5744),
    .X(net5750));
 sky130_fd_sc_hd__buf_1 fanout5751 (.A(\pid_d.mult0.b[10] ),
    .X(net5751));
 sky130_fd_sc_hd__clkbuf_1 wire5752 (.A(net5753),
    .X(net5752));
 sky130_fd_sc_hd__buf_1 wire5753 (.A(net5754),
    .X(net5753));
 sky130_fd_sc_hd__buf_1 wire5754 (.A(net5755),
    .X(net5754));
 sky130_fd_sc_hd__clkbuf_1 wire5755 (.A(net5756),
    .X(net5755));
 sky130_fd_sc_hd__buf_1 wire5756 (.A(net5757),
    .X(net5756));
 sky130_fd_sc_hd__clkbuf_1 wire5757 (.A(net5751),
    .X(net5757));
 sky130_fd_sc_hd__clkbuf_1 fanout5758 (.A(net5766),
    .X(net5758));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length5759 (.A(net5760),
    .X(net5759));
 sky130_fd_sc_hd__buf_1 wire5760 (.A(net5761),
    .X(net5760));
 sky130_fd_sc_hd__buf_1 wire5761 (.A(net5758),
    .X(net5761));
 sky130_fd_sc_hd__clkbuf_2 fanout5762 (.A(net5765),
    .X(net5762));
 sky130_fd_sc_hd__buf_1 wire5763 (.A(net5764),
    .X(net5763));
 sky130_fd_sc_hd__buf_1 wire5764 (.A(net5762),
    .X(net5764));
 sky130_fd_sc_hd__buf_1 fanout5765 (.A(net5767),
    .X(net5765));
 sky130_fd_sc_hd__buf_1 fanout5766 (.A(net5770),
    .X(net5766));
 sky130_fd_sc_hd__clkbuf_1 wire5767 (.A(net5768),
    .X(net5767));
 sky130_fd_sc_hd__buf_1 wire5768 (.A(net5769),
    .X(net5768));
 sky130_fd_sc_hd__buf_1 wire5769 (.A(net5766),
    .X(net5769));
 sky130_fd_sc_hd__clkbuf_1 wire5770 (.A(net5771),
    .X(net5770));
 sky130_fd_sc_hd__clkbuf_1 wire5771 (.A(net5772),
    .X(net5771));
 sky130_fd_sc_hd__clkbuf_1 wire5772 (.A(net5773),
    .X(net5772));
 sky130_fd_sc_hd__clkbuf_1 wire5773 (.A(\pid_d.mult0.b[9] ),
    .X(net5773));
 sky130_fd_sc_hd__buf_1 fanout5774 (.A(net5778),
    .X(net5774));
 sky130_fd_sc_hd__buf_1 max_length5775 (.A(net5776),
    .X(net5775));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5776 (.A(net5774),
    .X(net5776));
 sky130_fd_sc_hd__buf_1 fanout5777 (.A(net5788),
    .X(net5777));
 sky130_fd_sc_hd__buf_1 wire5778 (.A(net5777),
    .X(net5778));
 sky130_fd_sc_hd__buf_1 wire5779 (.A(net5780),
    .X(net5779));
 sky130_fd_sc_hd__buf_1 wire5780 (.A(net5781),
    .X(net5780));
 sky130_fd_sc_hd__clkbuf_1 wire5781 (.A(net5782),
    .X(net5781));
 sky130_fd_sc_hd__buf_1 wire5782 (.A(net5777),
    .X(net5782));
 sky130_fd_sc_hd__buf_1 fanout5783 (.A(net5786),
    .X(net5783));
 sky130_fd_sc_hd__buf_1 wire5784 (.A(net5785),
    .X(net5784));
 sky130_fd_sc_hd__buf_1 wire5785 (.A(net5783),
    .X(net5785));
 sky130_fd_sc_hd__clkbuf_1 wire5786 (.A(net5787),
    .X(net5786));
 sky130_fd_sc_hd__clkbuf_1 wire5787 (.A(net5788),
    .X(net5787));
 sky130_fd_sc_hd__buf_1 wire5788 (.A(net5789),
    .X(net5788));
 sky130_fd_sc_hd__clkbuf_1 wire5789 (.A(net5790),
    .X(net5789));
 sky130_fd_sc_hd__clkbuf_1 wire5790 (.A(net5791),
    .X(net5790));
 sky130_fd_sc_hd__clkbuf_1 wire5791 (.A(\pid_d.mult0.b[8] ),
    .X(net5791));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout5792 (.A(net5797),
    .X(net5792));
 sky130_fd_sc_hd__buf_1 wire5793 (.A(net5792),
    .X(net5793));
 sky130_fd_sc_hd__buf_1 wire5794 (.A(net5792),
    .X(net5794));
 sky130_fd_sc_hd__buf_1 fanout5795 (.A(net5803),
    .X(net5795));
 sky130_fd_sc_hd__clkbuf_1 wire5796 (.A(net5797),
    .X(net5796));
 sky130_fd_sc_hd__buf_1 wire5797 (.A(net5795),
    .X(net5797));
 sky130_fd_sc_hd__clkbuf_1 fanout5798 (.A(net5805),
    .X(net5798));
 sky130_fd_sc_hd__clkbuf_2 wire5799 (.A(net5801),
    .X(net5799));
 sky130_fd_sc_hd__buf_1 max_length5800 (.A(net5801),
    .X(net5800));
 sky130_fd_sc_hd__buf_1 wire5801 (.A(net5798),
    .X(net5801));
 sky130_fd_sc_hd__buf_1 fanout5802 (.A(\pid_d.mult0.b[7] ),
    .X(net5802));
 sky130_fd_sc_hd__buf_1 wire5803 (.A(net5807),
    .X(net5803));
 sky130_fd_sc_hd__clkbuf_1 wire5804 (.A(net5805),
    .X(net5804));
 sky130_fd_sc_hd__buf_1 wire5805 (.A(net5806),
    .X(net5805));
 sky130_fd_sc_hd__buf_1 wire5806 (.A(net5807),
    .X(net5806));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5807 (.A(net5808),
    .X(net5807));
 sky130_fd_sc_hd__clkbuf_1 wire5808 (.A(net5802),
    .X(net5808));
 sky130_fd_sc_hd__buf_1 fanout5809 (.A(net5829),
    .X(net5809));
 sky130_fd_sc_hd__buf_1 wire5810 (.A(net5811),
    .X(net5810));
 sky130_fd_sc_hd__buf_1 wire5811 (.A(net5815),
    .X(net5811));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5812 (.A(net5813),
    .X(net5812));
 sky130_fd_sc_hd__buf_1 wire5813 (.A(net5814),
    .X(net5813));
 sky130_fd_sc_hd__buf_1 wire5814 (.A(net5815),
    .X(net5814));
 sky130_fd_sc_hd__buf_1 wire5815 (.A(net5809),
    .X(net5815));
 sky130_fd_sc_hd__buf_1 fanout5816 (.A(net5819),
    .X(net5816));
 sky130_fd_sc_hd__buf_1 wire5817 (.A(net5818),
    .X(net5817));
 sky130_fd_sc_hd__clkbuf_1 wire5818 (.A(net5816),
    .X(net5818));
 sky130_fd_sc_hd__buf_1 fanout5819 (.A(net5827),
    .X(net5819));
 sky130_fd_sc_hd__buf_1 wire5820 (.A(net5821),
    .X(net5820));
 sky130_fd_sc_hd__clkbuf_2 wire5821 (.A(net5822),
    .X(net5821));
 sky130_fd_sc_hd__buf_1 wire5822 (.A(net5823),
    .X(net5822));
 sky130_fd_sc_hd__buf_1 wire5823 (.A(net5824),
    .X(net5823));
 sky130_fd_sc_hd__clkbuf_1 wire5824 (.A(net5825),
    .X(net5824));
 sky130_fd_sc_hd__clkbuf_1 wire5825 (.A(net5826),
    .X(net5825));
 sky130_fd_sc_hd__clkbuf_1 wire5826 (.A(net5819),
    .X(net5826));
 sky130_fd_sc_hd__clkbuf_1 wire5827 (.A(net5828),
    .X(net5827));
 sky130_fd_sc_hd__clkbuf_1 wire5828 (.A(net5829),
    .X(net5828));
 sky130_fd_sc_hd__buf_1 wire5829 (.A(\pid_d.mult0.b[6] ),
    .X(net5829));
 sky130_fd_sc_hd__buf_1 fanout5830 (.A(net5847),
    .X(net5830));
 sky130_fd_sc_hd__buf_1 wire5831 (.A(net5832),
    .X(net5831));
 sky130_fd_sc_hd__buf_1 wire5832 (.A(net5836),
    .X(net5832));
 sky130_fd_sc_hd__clkbuf_1 wire5833 (.A(net5834),
    .X(net5833));
 sky130_fd_sc_hd__clkbuf_1 wire5834 (.A(net5835),
    .X(net5834));
 sky130_fd_sc_hd__clkbuf_1 wire5835 (.A(net5837),
    .X(net5835));
 sky130_fd_sc_hd__buf_1 max_length5836 (.A(net5837),
    .X(net5836));
 sky130_fd_sc_hd__buf_1 wire5837 (.A(net5838),
    .X(net5837));
 sky130_fd_sc_hd__buf_1 wire5838 (.A(net5830),
    .X(net5838));
 sky130_fd_sc_hd__clkbuf_2 fanout5839 (.A(net5848),
    .X(net5839));
 sky130_fd_sc_hd__buf_1 fanout5840 (.A(\pid_d.mult0.b[5] ),
    .X(net5840));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5841 (.A(net5842),
    .X(net5841));
 sky130_fd_sc_hd__buf_1 wire5842 (.A(net5843),
    .X(net5842));
 sky130_fd_sc_hd__buf_1 wire5843 (.A(net5844),
    .X(net5843));
 sky130_fd_sc_hd__buf_1 wire5844 (.A(net5845),
    .X(net5844));
 sky130_fd_sc_hd__clkbuf_1 wire5845 (.A(net5846),
    .X(net5845));
 sky130_fd_sc_hd__clkbuf_1 wire5846 (.A(net5840),
    .X(net5846));
 sky130_fd_sc_hd__clkbuf_1 wire5847 (.A(net5853),
    .X(net5847));
 sky130_fd_sc_hd__clkbuf_1 wire5848 (.A(net5849),
    .X(net5848));
 sky130_fd_sc_hd__clkbuf_1 wire5849 (.A(net5850),
    .X(net5849));
 sky130_fd_sc_hd__clkbuf_1 wire5850 (.A(net5851),
    .X(net5850));
 sky130_fd_sc_hd__buf_1 wire5851 (.A(net5852),
    .X(net5851));
 sky130_fd_sc_hd__clkbuf_1 max_length5852 (.A(net5853),
    .X(net5852));
 sky130_fd_sc_hd__buf_1 wire5853 (.A(net5854),
    .X(net5853));
 sky130_fd_sc_hd__clkbuf_1 wire5854 (.A(net5855),
    .X(net5854));
 sky130_fd_sc_hd__clkbuf_1 wire5855 (.A(\pid_d.mult0.b[5] ),
    .X(net5855));
 sky130_fd_sc_hd__buf_1 fanout5856 (.A(net5864),
    .X(net5856));
 sky130_fd_sc_hd__buf_1 wire5857 (.A(net5858),
    .X(net5857));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5858 (.A(net5859),
    .X(net5858));
 sky130_fd_sc_hd__buf_1 wire5859 (.A(net5856),
    .X(net5859));
 sky130_fd_sc_hd__clkbuf_1 fanout5860 (.A(\pid_d.mult0.b[4] ),
    .X(net5860));
 sky130_fd_sc_hd__buf_1 wire5861 (.A(net5865),
    .X(net5861));
 sky130_fd_sc_hd__buf_1 wire5862 (.A(net5863),
    .X(net5862));
 sky130_fd_sc_hd__clkbuf_1 wire5863 (.A(net5864),
    .X(net5863));
 sky130_fd_sc_hd__buf_1 wire5864 (.A(net5865),
    .X(net5864));
 sky130_fd_sc_hd__buf_1 wire5865 (.A(net5866),
    .X(net5865));
 sky130_fd_sc_hd__clkbuf_1 wire5866 (.A(net5860),
    .X(net5866));
 sky130_fd_sc_hd__buf_1 fanout5867 (.A(net5875),
    .X(net5867));
 sky130_fd_sc_hd__buf_1 wire5868 (.A(net5869),
    .X(net5868));
 sky130_fd_sc_hd__buf_1 wire5869 (.A(net5873),
    .X(net5869));
 sky130_fd_sc_hd__clkbuf_1 wire5870 (.A(net5871),
    .X(net5870));
 sky130_fd_sc_hd__clkbuf_1 wire5871 (.A(net5872),
    .X(net5871));
 sky130_fd_sc_hd__buf_1 wire5872 (.A(net5874),
    .X(net5872));
 sky130_fd_sc_hd__buf_1 max_length5873 (.A(net5874),
    .X(net5873));
 sky130_fd_sc_hd__buf_1 wire5874 (.A(net5867),
    .X(net5874));
 sky130_fd_sc_hd__clkbuf_1 wire5875 (.A(net5876),
    .X(net5875));
 sky130_fd_sc_hd__clkbuf_1 wire5876 (.A(net5877),
    .X(net5876));
 sky130_fd_sc_hd__clkbuf_1 wire5877 (.A(\pid_d.mult0.b[4] ),
    .X(net5877));
 sky130_fd_sc_hd__buf_1 fanout5878 (.A(net5885),
    .X(net5878));
 sky130_fd_sc_hd__buf_1 wire5879 (.A(net5880),
    .X(net5879));
 sky130_fd_sc_hd__buf_1 wire5880 (.A(net5881),
    .X(net5880));
 sky130_fd_sc_hd__buf_1 wire5881 (.A(net5878),
    .X(net5881));
 sky130_fd_sc_hd__buf_1 fanout5882 (.A(net5885),
    .X(net5882));
 sky130_fd_sc_hd__clkbuf_2 fanout5883 (.A(net5899),
    .X(net5883));
 sky130_fd_sc_hd__buf_1 wire5884 (.A(net5883),
    .X(net5884));
 sky130_fd_sc_hd__clkbuf_1 wire5885 (.A(net5886),
    .X(net5885));
 sky130_fd_sc_hd__clkbuf_1 wire5886 (.A(net5887),
    .X(net5886));
 sky130_fd_sc_hd__clkbuf_1 max_length5887 (.A(net5883),
    .X(net5887));
 sky130_fd_sc_hd__clkbuf_1 fanout5888 (.A(net5895),
    .X(net5888));
 sky130_fd_sc_hd__clkbuf_1 wire5889 (.A(net5890),
    .X(net5889));
 sky130_fd_sc_hd__buf_1 wire5890 (.A(net5894),
    .X(net5890));
 sky130_fd_sc_hd__clkbuf_1 wire5891 (.A(net5892),
    .X(net5891));
 sky130_fd_sc_hd__buf_1 wire5892 (.A(net5893),
    .X(net5892));
 sky130_fd_sc_hd__buf_1 max_length5893 (.A(net5894),
    .X(net5893));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5894 (.A(net5888),
    .X(net5894));
 sky130_fd_sc_hd__buf_1 fanout5895 (.A(\pid_d.mult0.b[3] ),
    .X(net5895));
 sky130_fd_sc_hd__buf_1 wire5896 (.A(net5897),
    .X(net5896));
 sky130_fd_sc_hd__buf_1 wire5897 (.A(net5898),
    .X(net5897));
 sky130_fd_sc_hd__clkbuf_1 wire5898 (.A(net5895),
    .X(net5898));
 sky130_fd_sc_hd__clkbuf_1 wire5899 (.A(net5900),
    .X(net5899));
 sky130_fd_sc_hd__clkbuf_1 wire5900 (.A(net5901),
    .X(net5900));
 sky130_fd_sc_hd__clkbuf_1 wire5901 (.A(net5902),
    .X(net5901));
 sky130_fd_sc_hd__clkbuf_1 wire5902 (.A(net5895),
    .X(net5902));
 sky130_fd_sc_hd__clkbuf_1 fanout5903 (.A(net5916),
    .X(net5903));
 sky130_fd_sc_hd__clkbuf_1 wire5904 (.A(net5903),
    .X(net5904));
 sky130_fd_sc_hd__buf_1 wire5905 (.A(net5906),
    .X(net5905));
 sky130_fd_sc_hd__clkbuf_2 wire5906 (.A(net5907),
    .X(net5906));
 sky130_fd_sc_hd__clkbuf_1 wire5907 (.A(net5908),
    .X(net5907));
 sky130_fd_sc_hd__buf_1 max_length5908 (.A(net5903),
    .X(net5908));
 sky130_fd_sc_hd__buf_1 fanout5909 (.A(net5912),
    .X(net5909));
 sky130_fd_sc_hd__buf_1 max_length5910 (.A(net5911),
    .X(net5910));
 sky130_fd_sc_hd__clkbuf_2 wire5911 (.A(net5909),
    .X(net5911));
 sky130_fd_sc_hd__buf_1 fanout5912 (.A(net5918),
    .X(net5912));
 sky130_fd_sc_hd__clkbuf_1 wire5913 (.A(net5914),
    .X(net5913));
 sky130_fd_sc_hd__buf_1 wire5914 (.A(net5915),
    .X(net5914));
 sky130_fd_sc_hd__clkbuf_1 wire5915 (.A(net5916),
    .X(net5915));
 sky130_fd_sc_hd__buf_1 wire5916 (.A(net5912),
    .X(net5916));
 sky130_fd_sc_hd__clkbuf_1 fanout5917 (.A(net5925),
    .X(net5917));
 sky130_fd_sc_hd__clkbuf_1 wire5918 (.A(net5919),
    .X(net5918));
 sky130_fd_sc_hd__clkbuf_1 wire5919 (.A(net5920),
    .X(net5919));
 sky130_fd_sc_hd__buf_1 wire5920 (.A(net5921),
    .X(net5920));
 sky130_fd_sc_hd__buf_1 wire5921 (.A(net5922),
    .X(net5921));
 sky130_fd_sc_hd__buf_1 wire5922 (.A(net5923),
    .X(net5922));
 sky130_fd_sc_hd__clkbuf_1 wire5923 (.A(net5924),
    .X(net5923));
 sky130_fd_sc_hd__buf_1 wire5924 (.A(net5917),
    .X(net5924));
 sky130_fd_sc_hd__clkbuf_1 wire5925 (.A(net5926),
    .X(net5925));
 sky130_fd_sc_hd__clkbuf_1 wire5926 (.A(net5927),
    .X(net5926));
 sky130_fd_sc_hd__clkbuf_1 wire5927 (.A(\pid_d.mult0.b[2] ),
    .X(net5927));
 sky130_fd_sc_hd__buf_1 fanout5928 (.A(net5933),
    .X(net5928));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5929 (.A(net5930),
    .X(net5929));
 sky130_fd_sc_hd__buf_1 wire5930 (.A(net5928),
    .X(net5930));
 sky130_fd_sc_hd__buf_1 fanout5931 (.A(net5938),
    .X(net5931));
 sky130_fd_sc_hd__clkbuf_1 max_length5932 (.A(net5933),
    .X(net5932));
 sky130_fd_sc_hd__buf_1 wire5933 (.A(net5934),
    .X(net5933));
 sky130_fd_sc_hd__clkbuf_1 wire5934 (.A(net5931),
    .X(net5934));
 sky130_fd_sc_hd__clkbuf_1 wire5935 (.A(net5931),
    .X(net5935));
 sky130_fd_sc_hd__buf_1 fanout5936 (.A(net5942),
    .X(net5936));
 sky130_fd_sc_hd__buf_1 wire5937 (.A(net5939),
    .X(net5937));
 sky130_fd_sc_hd__clkbuf_1 max_length5938 (.A(net5940),
    .X(net5938));
 sky130_fd_sc_hd__clkbuf_1 max_length5939 (.A(net5940),
    .X(net5939));
 sky130_fd_sc_hd__buf_1 wire5940 (.A(net5936),
    .X(net5940));
 sky130_fd_sc_hd__clkbuf_1 fanout5941 (.A(\pid_d.mult0.b[1] ),
    .X(net5941));
 sky130_fd_sc_hd__clkbuf_1 wire5942 (.A(net5945),
    .X(net5942));
 sky130_fd_sc_hd__buf_1 wire5943 (.A(net5944),
    .X(net5943));
 sky130_fd_sc_hd__buf_1 max_length5944 (.A(net5945),
    .X(net5944));
 sky130_fd_sc_hd__buf_1 wire5945 (.A(net5946),
    .X(net5945));
 sky130_fd_sc_hd__clkbuf_1 wire5946 (.A(net5947),
    .X(net5946));
 sky130_fd_sc_hd__clkbuf_1 wire5947 (.A(net5941),
    .X(net5947));
 sky130_fd_sc_hd__clkbuf_1 fanout5948 (.A(net5955),
    .X(net5948));
 sky130_fd_sc_hd__buf_1 wire5949 (.A(net5951),
    .X(net5949));
 sky130_fd_sc_hd__buf_1 wire5950 (.A(net5951),
    .X(net5950));
 sky130_fd_sc_hd__buf_1 wire5951 (.A(net5952),
    .X(net5951));
 sky130_fd_sc_hd__buf_1 max_length5952 (.A(net5948),
    .X(net5952));
 sky130_fd_sc_hd__buf_1 fanout5953 (.A(net5959),
    .X(net5953));
 sky130_fd_sc_hd__buf_1 wire5954 (.A(net5953),
    .X(net5954));
 sky130_fd_sc_hd__buf_1 wire5955 (.A(net5956),
    .X(net5955));
 sky130_fd_sc_hd__clkbuf_1 wire5956 (.A(net5957),
    .X(net5956));
 sky130_fd_sc_hd__clkbuf_1 wire5957 (.A(net5953),
    .X(net5957));
 sky130_fd_sc_hd__buf_1 fanout5958 (.A(\pid_d.mult0.b[0] ),
    .X(net5958));
 sky130_fd_sc_hd__clkbuf_1 wire5959 (.A(net5960),
    .X(net5959));
 sky130_fd_sc_hd__buf_1 wire5960 (.A(net5962),
    .X(net5960));
 sky130_fd_sc_hd__buf_1 wire5961 (.A(net5963),
    .X(net5961));
 sky130_fd_sc_hd__clkbuf_1 max_length5962 (.A(net5963),
    .X(net5962));
 sky130_fd_sc_hd__buf_1 wire5963 (.A(net5958),
    .X(net5963));
 sky130_fd_sc_hd__buf_1 wire5964 (.A(\pid_d.curr_error[15] ),
    .X(net5964));
 sky130_fd_sc_hd__buf_1 wire5965 (.A(\pid_d.curr_error[13] ),
    .X(net5965));
 sky130_fd_sc_hd__buf_1 wire5966 (.A(\pid_d.curr_error[11] ),
    .X(net5966));
 sky130_fd_sc_hd__buf_1 wire5967 (.A(\pid_d.curr_error[9] ),
    .X(net5967));
 sky130_fd_sc_hd__clkbuf_2 wire5968 (.A(\pid_d.curr_error[6] ),
    .X(net5968));
 sky130_fd_sc_hd__buf_1 wire5969 (.A(\pid_d.curr_error[5] ),
    .X(net5969));
 sky130_fd_sc_hd__buf_1 wire5970 (.A(\pid_d.curr_error[3] ),
    .X(net5970));
 sky130_fd_sc_hd__clkbuf_2 wire5971 (.A(\pid_d.curr_error[2] ),
    .X(net5971));
 sky130_fd_sc_hd__buf_1 wire5972 (.A(\pid_d.curr_error[1] ),
    .X(net5972));
 sky130_fd_sc_hd__clkbuf_2 wire5973 (.A(\pid_d.curr_error[0] ),
    .X(net5973));
 sky130_fd_sc_hd__buf_1 wire5974 (.A(\pid_d.curr_int[15] ),
    .X(net5974));
 sky130_fd_sc_hd__buf_1 wire5975 (.A(\pid_d.curr_int[12] ),
    .X(net5975));
 sky130_fd_sc_hd__clkbuf_2 wire5976 (.A(\pid_d.curr_int[9] ),
    .X(net5976));
 sky130_fd_sc_hd__clkbuf_2 wire5977 (.A(\pid_d.curr_int[8] ),
    .X(net5977));
 sky130_fd_sc_hd__clkbuf_2 wire5978 (.A(\pid_d.curr_int[7] ),
    .X(net5978));
 sky130_fd_sc_hd__buf_1 wire5979 (.A(\pid_d.curr_int[6] ),
    .X(net5979));
 sky130_fd_sc_hd__buf_1 wire5980 (.A(\pid_d.curr_int[5] ),
    .X(net5980));
 sky130_fd_sc_hd__clkbuf_2 wire5981 (.A(\pid_d.curr_int[4] ),
    .X(net5981));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5982 (.A(\pid_d.curr_int[3] ),
    .X(net5982));
 sky130_fd_sc_hd__clkbuf_2 wire5983 (.A(\pid_d.curr_int[2] ),
    .X(net5983));
 sky130_fd_sc_hd__clkbuf_2 wire5984 (.A(net5985),
    .X(net5984));
 sky130_fd_sc_hd__buf_1 max_length5985 (.A(\pid_d.curr_int[1] ),
    .X(net5985));
 sky130_fd_sc_hd__buf_1 wire5986 (.A(\pid_d.curr_int[0] ),
    .X(net5986));
 sky130_fd_sc_hd__clkbuf_2 max_length5987 (.A(\pid_d.curr_int[0] ),
    .X(net5987));
 sky130_fd_sc_hd__buf_1 fanout5988 (.A(net5991),
    .X(net5988));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire5989 (.A(net5990),
    .X(net5989));
 sky130_fd_sc_hd__buf_1 wire5990 (.A(net5988),
    .X(net5990));
 sky130_fd_sc_hd__clkbuf_1 fanout5991 (.A(net5997),
    .X(net5991));
 sky130_fd_sc_hd__buf_1 max_length5992 (.A(net5993),
    .X(net5992));
 sky130_fd_sc_hd__buf_1 wire5993 (.A(net5991),
    .X(net5993));
 sky130_fd_sc_hd__clkbuf_1 fanout5994 (.A(net6015),
    .X(net5994));
 sky130_fd_sc_hd__buf_1 wire5995 (.A(net5996),
    .X(net5995));
 sky130_fd_sc_hd__buf_1 wire5996 (.A(net5997),
    .X(net5996));
 sky130_fd_sc_hd__buf_1 wire5997 (.A(net5998),
    .X(net5997));
 sky130_fd_sc_hd__buf_1 wire5998 (.A(net5994),
    .X(net5998));
 sky130_fd_sc_hd__buf_1 fanout5999 (.A(net6003),
    .X(net5999));
 sky130_fd_sc_hd__buf_1 wire6000 (.A(net6001),
    .X(net6000));
 sky130_fd_sc_hd__buf_1 wire6001 (.A(net6002),
    .X(net6001));
 sky130_fd_sc_hd__buf_1 max_length6002 (.A(net5999),
    .X(net6002));
 sky130_fd_sc_hd__buf_1 fanout6003 (.A(net6014),
    .X(net6003));
 sky130_fd_sc_hd__buf_1 wire6004 (.A(net6006),
    .X(net6004));
 sky130_fd_sc_hd__buf_1 max_length6005 (.A(net6006),
    .X(net6005));
 sky130_fd_sc_hd__buf_1 wire6006 (.A(net6003),
    .X(net6006));
 sky130_fd_sc_hd__buf_1 fanout6007 (.A(net6011),
    .X(net6007));
 sky130_fd_sc_hd__buf_1 max_length6008 (.A(net6009),
    .X(net6008));
 sky130_fd_sc_hd__buf_1 wire6009 (.A(net6010),
    .X(net6009));
 sky130_fd_sc_hd__buf_1 wire6010 (.A(net6007),
    .X(net6010));
 sky130_fd_sc_hd__buf_1 fanout6011 (.A(net6017),
    .X(net6011));
 sky130_fd_sc_hd__clkbuf_2 wire6012 (.A(net6013),
    .X(net6012));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6013 (.A(net6011),
    .X(net6013));
 sky130_fd_sc_hd__buf_1 fanout6014 (.A(\cordic0.vec[0][17] ),
    .X(net6014));
 sky130_fd_sc_hd__clkbuf_1 wire6015 (.A(net6014),
    .X(net6015));
 sky130_fd_sc_hd__clkbuf_1 wire6016 (.A(net6017),
    .X(net6016));
 sky130_fd_sc_hd__buf_1 wire6017 (.A(net6014),
    .X(net6017));
 sky130_fd_sc_hd__clkbuf_1 fanout6018 (.A(net6035),
    .X(net6018));
 sky130_fd_sc_hd__buf_1 wire6019 (.A(net6020),
    .X(net6019));
 sky130_fd_sc_hd__buf_1 wire6020 (.A(net6023),
    .X(net6020));
 sky130_fd_sc_hd__clkbuf_2 wire6021 (.A(net6022),
    .X(net6021));
 sky130_fd_sc_hd__buf_1 wire6022 (.A(net6018),
    .X(net6022));
 sky130_fd_sc_hd__buf_1 max_length6023 (.A(net6018),
    .X(net6023));
 sky130_fd_sc_hd__buf_1 fanout6024 (.A(net6036),
    .X(net6024));
 sky130_fd_sc_hd__buf_1 wire6025 (.A(net6026),
    .X(net6025));
 sky130_fd_sc_hd__buf_1 wire6026 (.A(net6024),
    .X(net6026));
 sky130_fd_sc_hd__clkbuf_2 max_length6027 (.A(net6024),
    .X(net6027));
 sky130_fd_sc_hd__buf_1 fanout6028 (.A(net6036),
    .X(net6028));
 sky130_fd_sc_hd__buf_1 max_length6029 (.A(net6030),
    .X(net6029));
 sky130_fd_sc_hd__clkbuf_2 wire6030 (.A(net6028),
    .X(net6030));
 sky130_fd_sc_hd__buf_1 fanout6031 (.A(net6038),
    .X(net6031));
 sky130_fd_sc_hd__buf_1 wire6032 (.A(net6033),
    .X(net6032));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6033 (.A(net6031),
    .X(net6033));
 sky130_fd_sc_hd__buf_1 wire6034 (.A(net6031),
    .X(net6034));
 sky130_fd_sc_hd__buf_1 fanout6035 (.A(\cordic0.vec[0][16] ),
    .X(net6035));
 sky130_fd_sc_hd__buf_1 wire6036 (.A(net6037),
    .X(net6036));
 sky130_fd_sc_hd__buf_1 wire6037 (.A(net6038),
    .X(net6037));
 sky130_fd_sc_hd__buf_1 wire6038 (.A(net6039),
    .X(net6038));
 sky130_fd_sc_hd__clkbuf_1 wire6039 (.A(net6040),
    .X(net6039));
 sky130_fd_sc_hd__clkbuf_1 max_length6040 (.A(net6035),
    .X(net6040));
 sky130_fd_sc_hd__buf_1 fanout6041 (.A(net6047),
    .X(net6041));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6042 (.A(net6041),
    .X(net6042));
 sky130_fd_sc_hd__buf_1 wire6043 (.A(net6041),
    .X(net6043));
 sky130_fd_sc_hd__clkbuf_1 fanout6044 (.A(net6047),
    .X(net6044));
 sky130_fd_sc_hd__buf_1 max_length6045 (.A(net6046),
    .X(net6045));
 sky130_fd_sc_hd__buf_1 wire6046 (.A(net6044),
    .X(net6046));
 sky130_fd_sc_hd__buf_1 fanout6047 (.A(net6053),
    .X(net6047));
 sky130_fd_sc_hd__buf_1 wire6048 (.A(net6049),
    .X(net6048));
 sky130_fd_sc_hd__buf_2 wire6049 (.A(net6050),
    .X(net6049));
 sky130_fd_sc_hd__buf_1 wire6050 (.A(net6047),
    .X(net6050));
 sky130_fd_sc_hd__buf_1 fanout6051 (.A(\cordic0.vec[0][15] ),
    .X(net6051));
 sky130_fd_sc_hd__buf_1 wire6052 (.A(net6057),
    .X(net6052));
 sky130_fd_sc_hd__clkbuf_1 wire6053 (.A(net6054),
    .X(net6053));
 sky130_fd_sc_hd__clkbuf_1 max_length6054 (.A(net6057),
    .X(net6054));
 sky130_fd_sc_hd__buf_1 wire6055 (.A(net6056),
    .X(net6055));
 sky130_fd_sc_hd__clkbuf_1 max_length6056 (.A(net6051),
    .X(net6056));
 sky130_fd_sc_hd__clkbuf_2 max_length6057 (.A(net6051),
    .X(net6057));
 sky130_fd_sc_hd__buf_1 fanout6058 (.A(net6076),
    .X(net6058));
 sky130_fd_sc_hd__clkbuf_1 wire6059 (.A(net6060),
    .X(net6059));
 sky130_fd_sc_hd__buf_1 wire6060 (.A(net6062),
    .X(net6060));
 sky130_fd_sc_hd__buf_1 wire6061 (.A(net6062),
    .X(net6061));
 sky130_fd_sc_hd__buf_1 wire6062 (.A(net6058),
    .X(net6062));
 sky130_fd_sc_hd__clkbuf_2 fanout6063 (.A(net6076),
    .X(net6063));
 sky130_fd_sc_hd__clkbuf_1 fanout6064 (.A(net6068),
    .X(net6064));
 sky130_fd_sc_hd__buf_1 wire6065 (.A(net6066),
    .X(net6065));
 sky130_fd_sc_hd__buf_1 wire6066 (.A(net6067),
    .X(net6066));
 sky130_fd_sc_hd__clkbuf_2 wire6067 (.A(net6064),
    .X(net6067));
 sky130_fd_sc_hd__buf_1 fanout6068 (.A(net6075),
    .X(net6068));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6069 (.A(net6071),
    .X(net6069));
 sky130_fd_sc_hd__buf_1 max_length6070 (.A(net6071),
    .X(net6070));
 sky130_fd_sc_hd__buf_1 wire6071 (.A(net6072),
    .X(net6071));
 sky130_fd_sc_hd__buf_1 wire6072 (.A(net6068),
    .X(net6072));
 sky130_fd_sc_hd__buf_1 wire6073 (.A(net6074),
    .X(net6073));
 sky130_fd_sc_hd__clkbuf_1 wire6074 (.A(net6075),
    .X(net6074));
 sky130_fd_sc_hd__buf_1 wire6075 (.A(net6076),
    .X(net6075));
 sky130_fd_sc_hd__buf_1 wire6076 (.A(\cordic0.vec[0][14] ),
    .X(net6076));
 sky130_fd_sc_hd__clkbuf_2 fanout6077 (.A(net6083),
    .X(net6077));
 sky130_fd_sc_hd__buf_1 max_length6078 (.A(net6079),
    .X(net6078));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6079 (.A(net6077),
    .X(net6079));
 sky130_fd_sc_hd__buf_1 fanout6080 (.A(\cordic0.vec[0][13] ),
    .X(net6080));
 sky130_fd_sc_hd__clkbuf_2 wire6081 (.A(net6080),
    .X(net6081));
 sky130_fd_sc_hd__clkbuf_1 wire6082 (.A(net6080),
    .X(net6082));
 sky130_fd_sc_hd__clkbuf_1 max_length6083 (.A(net6080),
    .X(net6083));
 sky130_fd_sc_hd__buf_1 fanout6084 (.A(net6089),
    .X(net6084));
 sky130_fd_sc_hd__clkbuf_2 wire6085 (.A(net6084),
    .X(net6085));
 sky130_fd_sc_hd__buf_1 wire6086 (.A(net6087),
    .X(net6086));
 sky130_fd_sc_hd__buf_1 wire6087 (.A(net6084),
    .X(net6087));
 sky130_fd_sc_hd__clkbuf_2 fanout6088 (.A(net6090),
    .X(net6088));
 sky130_fd_sc_hd__clkbuf_1 max_length6089 (.A(net6090),
    .X(net6089));
 sky130_fd_sc_hd__buf_1 wire6090 (.A(\cordic0.vec[0][13] ),
    .X(net6090));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout6091 (.A(net6104),
    .X(net6091));
 sky130_fd_sc_hd__buf_1 wire6092 (.A(net6091),
    .X(net6092));
 sky130_fd_sc_hd__buf_1 wire6093 (.A(net6094),
    .X(net6093));
 sky130_fd_sc_hd__buf_1 wire6094 (.A(net6095),
    .X(net6094));
 sky130_fd_sc_hd__buf_1 wire6095 (.A(net6091),
    .X(net6095));
 sky130_fd_sc_hd__buf_1 fanout6096 (.A(net6100),
    .X(net6096));
 sky130_fd_sc_hd__clkbuf_2 wire6097 (.A(net6098),
    .X(net6097));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6098 (.A(net6099),
    .X(net6098));
 sky130_fd_sc_hd__buf_1 wire6099 (.A(net6096),
    .X(net6099));
 sky130_fd_sc_hd__buf_1 fanout6100 (.A(net6108),
    .X(net6100));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6101 (.A(net6102),
    .X(net6101));
 sky130_fd_sc_hd__buf_1 wire6102 (.A(net6103),
    .X(net6102));
 sky130_fd_sc_hd__buf_1 wire6103 (.A(net6100),
    .X(net6103));
 sky130_fd_sc_hd__clkbuf_1 fanout6104 (.A(\cordic0.vec[0][12] ),
    .X(net6104));
 sky130_fd_sc_hd__clkbuf_2 wire6105 (.A(net6106),
    .X(net6105));
 sky130_fd_sc_hd__clkbuf_1 wire6106 (.A(net6107),
    .X(net6106));
 sky130_fd_sc_hd__buf_1 wire6107 (.A(net6108),
    .X(net6107));
 sky130_fd_sc_hd__buf_1 wire6108 (.A(net6104),
    .X(net6108));
 sky130_fd_sc_hd__buf_1 fanout6109 (.A(net6123),
    .X(net6109));
 sky130_fd_sc_hd__buf_1 wire6110 (.A(net6111),
    .X(net6110));
 sky130_fd_sc_hd__buf_1 wire6111 (.A(net6109),
    .X(net6111));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6112 (.A(net6109),
    .X(net6112));
 sky130_fd_sc_hd__buf_1 fanout6113 (.A(net6118),
    .X(net6113));
 sky130_fd_sc_hd__buf_1 max_length6114 (.A(net6115),
    .X(net6114));
 sky130_fd_sc_hd__buf_1 wire6115 (.A(net6116),
    .X(net6115));
 sky130_fd_sc_hd__buf_1 wire6116 (.A(net6113),
    .X(net6116));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length6117 (.A(net6113),
    .X(net6117));
 sky130_fd_sc_hd__clkbuf_1 fanout6118 (.A(net6124),
    .X(net6118));
 sky130_fd_sc_hd__clkbuf_2 wire6119 (.A(net6121),
    .X(net6119));
 sky130_fd_sc_hd__clkbuf_1 wire6120 (.A(net6121),
    .X(net6120));
 sky130_fd_sc_hd__buf_1 wire6121 (.A(net6118),
    .X(net6121));
 sky130_fd_sc_hd__clkbuf_1 fanout6122 (.A(\cordic0.vec[0][11] ),
    .X(net6122));
 sky130_fd_sc_hd__buf_1 wire6123 (.A(net6122),
    .X(net6123));
 sky130_fd_sc_hd__clkbuf_1 wire6124 (.A(net6125),
    .X(net6124));
 sky130_fd_sc_hd__clkbuf_1 wire6125 (.A(net6126),
    .X(net6125));
 sky130_fd_sc_hd__clkbuf_1 wire6126 (.A(net6122),
    .X(net6126));
 sky130_fd_sc_hd__buf_1 fanout6127 (.A(net6135),
    .X(net6127));
 sky130_fd_sc_hd__buf_1 wire6128 (.A(net6130),
    .X(net6128));
 sky130_fd_sc_hd__buf_1 wire6129 (.A(net6130),
    .X(net6129));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6130 (.A(net6127),
    .X(net6130));
 sky130_fd_sc_hd__buf_1 max_length6131 (.A(net6127),
    .X(net6131));
 sky130_fd_sc_hd__buf_1 fanout6132 (.A(net6146),
    .X(net6132));
 sky130_fd_sc_hd__buf_1 wire6133 (.A(net6132),
    .X(net6133));
 sky130_fd_sc_hd__buf_1 wire6134 (.A(net6132),
    .X(net6134));
 sky130_fd_sc_hd__buf_1 max_length6135 (.A(net6136),
    .X(net6135));
 sky130_fd_sc_hd__buf_1 wire6136 (.A(net6137),
    .X(net6136));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6137 (.A(net6132),
    .X(net6137));
 sky130_fd_sc_hd__clkbuf_1 fanout6138 (.A(net6147),
    .X(net6138));
 sky130_fd_sc_hd__buf_1 wire6139 (.A(net6140),
    .X(net6139));
 sky130_fd_sc_hd__clkbuf_1 wire6140 (.A(net6145),
    .X(net6140));
 sky130_fd_sc_hd__clkbuf_1 wire6141 (.A(net6142),
    .X(net6141));
 sky130_fd_sc_hd__buf_1 wire6142 (.A(net6143),
    .X(net6142));
 sky130_fd_sc_hd__clkbuf_1 wire6143 (.A(net6144),
    .X(net6143));
 sky130_fd_sc_hd__clkbuf_1 wire6144 (.A(net6145),
    .X(net6144));
 sky130_fd_sc_hd__buf_1 wire6145 (.A(net6138),
    .X(net6145));
 sky130_fd_sc_hd__buf_1 fanout6146 (.A(\cordic0.vec[0][10] ),
    .X(net6146));
 sky130_fd_sc_hd__clkbuf_2 wire6147 (.A(net6148),
    .X(net6147));
 sky130_fd_sc_hd__buf_1 wire6148 (.A(net6149),
    .X(net6148));
 sky130_fd_sc_hd__clkbuf_1 wire6149 (.A(net6150),
    .X(net6149));
 sky130_fd_sc_hd__clkbuf_1 wire6150 (.A(net6146),
    .X(net6150));
 sky130_fd_sc_hd__clkbuf_2 fanout6151 (.A(net6160),
    .X(net6151));
 sky130_fd_sc_hd__clkbuf_2 wire6152 (.A(net6151),
    .X(net6152));
 sky130_fd_sc_hd__buf_1 fanout6153 (.A(net6158),
    .X(net6153));
 sky130_fd_sc_hd__buf_1 wire6154 (.A(net6153),
    .X(net6154));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6155 (.A(net6153),
    .X(net6155));
 sky130_fd_sc_hd__clkbuf_2 fanout6156 (.A(net6159),
    .X(net6156));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6157 (.A(net6156),
    .X(net6157));
 sky130_fd_sc_hd__buf_1 wire6158 (.A(net6156),
    .X(net6158));
 sky130_fd_sc_hd__buf_1 fanout6159 (.A(net6165),
    .X(net6159));
 sky130_fd_sc_hd__clkbuf_1 wire6160 (.A(net6161),
    .X(net6160));
 sky130_fd_sc_hd__clkbuf_1 wire6161 (.A(net6159),
    .X(net6161));
 sky130_fd_sc_hd__clkbuf_2 wire6162 (.A(net6163),
    .X(net6162));
 sky130_fd_sc_hd__buf_1 wire6163 (.A(net6159),
    .X(net6163));
 sky130_fd_sc_hd__buf_1 fanout6164 (.A(\cordic0.vec[0][9] ),
    .X(net6164));
 sky130_fd_sc_hd__clkbuf_1 wire6165 (.A(net6166),
    .X(net6165));
 sky130_fd_sc_hd__buf_1 wire6166 (.A(net6168),
    .X(net6166));
 sky130_fd_sc_hd__clkbuf_1 wire6167 (.A(net6164),
    .X(net6167));
 sky130_fd_sc_hd__clkbuf_2 max_length6168 (.A(net6164),
    .X(net6168));
 sky130_fd_sc_hd__clkbuf_2 fanout6169 (.A(net6193),
    .X(net6169));
 sky130_fd_sc_hd__buf_1 wire6170 (.A(net6171),
    .X(net6170));
 sky130_fd_sc_hd__clkbuf_1 wire6171 (.A(net6169),
    .X(net6171));
 sky130_fd_sc_hd__buf_1 wire6172 (.A(net6173),
    .X(net6172));
 sky130_fd_sc_hd__buf_1 wire6173 (.A(net6169),
    .X(net6173));
 sky130_fd_sc_hd__buf_1 wire6174 (.A(net6169),
    .X(net6174));
 sky130_fd_sc_hd__buf_1 fanout6175 (.A(net6192),
    .X(net6175));
 sky130_fd_sc_hd__buf_1 max_length6176 (.A(net6175),
    .X(net6176));
 sky130_fd_sc_hd__clkbuf_2 fanout6177 (.A(net6185),
    .X(net6177));
 sky130_fd_sc_hd__clkbuf_2 wire6178 (.A(net6177),
    .X(net6178));
 sky130_fd_sc_hd__buf_1 wire6179 (.A(net6177),
    .X(net6179));
 sky130_fd_sc_hd__clkbuf_1 max_length6180 (.A(net6177),
    .X(net6180));
 sky130_fd_sc_hd__clkbuf_2 max_length6181 (.A(net6177),
    .X(net6181));
 sky130_fd_sc_hd__buf_1 fanout6182 (.A(net6185),
    .X(net6182));
 sky130_fd_sc_hd__buf_1 max_length6183 (.A(net6184),
    .X(net6183));
 sky130_fd_sc_hd__buf_1 wire6184 (.A(net6182),
    .X(net6184));
 sky130_fd_sc_hd__buf_1 fanout6185 (.A(net6191),
    .X(net6185));
 sky130_fd_sc_hd__buf_1 wire6186 (.A(net6187),
    .X(net6186));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6187 (.A(net6188),
    .X(net6187));
 sky130_fd_sc_hd__clkbuf_1 max_length6188 (.A(net6189),
    .X(net6188));
 sky130_fd_sc_hd__buf_1 wire6189 (.A(net6190),
    .X(net6189));
 sky130_fd_sc_hd__clkbuf_1 wire6190 (.A(net6185),
    .X(net6190));
 sky130_fd_sc_hd__clkbuf_1 wire6191 (.A(net6193),
    .X(net6191));
 sky130_fd_sc_hd__clkbuf_1 max_length6192 (.A(net6193),
    .X(net6192));
 sky130_fd_sc_hd__buf_1 wire6193 (.A(\cordic0.vec[0][8] ),
    .X(net6193));
 sky130_fd_sc_hd__buf_1 fanout6194 (.A(net6214),
    .X(net6194));
 sky130_fd_sc_hd__buf_1 wire6195 (.A(net6196),
    .X(net6195));
 sky130_fd_sc_hd__buf_1 wire6196 (.A(net6197),
    .X(net6196));
 sky130_fd_sc_hd__clkbuf_1 max_length6197 (.A(net6198),
    .X(net6197));
 sky130_fd_sc_hd__buf_1 wire6198 (.A(net6199),
    .X(net6198));
 sky130_fd_sc_hd__buf_1 wire6199 (.A(net6194),
    .X(net6199));
 sky130_fd_sc_hd__buf_1 fanout6200 (.A(net6206),
    .X(net6200));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6201 (.A(net6200),
    .X(net6201));
 sky130_fd_sc_hd__buf_1 wire6202 (.A(net6203),
    .X(net6202));
 sky130_fd_sc_hd__buf_1 max_length6203 (.A(net6200),
    .X(net6203));
 sky130_fd_sc_hd__buf_1 fanout6204 (.A(net6206),
    .X(net6204));
 sky130_fd_sc_hd__buf_1 wire6205 (.A(net6204),
    .X(net6205));
 sky130_fd_sc_hd__buf_1 fanout6206 (.A(net6213),
    .X(net6206));
 sky130_fd_sc_hd__clkbuf_1 wire6207 (.A(net6208),
    .X(net6207));
 sky130_fd_sc_hd__buf_1 wire6208 (.A(net6209),
    .X(net6208));
 sky130_fd_sc_hd__buf_2 wire6209 (.A(net6210),
    .X(net6209));
 sky130_fd_sc_hd__clkbuf_1 wire6210 (.A(net6211),
    .X(net6210));
 sky130_fd_sc_hd__clkbuf_1 max_length6211 (.A(net6206),
    .X(net6211));
 sky130_fd_sc_hd__clkbuf_2 fanout6212 (.A(\cordic0.vec[0][7] ),
    .X(net6212));
 sky130_fd_sc_hd__clkbuf_1 wire6213 (.A(net6212),
    .X(net6213));
 sky130_fd_sc_hd__buf_1 wire6214 (.A(net6212),
    .X(net6214));
 sky130_fd_sc_hd__buf_1 fanout6215 (.A(net6239),
    .X(net6215));
 sky130_fd_sc_hd__buf_1 wire6216 (.A(net6217),
    .X(net6216));
 sky130_fd_sc_hd__buf_1 wire6217 (.A(net6215),
    .X(net6217));
 sky130_fd_sc_hd__buf_1 wire6218 (.A(net6219),
    .X(net6218));
 sky130_fd_sc_hd__buf_1 wire6219 (.A(net6215),
    .X(net6219));
 sky130_fd_sc_hd__clkbuf_2 fanout6220 (.A(net6223),
    .X(net6220));
 sky130_fd_sc_hd__clkbuf_1 max_length6221 (.A(net6222),
    .X(net6221));
 sky130_fd_sc_hd__buf_1 wire6222 (.A(net6220),
    .X(net6222));
 sky130_fd_sc_hd__clkbuf_1 fanout6223 (.A(net6228),
    .X(net6223));
 sky130_fd_sc_hd__buf_1 wire6224 (.A(net6227),
    .X(net6224));
 sky130_fd_sc_hd__buf_1 wire6225 (.A(net6226),
    .X(net6225));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6226 (.A(net6227),
    .X(net6226));
 sky130_fd_sc_hd__buf_1 wire6227 (.A(net6223),
    .X(net6227));
 sky130_fd_sc_hd__buf_1 fanout6228 (.A(net6237),
    .X(net6228));
 sky130_fd_sc_hd__clkbuf_2 wire6229 (.A(net6230),
    .X(net6229));
 sky130_fd_sc_hd__buf_1 wire6230 (.A(net6232),
    .X(net6230));
 sky130_fd_sc_hd__clkbuf_1 wire6231 (.A(net6232),
    .X(net6231));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6232 (.A(net6228),
    .X(net6232));
 sky130_fd_sc_hd__clkbuf_1 fanout6233 (.A(\cordic0.vec[0][6] ),
    .X(net6233));
 sky130_fd_sc_hd__clkbuf_1 wire6234 (.A(net6235),
    .X(net6234));
 sky130_fd_sc_hd__clkbuf_1 wire6235 (.A(net6236),
    .X(net6235));
 sky130_fd_sc_hd__clkbuf_1 wire6236 (.A(net6238),
    .X(net6236));
 sky130_fd_sc_hd__clkbuf_1 max_length6237 (.A(net6238),
    .X(net6237));
 sky130_fd_sc_hd__buf_1 wire6238 (.A(net6233),
    .X(net6238));
 sky130_fd_sc_hd__buf_1 wire6239 (.A(net6233),
    .X(net6239));
 sky130_fd_sc_hd__clkbuf_2 fanout6240 (.A(net6250),
    .X(net6240));
 sky130_fd_sc_hd__buf_1 wire6241 (.A(net6242),
    .X(net6241));
 sky130_fd_sc_hd__clkbuf_1 max_length6242 (.A(net6240),
    .X(net6242));
 sky130_fd_sc_hd__buf_1 fanout6243 (.A(net6251),
    .X(net6243));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6244 (.A(net6246),
    .X(net6244));
 sky130_fd_sc_hd__clkbuf_2 wire6245 (.A(net6246),
    .X(net6245));
 sky130_fd_sc_hd__buf_1 wire6246 (.A(net6243),
    .X(net6246));
 sky130_fd_sc_hd__buf_1 fanout6247 (.A(net6251),
    .X(net6247));
 sky130_fd_sc_hd__buf_1 wire6248 (.A(net6249),
    .X(net6248));
 sky130_fd_sc_hd__buf_1 wire6249 (.A(net6247),
    .X(net6249));
 sky130_fd_sc_hd__clkbuf_1 fanout6250 (.A(net6256),
    .X(net6250));
 sky130_fd_sc_hd__buf_1 wire6251 (.A(net6252),
    .X(net6251));
 sky130_fd_sc_hd__clkbuf_2 wire6252 (.A(net6250),
    .X(net6252));
 sky130_fd_sc_hd__buf_1 fanout6253 (.A(\cordic0.vec[0][5] ),
    .X(net6253));
 sky130_fd_sc_hd__buf_1 wire6254 (.A(net6255),
    .X(net6254));
 sky130_fd_sc_hd__buf_1 wire6255 (.A(net6253),
    .X(net6255));
 sky130_fd_sc_hd__clkbuf_1 max_length6256 (.A(net6257),
    .X(net6256));
 sky130_fd_sc_hd__buf_1 wire6257 (.A(net6253),
    .X(net6257));
 sky130_fd_sc_hd__clkbuf_2 fanout6258 (.A(net6283),
    .X(net6258));
 sky130_fd_sc_hd__buf_1 wire6259 (.A(net6258),
    .X(net6259));
 sky130_fd_sc_hd__buf_1 wire6260 (.A(net6258),
    .X(net6260));
 sky130_fd_sc_hd__clkbuf_2 fanout6261 (.A(net6282),
    .X(net6261));
 sky130_fd_sc_hd__buf_1 wire6262 (.A(net6261),
    .X(net6262));
 sky130_fd_sc_hd__clkbuf_1 max_length6263 (.A(net6261),
    .X(net6263));
 sky130_fd_sc_hd__clkbuf_1 fanout6264 (.A(net6273),
    .X(net6264));
 sky130_fd_sc_hd__buf_1 max_length6265 (.A(net6266),
    .X(net6265));
 sky130_fd_sc_hd__buf_1 wire6266 (.A(net6267),
    .X(net6266));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6267 (.A(net6264),
    .X(net6267));
 sky130_fd_sc_hd__clkbuf_2 fanout6268 (.A(net6282),
    .X(net6268));
 sky130_fd_sc_hd__buf_1 fanout6269 (.A(net6281),
    .X(net6269));
 sky130_fd_sc_hd__clkbuf_1 max_length6270 (.A(net6271),
    .X(net6270));
 sky130_fd_sc_hd__buf_2 wire6271 (.A(net6274),
    .X(net6271));
 sky130_fd_sc_hd__buf_1 wire6272 (.A(net6274),
    .X(net6272));
 sky130_fd_sc_hd__buf_1 wire6273 (.A(net6274),
    .X(net6273));
 sky130_fd_sc_hd__buf_1 wire6274 (.A(net6269),
    .X(net6274));
 sky130_fd_sc_hd__buf_1 fanout6275 (.A(net6285),
    .X(net6275));
 sky130_fd_sc_hd__buf_1 max_length6276 (.A(net6275),
    .X(net6276));
 sky130_fd_sc_hd__buf_1 wire6277 (.A(net6278),
    .X(net6277));
 sky130_fd_sc_hd__clkbuf_1 wire6278 (.A(net6279),
    .X(net6278));
 sky130_fd_sc_hd__clkbuf_1 wire6279 (.A(net6280),
    .X(net6279));
 sky130_fd_sc_hd__clkbuf_1 max_length6280 (.A(net6281),
    .X(net6280));
 sky130_fd_sc_hd__clkbuf_1 max_length6281 (.A(net6275),
    .X(net6281));
 sky130_fd_sc_hd__buf_1 wire6282 (.A(net6283),
    .X(net6282));
 sky130_fd_sc_hd__buf_1 wire6283 (.A(net6284),
    .X(net6283));
 sky130_fd_sc_hd__clkbuf_1 wire6284 (.A(net6285),
    .X(net6284));
 sky130_fd_sc_hd__buf_1 wire6285 (.A(\cordic0.vec[0][4] ),
    .X(net6285));
 sky130_fd_sc_hd__clkbuf_1 fanout6286 (.A(net6301),
    .X(net6286));
 sky130_fd_sc_hd__buf_1 max_length6287 (.A(net6289),
    .X(net6287));
 sky130_fd_sc_hd__buf_1 wire6288 (.A(net6289),
    .X(net6288));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6289 (.A(net6286),
    .X(net6289));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout6290 (.A(net6305),
    .X(net6290));
 sky130_fd_sc_hd__buf_1 fanout6291 (.A(net6304),
    .X(net6291));
 sky130_fd_sc_hd__clkbuf_2 max_length6292 (.A(net6293),
    .X(net6292));
 sky130_fd_sc_hd__buf_1 wire6293 (.A(net6291),
    .X(net6293));
 sky130_fd_sc_hd__buf_1 max_length6294 (.A(net6291),
    .X(net6294));
 sky130_fd_sc_hd__clkbuf_2 fanout6295 (.A(net6303),
    .X(net6295));
 sky130_fd_sc_hd__buf_1 wire6296 (.A(net6295),
    .X(net6296));
 sky130_fd_sc_hd__clkbuf_1 fanout6297 (.A(net6302),
    .X(net6297));
 sky130_fd_sc_hd__buf_1 wire6298 (.A(net6300),
    .X(net6298));
 sky130_fd_sc_hd__buf_1 wire6299 (.A(net6300),
    .X(net6299));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6300 (.A(net6297),
    .X(net6300));
 sky130_fd_sc_hd__buf_1 fanout6301 (.A(net6307),
    .X(net6301));
 sky130_fd_sc_hd__buf_1 wire6302 (.A(net6304),
    .X(net6302));
 sky130_fd_sc_hd__buf_1 wire6303 (.A(net6304),
    .X(net6303));
 sky130_fd_sc_hd__buf_1 wire6304 (.A(net6305),
    .X(net6304));
 sky130_fd_sc_hd__buf_1 max_length6305 (.A(net6301),
    .X(net6305));
 sky130_fd_sc_hd__buf_1 fanout6306 (.A(\cordic0.vec[0][3] ),
    .X(net6306));
 sky130_fd_sc_hd__clkbuf_1 wire6307 (.A(net6308),
    .X(net6307));
 sky130_fd_sc_hd__buf_1 wire6308 (.A(net6306),
    .X(net6308));
 sky130_fd_sc_hd__buf_1 wire6309 (.A(net6310),
    .X(net6309));
 sky130_fd_sc_hd__buf_1 wire6310 (.A(net6306),
    .X(net6310));
 sky130_fd_sc_hd__buf_1 fanout6311 (.A(net6314),
    .X(net6311));
 sky130_fd_sc_hd__buf_2 wire6312 (.A(net6311),
    .X(net6312));
 sky130_fd_sc_hd__clkbuf_2 fanout6313 (.A(net6316),
    .X(net6313));
 sky130_fd_sc_hd__buf_1 wire6314 (.A(net6313),
    .X(net6314));
 sky130_fd_sc_hd__buf_1 max_length6315 (.A(net6313),
    .X(net6315));
 sky130_fd_sc_hd__clkbuf_1 fanout6316 (.A(net6322),
    .X(net6316));
 sky130_fd_sc_hd__buf_1 wire6317 (.A(net6319),
    .X(net6317));
 sky130_fd_sc_hd__buf_1 max_length6318 (.A(net6319),
    .X(net6318));
 sky130_fd_sc_hd__clkbuf_2 wire6319 (.A(net6316),
    .X(net6319));
 sky130_fd_sc_hd__buf_1 fanout6320 (.A(net6330),
    .X(net6320));
 sky130_fd_sc_hd__buf_1 max_length6321 (.A(net6322),
    .X(net6321));
 sky130_fd_sc_hd__buf_1 max_length6322 (.A(net6323),
    .X(net6322));
 sky130_fd_sc_hd__buf_1 wire6323 (.A(net6320),
    .X(net6323));
 sky130_fd_sc_hd__clkbuf_2 fanout6324 (.A(\cordic0.vec[0][2] ),
    .X(net6324));
 sky130_fd_sc_hd__buf_1 wire6325 (.A(net6326),
    .X(net6325));
 sky130_fd_sc_hd__clkbuf_2 max_length6326 (.A(net6324),
    .X(net6326));
 sky130_fd_sc_hd__buf_1 wire6327 (.A(net6328),
    .X(net6327));
 sky130_fd_sc_hd__buf_1 wire6328 (.A(net6329),
    .X(net6328));
 sky130_fd_sc_hd__clkbuf_1 wire6329 (.A(net6330),
    .X(net6329));
 sky130_fd_sc_hd__buf_1 wire6330 (.A(net6331),
    .X(net6330));
 sky130_fd_sc_hd__clkbuf_1 wire6331 (.A(net6332),
    .X(net6331));
 sky130_fd_sc_hd__clkbuf_1 max_length6332 (.A(\cordic0.vec[0][2] ),
    .X(net6332));
 sky130_fd_sc_hd__clkbuf_1 fanout6333 (.A(net6346),
    .X(net6333));
 sky130_fd_sc_hd__buf_1 max_length6334 (.A(net6335),
    .X(net6334));
 sky130_fd_sc_hd__buf_1 wire6335 (.A(net6336),
    .X(net6335));
 sky130_fd_sc_hd__buf_1 wire6336 (.A(net6333),
    .X(net6336));
 sky130_fd_sc_hd__clkbuf_1 fanout6337 (.A(net6341),
    .X(net6337));
 sky130_fd_sc_hd__buf_1 wire6338 (.A(net6340),
    .X(net6338));
 sky130_fd_sc_hd__buf_1 wire6339 (.A(net6340),
    .X(net6339));
 sky130_fd_sc_hd__clkbuf_2 wire6340 (.A(net6337),
    .X(net6340));
 sky130_fd_sc_hd__buf_1 fanout6341 (.A(net6345),
    .X(net6341));
 sky130_fd_sc_hd__buf_1 wire6342 (.A(net6341),
    .X(net6342));
 sky130_fd_sc_hd__buf_1 wire6343 (.A(net6341),
    .X(net6343));
 sky130_fd_sc_hd__buf_1 fanout6344 (.A(\cordic0.vec[0][1] ),
    .X(net6344));
 sky130_fd_sc_hd__clkbuf_1 wire6345 (.A(net6346),
    .X(net6345));
 sky130_fd_sc_hd__clkbuf_2 wire6346 (.A(net6347),
    .X(net6346));
 sky130_fd_sc_hd__clkbuf_1 wire6347 (.A(net6348),
    .X(net6347));
 sky130_fd_sc_hd__clkbuf_1 wire6348 (.A(net6349),
    .X(net6348));
 sky130_fd_sc_hd__clkbuf_1 wire6349 (.A(net6350),
    .X(net6349));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length6350 (.A(net6344),
    .X(net6350));
 sky130_fd_sc_hd__clkbuf_1 fanout6351 (.A(net6354),
    .X(net6351));
 sky130_fd_sc_hd__buf_2 wire6352 (.A(net6351),
    .X(net6352));
 sky130_fd_sc_hd__buf_1 fanout6353 (.A(net6361),
    .X(net6353));
 sky130_fd_sc_hd__buf_1 wire6354 (.A(net6353),
    .X(net6354));
 sky130_fd_sc_hd__buf_1 wire6355 (.A(net6357),
    .X(net6355));
 sky130_fd_sc_hd__buf_1 max_length6356 (.A(net6357),
    .X(net6356));
 sky130_fd_sc_hd__buf_1 wire6357 (.A(net6353),
    .X(net6357));
 sky130_fd_sc_hd__buf_1 fanout6358 (.A(net6365),
    .X(net6358));
 sky130_fd_sc_hd__buf_1 wire6359 (.A(net6361),
    .X(net6359));
 sky130_fd_sc_hd__clkbuf_1 wire6360 (.A(net6361),
    .X(net6360));
 sky130_fd_sc_hd__buf_1 wire6361 (.A(net6362),
    .X(net6361));
 sky130_fd_sc_hd__buf_1 wire6362 (.A(net6358),
    .X(net6362));
 sky130_fd_sc_hd__buf_1 wire6363 (.A(net6364),
    .X(net6363));
 sky130_fd_sc_hd__clkbuf_1 wire6364 (.A(\cordic0.vec[0][0] ),
    .X(net6364));
 sky130_fd_sc_hd__clkbuf_1 wire6365 (.A(net6366),
    .X(net6365));
 sky130_fd_sc_hd__clkbuf_1 wire6366 (.A(net6367),
    .X(net6366));
 sky130_fd_sc_hd__clkbuf_1 max_length6367 (.A(\cordic0.vec[0][0] ),
    .X(net6367));
 sky130_fd_sc_hd__buf_1 wire6368 (.A(\cordic0.slte0.opA[15] ),
    .X(net6368));
 sky130_fd_sc_hd__clkbuf_2 wire6369 (.A(\cordic0.slte0.opA[13] ),
    .X(net6369));
 sky130_fd_sc_hd__buf_1 wire6370 (.A(\cordic0.slte0.opA[12] ),
    .X(net6370));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6371 (.A(\cordic0.slte0.opA[11] ),
    .X(net6371));
 sky130_fd_sc_hd__buf_1 wire6372 (.A(\cordic0.slte0.opA[10] ),
    .X(net6372));
 sky130_fd_sc_hd__buf_1 wire6373 (.A(\cordic0.slte0.opA[7] ),
    .X(net6373));
 sky130_fd_sc_hd__clkbuf_2 wire6374 (.A(\cordic0.slte0.opA[6] ),
    .X(net6374));
 sky130_fd_sc_hd__buf_1 fanout6375 (.A(net6378),
    .X(net6375));
 sky130_fd_sc_hd__clkbuf_2 wire6376 (.A(net6375),
    .X(net6376));
 sky130_fd_sc_hd__buf_1 fanout6377 (.A(net6380),
    .X(net6377));
 sky130_fd_sc_hd__buf_1 wire6378 (.A(net6377),
    .X(net6378));
 sky130_fd_sc_hd__buf_1 wire6379 (.A(net6377),
    .X(net6379));
 sky130_fd_sc_hd__clkbuf_1 wire6380 (.A(net6381),
    .X(net6380));
 sky130_fd_sc_hd__clkbuf_1 wire6381 (.A(net6382),
    .X(net6381));
 sky130_fd_sc_hd__buf_1 wire6382 (.A(net6383),
    .X(net6382));
 sky130_fd_sc_hd__clkbuf_1 wire6383 (.A(net6384),
    .X(net6383));
 sky130_fd_sc_hd__clkbuf_1 wire6384 (.A(net6385),
    .X(net6384));
 sky130_fd_sc_hd__clkbuf_1 wire6385 (.A(\cordic0.domain[1] ),
    .X(net6385));
 sky130_fd_sc_hd__buf_1 wire6386 (.A(net6387),
    .X(net6386));
 sky130_fd_sc_hd__clkbuf_1 wire6387 (.A(net6388),
    .X(net6387));
 sky130_fd_sc_hd__clkbuf_1 wire6388 (.A(net6389),
    .X(net6388));
 sky130_fd_sc_hd__clkbuf_1 wire6389 (.A(\cordic0.domain[0] ),
    .X(net6389));
 sky130_fd_sc_hd__clkbuf_1 wire6390 (.A(net6391),
    .X(net6390));
 sky130_fd_sc_hd__clkbuf_1 wire6391 (.A(net6392),
    .X(net6391));
 sky130_fd_sc_hd__clkbuf_1 wire6392 (.A(\cordic0.slte0.opB[15] ),
    .X(net6392));
 sky130_fd_sc_hd__buf_1 wire6393 (.A(net6394),
    .X(net6393));
 sky130_fd_sc_hd__clkbuf_1 wire6394 (.A(net6395),
    .X(net6394));
 sky130_fd_sc_hd__clkbuf_1 wire6395 (.A(\cordic0.slte0.opB[14] ),
    .X(net6395));
 sky130_fd_sc_hd__buf_1 wire6396 (.A(net6397),
    .X(net6396));
 sky130_fd_sc_hd__clkbuf_1 wire6397 (.A(net6398),
    .X(net6397));
 sky130_fd_sc_hd__clkbuf_1 wire6398 (.A(\cordic0.slte0.opB[13] ),
    .X(net6398));
 sky130_fd_sc_hd__buf_1 wire6399 (.A(net6400),
    .X(net6399));
 sky130_fd_sc_hd__clkbuf_1 wire6400 (.A(net6401),
    .X(net6400));
 sky130_fd_sc_hd__clkbuf_1 wire6401 (.A(\cordic0.slte0.opB[12] ),
    .X(net6401));
 sky130_fd_sc_hd__buf_1 wire6402 (.A(net6403),
    .X(net6402));
 sky130_fd_sc_hd__clkbuf_1 wire6403 (.A(\cordic0.slte0.opB[10] ),
    .X(net6403));
 sky130_fd_sc_hd__buf_1 wire6404 (.A(net6405),
    .X(net6404));
 sky130_fd_sc_hd__clkbuf_1 wire6405 (.A(net6406),
    .X(net6405));
 sky130_fd_sc_hd__clkbuf_1 wire6406 (.A(\cordic0.slte0.opB[9] ),
    .X(net6406));
 sky130_fd_sc_hd__buf_1 wire6407 (.A(net6408),
    .X(net6407));
 sky130_fd_sc_hd__clkbuf_1 wire6408 (.A(net6409),
    .X(net6408));
 sky130_fd_sc_hd__clkbuf_1 wire6409 (.A(\cordic0.slte0.opB[8] ),
    .X(net6409));
 sky130_fd_sc_hd__buf_1 wire6410 (.A(net6411),
    .X(net6410));
 sky130_fd_sc_hd__clkbuf_1 wire6411 (.A(net6412),
    .X(net6411));
 sky130_fd_sc_hd__buf_1 wire6412 (.A(\cordic0.slte0.opB[7] ),
    .X(net6412));
 sky130_fd_sc_hd__clkbuf_1 wire6413 (.A(net6414),
    .X(net6413));
 sky130_fd_sc_hd__clkbuf_1 wire6414 (.A(net6415),
    .X(net6414));
 sky130_fd_sc_hd__buf_1 wire6415 (.A(\cordic0.slte0.opB[6] ),
    .X(net6415));
 sky130_fd_sc_hd__buf_1 wire6416 (.A(net6417),
    .X(net6416));
 sky130_fd_sc_hd__clkbuf_1 max_length6417 (.A(\cordic0.slte0.opB[5] ),
    .X(net6417));
 sky130_fd_sc_hd__buf_1 wire6418 (.A(\cordic0.slte0.opB[4] ),
    .X(net6418));
 sky130_fd_sc_hd__clkbuf_1 wire6419 (.A(\cordic0.slte0.opB[3] ),
    .X(net6419));
 sky130_fd_sc_hd__clkbuf_1 wire6420 (.A(\cordic0.slte0.opB[2] ),
    .X(net6420));
 sky130_fd_sc_hd__clkbuf_1 wire6421 (.A(\cordic0.sin[11] ),
    .X(net6421));
 sky130_fd_sc_hd__clkbuf_1 wire6422 (.A(\cordic0.sin[10] ),
    .X(net6422));
 sky130_fd_sc_hd__clkbuf_1 wire6423 (.A(\cordic0.sin[8] ),
    .X(net6423));
 sky130_fd_sc_hd__clkbuf_1 wire6424 (.A(\cordic0.sin[7] ),
    .X(net6424));
 sky130_fd_sc_hd__clkbuf_1 wire6425 (.A(net6426),
    .X(net6425));
 sky130_fd_sc_hd__clkbuf_1 max_length6426 (.A(\cordic0.sin[5] ),
    .X(net6426));
 sky130_fd_sc_hd__clkbuf_1 wire6427 (.A(\cordic0.sin[4] ),
    .X(net6427));
 sky130_fd_sc_hd__clkbuf_1 wire6428 (.A(net6429),
    .X(net6428));
 sky130_fd_sc_hd__clkbuf_1 wire6429 (.A(\cordic0.sin[3] ),
    .X(net6429));
 sky130_fd_sc_hd__clkbuf_1 wire6430 (.A(\cordic0.sin[1] ),
    .X(net6430));
 sky130_fd_sc_hd__clkbuf_1 wire6431 (.A(\cordic0.sin[0] ),
    .X(net6431));
 sky130_fd_sc_hd__buf_1 wire6432 (.A(net6433),
    .X(net6432));
 sky130_fd_sc_hd__clkbuf_1 wire6433 (.A(net6434),
    .X(net6433));
 sky130_fd_sc_hd__clkbuf_1 wire6434 (.A(net6435),
    .X(net6434));
 sky130_fd_sc_hd__clkbuf_1 wire6435 (.A(net6436),
    .X(net6435));
 sky130_fd_sc_hd__clkbuf_1 wire6436 (.A(net6437),
    .X(net6436));
 sky130_fd_sc_hd__clkbuf_1 wire6437 (.A(net6438),
    .X(net6437));
 sky130_fd_sc_hd__clkbuf_1 wire6438 (.A(net6439),
    .X(net6438));
 sky130_fd_sc_hd__clkbuf_1 wire6439 (.A(net6440),
    .X(net6439));
 sky130_fd_sc_hd__clkbuf_1 wire6440 (.A(net6441),
    .X(net6440));
 sky130_fd_sc_hd__clkbuf_1 wire6441 (.A(net6442),
    .X(net6441));
 sky130_fd_sc_hd__clkbuf_1 wire6442 (.A(\cordic0.out_valid ),
    .X(net6442));
 sky130_fd_sc_hd__buf_2 fanout6443 (.A(net6444),
    .X(net6443));
 sky130_fd_sc_hd__buf_1 fanout6444 (.A(\state[2] ),
    .X(net6444));
 sky130_fd_sc_hd__buf_1 wire6445 (.A(net6446),
    .X(net6445));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6446 (.A(net6444),
    .X(net6446));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout6447 (.A(\state[1] ),
    .X(net6447));
 sky130_fd_sc_hd__buf_1 max_length6448 (.A(net6449),
    .X(net6448));
 sky130_fd_sc_hd__buf_1 wire6449 (.A(net6447),
    .X(net6449));
 sky130_fd_sc_hd__clkbuf_1 fanout6450 (.A(\state[1] ),
    .X(net6450));
 sky130_fd_sc_hd__clkbuf_2 wire6451 (.A(net6450),
    .X(net6451));
 sky130_fd_sc_hd__clkbuf_1 fanout6452 (.A(\state[0] ),
    .X(net6452));
 sky130_fd_sc_hd__clkbuf_2 max_length6453 (.A(net6454),
    .X(net6453));
 sky130_fd_sc_hd__clkbuf_2 wire6454 (.A(net6452),
    .X(net6454));
 sky130_fd_sc_hd__buf_1 fanout6455 (.A(\state[0] ),
    .X(net6455));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6456 (.A(net6455),
    .X(net6456));
 sky130_fd_sc_hd__buf_1 fanout6457 (.A(net6463),
    .X(net6457));
 sky130_fd_sc_hd__buf_1 wire6458 (.A(net6459),
    .X(net6458));
 sky130_fd_sc_hd__clkbuf_2 max_length6459 (.A(net6457),
    .X(net6459));
 sky130_fd_sc_hd__clkbuf_2 fanout6460 (.A(net6465),
    .X(net6460));
 sky130_fd_sc_hd__buf_1 wire6461 (.A(net6460),
    .X(net6461));
 sky130_fd_sc_hd__buf_1 max_length6462 (.A(net6460),
    .X(net6462));
 sky130_fd_sc_hd__buf_1 fanout6463 (.A(\cordic0.gm0.iter[4] ),
    .X(net6463));
 sky130_fd_sc_hd__clkbuf_1 wire6464 (.A(net6465),
    .X(net6464));
 sky130_fd_sc_hd__buf_1 wire6465 (.A(net6463),
    .X(net6465));
 sky130_fd_sc_hd__buf_1 wire6466 (.A(net6463),
    .X(net6466));
 sky130_fd_sc_hd__clkbuf_2 fanout6467 (.A(net6469),
    .X(net6467));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6468 (.A(net6467),
    .X(net6468));
 sky130_fd_sc_hd__buf_1 fanout6469 (.A(\cordic0.gm0.iter[3] ),
    .X(net6469));
 sky130_fd_sc_hd__buf_1 wire6470 (.A(net6473),
    .X(net6470));
 sky130_fd_sc_hd__buf_1 wire6471 (.A(net6472),
    .X(net6471));
 sky130_fd_sc_hd__buf_1 wire6472 (.A(net6473),
    .X(net6472));
 sky130_fd_sc_hd__buf_1 wire6473 (.A(net6469),
    .X(net6473));
 sky130_fd_sc_hd__clkbuf_1 wire6474 (.A(\cordic0.gm0.iter[3] ),
    .X(net6474));
 sky130_fd_sc_hd__buf_1 fanout6475 (.A(net6481),
    .X(net6475));
 sky130_fd_sc_hd__clkbuf_1 max_length6476 (.A(net6477),
    .X(net6476));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6477 (.A(net6478),
    .X(net6477));
 sky130_fd_sc_hd__buf_1 max_length6478 (.A(net6475),
    .X(net6478));
 sky130_fd_sc_hd__buf_1 fanout6479 (.A(net6482),
    .X(net6479));
 sky130_fd_sc_hd__buf_1 wire6480 (.A(net6479),
    .X(net6480));
 sky130_fd_sc_hd__buf_1 fanout6481 (.A(\cordic0.gm0.iter[2] ),
    .X(net6481));
 sky130_fd_sc_hd__clkbuf_1 wire6482 (.A(net6481),
    .X(net6482));
 sky130_fd_sc_hd__buf_1 wire6483 (.A(net6484),
    .X(net6483));
 sky130_fd_sc_hd__buf_1 wire6484 (.A(net6485),
    .X(net6484));
 sky130_fd_sc_hd__buf_1 wire6485 (.A(net6481),
    .X(net6485));
 sky130_fd_sc_hd__clkbuf_1 wire6486 (.A(net6487),
    .X(net6486));
 sky130_fd_sc_hd__clkbuf_1 wire6487 (.A(\cordic0.gm0.iter[2] ),
    .X(net6487));
 sky130_fd_sc_hd__clkbuf_1 fanout6488 (.A(net6492),
    .X(net6488));
 sky130_fd_sc_hd__clkbuf_2 wire6489 (.A(net6490),
    .X(net6489));
 sky130_fd_sc_hd__clkbuf_2 wire6490 (.A(net6488),
    .X(net6490));
 sky130_fd_sc_hd__clkbuf_2 fanout6491 (.A(net6497),
    .X(net6491));
 sky130_fd_sc_hd__clkbuf_1 fanout6492 (.A(net6505),
    .X(net6492));
 sky130_fd_sc_hd__buf_1 wire6493 (.A(net6495),
    .X(net6493));
 sky130_fd_sc_hd__buf_1 max_length6494 (.A(net6495),
    .X(net6494));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length6495 (.A(net6496),
    .X(net6495));
 sky130_fd_sc_hd__clkbuf_1 wire6496 (.A(net6497),
    .X(net6496));
 sky130_fd_sc_hd__buf_1 wire6497 (.A(net6492),
    .X(net6497));
 sky130_fd_sc_hd__buf_2 fanout6498 (.A(net6504),
    .X(net6498));
 sky130_fd_sc_hd__buf_1 wire6499 (.A(net6500),
    .X(net6499));
 sky130_fd_sc_hd__buf_1 wire6500 (.A(net6498),
    .X(net6500));
 sky130_fd_sc_hd__buf_2 fanout6501 (.A(net6503),
    .X(net6501));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6502 (.A(net6501),
    .X(net6502));
 sky130_fd_sc_hd__clkbuf_1 fanout6503 (.A(\cordic0.gm0.iter[1] ),
    .X(net6503));
 sky130_fd_sc_hd__clkbuf_2 wire6504 (.A(net6503),
    .X(net6504));
 sky130_fd_sc_hd__clkbuf_1 wire6505 (.A(\cordic0.gm0.iter[1] ),
    .X(net6505));
 sky130_fd_sc_hd__buf_1 fanout6506 (.A(\cordic0.gm0.iter[0] ),
    .X(net6506));
 sky130_fd_sc_hd__clkbuf_1 wire6507 (.A(net6510),
    .X(net6507));
 sky130_fd_sc_hd__buf_1 wire6508 (.A(net6509),
    .X(net6508));
 sky130_fd_sc_hd__buf_1 wire6509 (.A(net6510),
    .X(net6509));
 sky130_fd_sc_hd__buf_1 wire6510 (.A(net6511),
    .X(net6510));
 sky130_fd_sc_hd__buf_1 wire6511 (.A(net6506),
    .X(net6511));
 sky130_fd_sc_hd__buf_1 fanout6512 (.A(net6528),
    .X(net6512));
 sky130_fd_sc_hd__buf_1 max_length6513 (.A(net6514),
    .X(net6513));
 sky130_fd_sc_hd__clkbuf_2 max_length6514 (.A(net6512),
    .X(net6514));
 sky130_fd_sc_hd__clkbuf_2 fanout6515 (.A(net6517),
    .X(net6515));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6516 (.A(net6515),
    .X(net6516));
 sky130_fd_sc_hd__clkbuf_1 fanout6517 (.A(net6524),
    .X(net6517));
 sky130_fd_sc_hd__clkbuf_2 max_length6518 (.A(net6519),
    .X(net6518));
 sky130_fd_sc_hd__buf_1 wire6519 (.A(net6520),
    .X(net6519));
 sky130_fd_sc_hd__buf_1 wire6520 (.A(net6517),
    .X(net6520));
 sky130_fd_sc_hd__clkbuf_2 fanout6521 (.A(net6526),
    .X(net6521));
 sky130_fd_sc_hd__buf_1 max_length6522 (.A(net6523),
    .X(net6522));
 sky130_fd_sc_hd__buf_1 max_length6523 (.A(net6521),
    .X(net6523));
 sky130_fd_sc_hd__clkbuf_1 fanout6524 (.A(net6529),
    .X(net6524));
 sky130_fd_sc_hd__clkbuf_2 wire6525 (.A(net6526),
    .X(net6525));
 sky130_fd_sc_hd__buf_1 wire6526 (.A(net6527),
    .X(net6526));
 sky130_fd_sc_hd__clkbuf_1 max_length6527 (.A(net6524),
    .X(net6527));
 sky130_fd_sc_hd__clkbuf_1 wire6528 (.A(net6530),
    .X(net6528));
 sky130_fd_sc_hd__clkbuf_1 wire6529 (.A(net6530),
    .X(net6529));
 sky130_fd_sc_hd__buf_1 wire6530 (.A(\cordic0.gm0.iter[0] ),
    .X(net6530));
 sky130_fd_sc_hd__buf_1 fanout6531 (.A(net6538),
    .X(net6531));
 sky130_fd_sc_hd__buf_1 wire6532 (.A(net6533),
    .X(net6532));
 sky130_fd_sc_hd__clkbuf_2 wire6533 (.A(net6531),
    .X(net6533));
 sky130_fd_sc_hd__buf_1 wire6534 (.A(net6531),
    .X(net6534));
 sky130_fd_sc_hd__buf_1 fanout6535 (.A(net6545),
    .X(net6535));
 sky130_fd_sc_hd__clkbuf_1 max_length6536 (.A(net6537),
    .X(net6536));
 sky130_fd_sc_hd__buf_1 wire6537 (.A(net6535),
    .X(net6537));
 sky130_fd_sc_hd__buf_1 wire6538 (.A(net6535),
    .X(net6538));
 sky130_fd_sc_hd__buf_1 fanout6539 (.A(net6544),
    .X(net6539));
 sky130_fd_sc_hd__buf_1 max_length6540 (.A(net6541),
    .X(net6540));
 sky130_fd_sc_hd__buf_1 wire6541 (.A(net6539),
    .X(net6541));
 sky130_fd_sc_hd__buf_1 wire6542 (.A(net6539),
    .X(net6542));
 sky130_fd_sc_hd__buf_1 max_length6543 (.A(net6539),
    .X(net6543));
 sky130_fd_sc_hd__buf_1 fanout6544 (.A(net6566),
    .X(net6544));
 sky130_fd_sc_hd__buf_1 wire6545 (.A(net6544),
    .X(net6545));
 sky130_fd_sc_hd__buf_1 wire6546 (.A(net6544),
    .X(net6546));
 sky130_fd_sc_hd__buf_1 fanout6547 (.A(net6562),
    .X(net6547));
 sky130_fd_sc_hd__buf_1 wire6548 (.A(net6549),
    .X(net6548));
 sky130_fd_sc_hd__buf_1 wire6549 (.A(net6551),
    .X(net6549));
 sky130_fd_sc_hd__buf_1 wire6550 (.A(net6551),
    .X(net6550));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6551 (.A(net6552),
    .X(net6551));
 sky130_fd_sc_hd__buf_1 wire6552 (.A(net6547),
    .X(net6552));
 sky130_fd_sc_hd__clkbuf_1 fanout6553 (.A(net6564),
    .X(net6553));
 sky130_fd_sc_hd__clkbuf_1 wire6554 (.A(net6562),
    .X(net6554));
 sky130_fd_sc_hd__clkbuf_1 wire6555 (.A(net6556),
    .X(net6555));
 sky130_fd_sc_hd__buf_1 wire6556 (.A(net6559),
    .X(net6556));
 sky130_fd_sc_hd__buf_1 wire6557 (.A(net6558),
    .X(net6557));
 sky130_fd_sc_hd__buf_1 wire6558 (.A(net6559),
    .X(net6558));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6559 (.A(net6560),
    .X(net6559));
 sky130_fd_sc_hd__clkbuf_1 wire6560 (.A(net6561),
    .X(net6560));
 sky130_fd_sc_hd__clkbuf_1 wire6561 (.A(net6562),
    .X(net6561));
 sky130_fd_sc_hd__buf_1 wire6562 (.A(net6553),
    .X(net6562));
 sky130_fd_sc_hd__buf_1 wire6563 (.A(net6564),
    .X(net6563));
 sky130_fd_sc_hd__buf_1 wire6564 (.A(net6565),
    .X(net6564));
 sky130_fd_sc_hd__clkbuf_1 wire6565 (.A(net6566),
    .X(net6565));
 sky130_fd_sc_hd__buf_1 wire6566 (.A(\matmul0.matmul_stage_inst.state[6] ),
    .X(net6566));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout6567 (.A(net6576),
    .X(net6567));
 sky130_fd_sc_hd__buf_1 wire6568 (.A(net6569),
    .X(net6568));
 sky130_fd_sc_hd__buf_1 wire6569 (.A(net6567),
    .X(net6569));
 sky130_fd_sc_hd__buf_1 max_length6570 (.A(net6571),
    .X(net6570));
 sky130_fd_sc_hd__buf_1 max_length6571 (.A(net6567),
    .X(net6571));
 sky130_fd_sc_hd__buf_1 fanout6572 (.A(net6579),
    .X(net6572));
 sky130_fd_sc_hd__clkbuf_1 wire6573 (.A(net6574),
    .X(net6573));
 sky130_fd_sc_hd__buf_1 max_length6574 (.A(net6575),
    .X(net6574));
 sky130_fd_sc_hd__buf_1 wire6575 (.A(net6578),
    .X(net6575));
 sky130_fd_sc_hd__clkbuf_1 wire6576 (.A(net6577),
    .X(net6576));
 sky130_fd_sc_hd__clkbuf_1 wire6577 (.A(net6578),
    .X(net6577));
 sky130_fd_sc_hd__buf_1 wire6578 (.A(net6572),
    .X(net6578));
 sky130_fd_sc_hd__clkbuf_1 wire6579 (.A(\matmul0.matmul_stage_inst.state[5] ),
    .X(net6579));
 sky130_fd_sc_hd__buf_1 fanout6580 (.A(net6585),
    .X(net6580));
 sky130_fd_sc_hd__buf_1 wire6581 (.A(net6580),
    .X(net6581));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6582 (.A(net6583),
    .X(net6582));
 sky130_fd_sc_hd__buf_1 wire6583 (.A(net6580),
    .X(net6583));
 sky130_fd_sc_hd__clkbuf_1 fanout6584 (.A(net6586),
    .X(net6584));
 sky130_fd_sc_hd__clkbuf_2 wire6585 (.A(net6584),
    .X(net6585));
 sky130_fd_sc_hd__buf_1 fanout6586 (.A(net6591),
    .X(net6586));
 sky130_fd_sc_hd__buf_1 wire6587 (.A(net6588),
    .X(net6587));
 sky130_fd_sc_hd__buf_1 wire6588 (.A(net6590),
    .X(net6588));
 sky130_fd_sc_hd__clkbuf_1 wire6589 (.A(net6586),
    .X(net6589));
 sky130_fd_sc_hd__clkbuf_1 max_length6590 (.A(net6586),
    .X(net6590));
 sky130_fd_sc_hd__buf_1 fanout6591 (.A(\matmul0.matmul_stage_inst.state[4] ),
    .X(net6591));
 sky130_fd_sc_hd__buf_1 max_length6592 (.A(net6594),
    .X(net6592));
 sky130_fd_sc_hd__clkbuf_1 wire6593 (.A(net6595),
    .X(net6593));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length6594 (.A(net6595),
    .X(net6594));
 sky130_fd_sc_hd__buf_1 wire6595 (.A(net6596),
    .X(net6595));
 sky130_fd_sc_hd__clkbuf_1 wire6596 (.A(net6591),
    .X(net6596));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout6597 (.A(net6608),
    .X(net6597));
 sky130_fd_sc_hd__clkbuf_1 wire6598 (.A(net6599),
    .X(net6598));
 sky130_fd_sc_hd__buf_1 wire6599 (.A(net6600),
    .X(net6599));
 sky130_fd_sc_hd__buf_1 wire6600 (.A(net6601),
    .X(net6600));
 sky130_fd_sc_hd__clkbuf_1 wire6601 (.A(net6602),
    .X(net6601));
 sky130_fd_sc_hd__clkbuf_1 wire6602 (.A(net6603),
    .X(net6602));
 sky130_fd_sc_hd__buf_1 wire6603 (.A(net6597),
    .X(net6603));
 sky130_fd_sc_hd__clkbuf_1 wire6604 (.A(net6605),
    .X(net6604));
 sky130_fd_sc_hd__clkbuf_1 wire6605 (.A(net6606),
    .X(net6605));
 sky130_fd_sc_hd__clkbuf_1 wire6606 (.A(net6607),
    .X(net6606));
 sky130_fd_sc_hd__clkbuf_1 wire6607 (.A(net6608),
    .X(net6607));
 sky130_fd_sc_hd__buf_1 wire6608 (.A(\matmul0.done_pass ),
    .X(net6608));
 sky130_fd_sc_hd__clkbuf_1 fanout6609 (.A(net6623),
    .X(net6609));
 sky130_fd_sc_hd__buf_1 wire6610 (.A(net6612),
    .X(net6610));
 sky130_fd_sc_hd__buf_1 max_length6611 (.A(net6612),
    .X(net6611));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6612 (.A(net6609),
    .X(net6612));
 sky130_fd_sc_hd__buf_1 fanout6613 (.A(net6625),
    .X(net6613));
 sky130_fd_sc_hd__buf_1 wire6614 (.A(net6615),
    .X(net6614));
 sky130_fd_sc_hd__buf_1 wire6615 (.A(net6613),
    .X(net6615));
 sky130_fd_sc_hd__buf_1 wire6616 (.A(net6617),
    .X(net6616));
 sky130_fd_sc_hd__buf_1 wire6617 (.A(net6613),
    .X(net6617));
 sky130_fd_sc_hd__clkbuf_1 fanout6618 (.A(net6622),
    .X(net6618));
 sky130_fd_sc_hd__buf_1 wire6619 (.A(net6620),
    .X(net6619));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6620 (.A(net6621),
    .X(net6620));
 sky130_fd_sc_hd__buf_1 wire6621 (.A(net6618),
    .X(net6621));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout6622 (.A(\matmul0.matmul_stage_inst.state[2] ),
    .X(net6622));
 sky130_fd_sc_hd__clkbuf_1 wire6623 (.A(net6624),
    .X(net6623));
 sky130_fd_sc_hd__clkbuf_1 max_length6624 (.A(net6625),
    .X(net6624));
 sky130_fd_sc_hd__buf_1 wire6625 (.A(\matmul0.matmul_stage_inst.state[2] ),
    .X(net6625));
 sky130_fd_sc_hd__clkbuf_1 fanout6626 (.A(net6633),
    .X(net6626));
 sky130_fd_sc_hd__clkbuf_1 wire6627 (.A(net6628),
    .X(net6627));
 sky130_fd_sc_hd__clkbuf_1 wire6628 (.A(net6626),
    .X(net6628));
 sky130_fd_sc_hd__buf_1 max_length6629 (.A(net6630),
    .X(net6629));
 sky130_fd_sc_hd__buf_1 wire6630 (.A(net6631),
    .X(net6630));
 sky130_fd_sc_hd__clkbuf_2 wire6631 (.A(net6626),
    .X(net6631));
 sky130_fd_sc_hd__clkbuf_1 fanout6632 (.A(net6648),
    .X(net6632));
 sky130_fd_sc_hd__clkbuf_1 wire6633 (.A(net6636),
    .X(net6633));
 sky130_fd_sc_hd__buf_1 wire6634 (.A(net6636),
    .X(net6634));
 sky130_fd_sc_hd__clkbuf_1 max_length6635 (.A(net6636),
    .X(net6635));
 sky130_fd_sc_hd__buf_1 wire6636 (.A(net6637),
    .X(net6636));
 sky130_fd_sc_hd__clkbuf_1 wire6637 (.A(net6632),
    .X(net6637));
 sky130_fd_sc_hd__buf_1 fanout6638 (.A(net6641),
    .X(net6638));
 sky130_fd_sc_hd__buf_1 wire6639 (.A(net6640),
    .X(net6639));
 sky130_fd_sc_hd__buf_1 wire6640 (.A(net6638),
    .X(net6640));
 sky130_fd_sc_hd__clkbuf_1 fanout6641 (.A(net6645),
    .X(net6641));
 sky130_fd_sc_hd__clkbuf_1 wire6642 (.A(net6643),
    .X(net6642));
 sky130_fd_sc_hd__buf_1 wire6643 (.A(net6644),
    .X(net6643));
 sky130_fd_sc_hd__clkbuf_2 wire6644 (.A(net6641),
    .X(net6644));
 sky130_fd_sc_hd__clkbuf_1 wire6645 (.A(net6646),
    .X(net6645));
 sky130_fd_sc_hd__clkbuf_1 wire6646 (.A(net6647),
    .X(net6646));
 sky130_fd_sc_hd__clkbuf_1 max_length6647 (.A(net6648),
    .X(net6647));
 sky130_fd_sc_hd__buf_1 wire6648 (.A(\matmul0.matmul_stage_inst.state[1] ),
    .X(net6648));
 sky130_fd_sc_hd__buf_1 wire6649 (.A(net6650),
    .X(net6649));
 sky130_fd_sc_hd__buf_1 wire6650 (.A(net6651),
    .X(net6650));
 sky130_fd_sc_hd__clkbuf_1 wire6651 (.A(net6652),
    .X(net6651));
 sky130_fd_sc_hd__clkbuf_1 wire6652 (.A(net6653),
    .X(net6652));
 sky130_fd_sc_hd__clkbuf_1 wire6653 (.A(net6654),
    .X(net6653));
 sky130_fd_sc_hd__clkbuf_1 wire6654 (.A(net6655),
    .X(net6654));
 sky130_fd_sc_hd__clkbuf_1 wire6655 (.A(\svm0.ready ),
    .X(net6655));
 sky130_fd_sc_hd__buf_1 fanout6656 (.A(net6671),
    .X(net6656));
 sky130_fd_sc_hd__buf_1 wire6657 (.A(net6659),
    .X(net6657));
 sky130_fd_sc_hd__buf_1 wire6658 (.A(net6659),
    .X(net6658));
 sky130_fd_sc_hd__buf_1 wire6659 (.A(net6656),
    .X(net6659));
 sky130_fd_sc_hd__buf_1 fanout6660 (.A(net6671),
    .X(net6660));
 sky130_fd_sc_hd__buf_1 wire6661 (.A(net6662),
    .X(net6661));
 sky130_fd_sc_hd__buf_1 wire6662 (.A(net6660),
    .X(net6662));
 sky130_fd_sc_hd__clkbuf_1 fanout6663 (.A(\svm0.state[2] ),
    .X(net6663));
 sky130_fd_sc_hd__buf_1 wire6664 (.A(net6665),
    .X(net6664));
 sky130_fd_sc_hd__clkbuf_1 wire6665 (.A(net6666),
    .X(net6665));
 sky130_fd_sc_hd__clkbuf_1 wire6666 (.A(net6667),
    .X(net6666));
 sky130_fd_sc_hd__clkbuf_1 wire6667 (.A(net6668),
    .X(net6667));
 sky130_fd_sc_hd__clkbuf_1 wire6668 (.A(net6669),
    .X(net6668));
 sky130_fd_sc_hd__buf_1 wire6669 (.A(net6670),
    .X(net6669));
 sky130_fd_sc_hd__clkbuf_1 wire6670 (.A(net6663),
    .X(net6670));
 sky130_fd_sc_hd__clkbuf_1 max_length6671 (.A(net6663),
    .X(net6671));
 sky130_fd_sc_hd__buf_1 fanout6672 (.A(net6674),
    .X(net6672));
 sky130_fd_sc_hd__clkbuf_2 wire6673 (.A(net6672),
    .X(net6673));
 sky130_fd_sc_hd__clkbuf_1 wire6674 (.A(net6675),
    .X(net6674));
 sky130_fd_sc_hd__clkbuf_1 wire6675 (.A(net6676),
    .X(net6675));
 sky130_fd_sc_hd__clkbuf_1 max_length6676 (.A(\svm0.state[1] ),
    .X(net6676));
 sky130_fd_sc_hd__clkbuf_2 fanout6677 (.A(net6679),
    .X(net6677));
 sky130_fd_sc_hd__clkbuf_2 max_length6678 (.A(net6677),
    .X(net6678));
 sky130_fd_sc_hd__clkbuf_1 wire6679 (.A(net6680),
    .X(net6679));
 sky130_fd_sc_hd__clkbuf_1 wire6680 (.A(net6681),
    .X(net6680));
 sky130_fd_sc_hd__clkbuf_1 wire6681 (.A(\svm0.state[0] ),
    .X(net6681));
 sky130_fd_sc_hd__clkbuf_1 wire6682 (.A(net149),
    .X(net6682));
 sky130_fd_sc_hd__clkbuf_1 wire6683 (.A(net151),
    .X(net6683));
 sky130_fd_sc_hd__buf_1 wire6684 (.A(net6685),
    .X(net6684));
 sky130_fd_sc_hd__clkbuf_2 max_length6685 (.A(\svm0.counter[15] ),
    .X(net6685));
 sky130_fd_sc_hd__clkbuf_2 fanout6686 (.A(\svm0.counter[14] ),
    .X(net6686));
 sky130_fd_sc_hd__buf_1 wire6687 (.A(net6686),
    .X(net6687));
 sky130_fd_sc_hd__buf_1 wire6688 (.A(net6686),
    .X(net6688));
 sky130_fd_sc_hd__buf_1 wire6689 (.A(\svm0.counter[14] ),
    .X(net6689));
 sky130_fd_sc_hd__buf_1 fanout6690 (.A(\svm0.counter[13] ),
    .X(net6690));
 sky130_fd_sc_hd__buf_1 wire6691 (.A(net6692),
    .X(net6691));
 sky130_fd_sc_hd__buf_1 wire6692 (.A(net6690),
    .X(net6692));
 sky130_fd_sc_hd__clkbuf_1 max_length6693 (.A(net6690),
    .X(net6693));
 sky130_fd_sc_hd__clkbuf_2 max_length6694 (.A(net6690),
    .X(net6694));
 sky130_fd_sc_hd__clkbuf_1 wire6695 (.A(net6696),
    .X(net6695));
 sky130_fd_sc_hd__clkbuf_1 wire6696 (.A(\svm0.counter[13] ),
    .X(net6696));
 sky130_fd_sc_hd__buf_1 fanout6697 (.A(\svm0.counter[12] ),
    .X(net6697));
 sky130_fd_sc_hd__buf_1 wire6698 (.A(net6699),
    .X(net6698));
 sky130_fd_sc_hd__buf_1 wire6699 (.A(net6700),
    .X(net6699));
 sky130_fd_sc_hd__clkbuf_1 max_length6700 (.A(net6697),
    .X(net6700));
 sky130_fd_sc_hd__clkbuf_2 wire6701 (.A(net6702),
    .X(net6701));
 sky130_fd_sc_hd__clkbuf_1 max_length6702 (.A(\svm0.counter[12] ),
    .X(net6702));
 sky130_fd_sc_hd__buf_1 wire6703 (.A(net6704),
    .X(net6703));
 sky130_fd_sc_hd__buf_1 wire6704 (.A(\svm0.counter[11] ),
    .X(net6704));
 sky130_fd_sc_hd__buf_1 fanout6705 (.A(\svm0.counter[9] ),
    .X(net6705));
 sky130_fd_sc_hd__buf_1 wire6706 (.A(net6707),
    .X(net6706));
 sky130_fd_sc_hd__buf_1 wire6707 (.A(net6708),
    .X(net6707));
 sky130_fd_sc_hd__buf_1 wire6708 (.A(net6705),
    .X(net6708));
 sky130_fd_sc_hd__clkbuf_1 wire6709 (.A(net6710),
    .X(net6709));
 sky130_fd_sc_hd__buf_1 wire6710 (.A(\svm0.counter[9] ),
    .X(net6710));
 sky130_fd_sc_hd__clkbuf_1 max_length6711 (.A(net6712),
    .X(net6711));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6712 (.A(net6713),
    .X(net6712));
 sky130_fd_sc_hd__clkbuf_1 wire6713 (.A(\svm0.counter[8] ),
    .X(net6713));
 sky130_fd_sc_hd__buf_1 wire6714 (.A(net6715),
    .X(net6714));
 sky130_fd_sc_hd__clkbuf_1 wire6715 (.A(net6716),
    .X(net6715));
 sky130_fd_sc_hd__buf_1 wire6716 (.A(net6717),
    .X(net6716));
 sky130_fd_sc_hd__clkbuf_2 max_length6717 (.A(\svm0.counter[7] ),
    .X(net6717));
 sky130_fd_sc_hd__buf_1 fanout6718 (.A(\svm0.counter[6] ),
    .X(net6718));
 sky130_fd_sc_hd__clkbuf_1 wire6719 (.A(net6724),
    .X(net6719));
 sky130_fd_sc_hd__buf_1 wire6720 (.A(net6721),
    .X(net6720));
 sky130_fd_sc_hd__buf_1 wire6721 (.A(net6722),
    .X(net6721));
 sky130_fd_sc_hd__buf_1 wire6722 (.A(net6723),
    .X(net6722));
 sky130_fd_sc_hd__clkbuf_1 wire6723 (.A(net6724),
    .X(net6723));
 sky130_fd_sc_hd__buf_1 wire6724 (.A(net6718),
    .X(net6724));
 sky130_fd_sc_hd__clkbuf_1 wire6725 (.A(net6726),
    .X(net6725));
 sky130_fd_sc_hd__clkbuf_1 wire6726 (.A(\svm0.counter[6] ),
    .X(net6726));
 sky130_fd_sc_hd__clkbuf_1 wire6727 (.A(net6729),
    .X(net6727));
 sky130_fd_sc_hd__buf_1 wire6728 (.A(\svm0.counter[5] ),
    .X(net6728));
 sky130_fd_sc_hd__buf_1 max_length6729 (.A(\svm0.counter[5] ),
    .X(net6729));
 sky130_fd_sc_hd__clkbuf_1 wire6730 (.A(net6731),
    .X(net6730));
 sky130_fd_sc_hd__clkbuf_1 wire6731 (.A(net6732),
    .X(net6731));
 sky130_fd_sc_hd__buf_1 wire6732 (.A(\svm0.counter[4] ),
    .X(net6732));
 sky130_fd_sc_hd__buf_1 wire6733 (.A(net6734),
    .X(net6733));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6734 (.A(net6735),
    .X(net6734));
 sky130_fd_sc_hd__buf_1 wire6735 (.A(\svm0.counter[2] ),
    .X(net6735));
 sky130_fd_sc_hd__buf_1 wire6736 (.A(\svm0.counter[2] ),
    .X(net6736));
 sky130_fd_sc_hd__buf_1 wire6737 (.A(\svm0.counter[1] ),
    .X(net6737));
 sky130_fd_sc_hd__buf_1 wire6738 (.A(\svm0.counter[1] ),
    .X(net6738));
 sky130_fd_sc_hd__buf_1 wire6739 (.A(net6740),
    .X(net6739));
 sky130_fd_sc_hd__buf_1 wire6740 (.A(net6741),
    .X(net6740));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6741 (.A(\svm0.counter[0] ),
    .X(net6741));
 sky130_fd_sc_hd__clkbuf_2 wire6742 (.A(\svm0.delta[13] ),
    .X(net6742));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6743 (.A(\svm0.delta[2] ),
    .X(net6743));
 sky130_fd_sc_hd__buf_1 max_length6744 (.A(\svm0.delta[1] ),
    .X(net6744));
 sky130_fd_sc_hd__clkbuf_1 wire6745 (.A(\svm0.rising ),
    .X(net6745));
 sky130_fd_sc_hd__buf_1 wire6746 (.A(\svm0.tA[9] ),
    .X(net6746));
 sky130_fd_sc_hd__buf_1 wire6747 (.A(\svm0.tB[13] ),
    .X(net6747));
 sky130_fd_sc_hd__clkbuf_1 wire6748 (.A(net6749),
    .X(net6748));
 sky130_fd_sc_hd__buf_1 wire6749 (.A(net6750),
    .X(net6749));
 sky130_fd_sc_hd__buf_1 wire6750 (.A(net6751),
    .X(net6750));
 sky130_fd_sc_hd__clkbuf_1 wire6751 (.A(net6752),
    .X(net6751));
 sky130_fd_sc_hd__clkbuf_1 wire6752 (.A(net6753),
    .X(net6752));
 sky130_fd_sc_hd__clkbuf_1 wire6753 (.A(net6754),
    .X(net6753));
 sky130_fd_sc_hd__buf_1 wire6754 (.A(\matmul0.state[1] ),
    .X(net6754));
 sky130_fd_sc_hd__buf_1 fanout6755 (.A(net6767),
    .X(net6755));
 sky130_fd_sc_hd__buf_1 wire6756 (.A(net6757),
    .X(net6756));
 sky130_fd_sc_hd__buf_1 wire6757 (.A(net6755),
    .X(net6757));
 sky130_fd_sc_hd__clkbuf_1 wire6758 (.A(net6755),
    .X(net6758));
 sky130_fd_sc_hd__buf_1 fanout6759 (.A(net6768),
    .X(net6759));
 sky130_fd_sc_hd__buf_1 wire6760 (.A(net6761),
    .X(net6760));
 sky130_fd_sc_hd__clkbuf_1 wire6761 (.A(net6764),
    .X(net6761));
 sky130_fd_sc_hd__buf_1 wire6762 (.A(net6763),
    .X(net6762));
 sky130_fd_sc_hd__buf_1 max_length6763 (.A(net6764),
    .X(net6763));
 sky130_fd_sc_hd__buf_1 wire6764 (.A(net6759),
    .X(net6764));
 sky130_fd_sc_hd__clkbuf_1 fanout6765 (.A(\cordic0.vec[1][17] ),
    .X(net6765));
 sky130_fd_sc_hd__buf_1 wire6766 (.A(net6767),
    .X(net6766));
 sky130_fd_sc_hd__buf_1 wire6767 (.A(net6768),
    .X(net6767));
 sky130_fd_sc_hd__buf_1 wire6768 (.A(net6765),
    .X(net6768));
 sky130_fd_sc_hd__buf_1 fanout6769 (.A(net6772),
    .X(net6769));
 sky130_fd_sc_hd__buf_1 wire6770 (.A(net6769),
    .X(net6770));
 sky130_fd_sc_hd__buf_1 wire6771 (.A(net6769),
    .X(net6771));
 sky130_fd_sc_hd__buf_1 fanout6772 (.A(net6787),
    .X(net6772));
 sky130_fd_sc_hd__buf_1 wire6773 (.A(net6774),
    .X(net6773));
 sky130_fd_sc_hd__clkbuf_2 wire6774 (.A(net6775),
    .X(net6774));
 sky130_fd_sc_hd__clkbuf_1 wire6775 (.A(net6776),
    .X(net6775));
 sky130_fd_sc_hd__clkbuf_1 max_length6776 (.A(net6772),
    .X(net6776));
 sky130_fd_sc_hd__clkbuf_1 fanout6777 (.A(net6782),
    .X(net6777));
 sky130_fd_sc_hd__clkbuf_1 max_length6778 (.A(net6779),
    .X(net6778));
 sky130_fd_sc_hd__buf_2 wire6779 (.A(net6777),
    .X(net6779));
 sky130_fd_sc_hd__clkbuf_1 fanout6780 (.A(net6783),
    .X(net6780));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6781 (.A(net6780),
    .X(net6781));
 sky130_fd_sc_hd__buf_1 fanout6782 (.A(net6786),
    .X(net6782));
 sky130_fd_sc_hd__clkbuf_1 wire6783 (.A(net6782),
    .X(net6783));
 sky130_fd_sc_hd__buf_1 wire6784 (.A(net6785),
    .X(net6784));
 sky130_fd_sc_hd__buf_1 wire6785 (.A(net6782),
    .X(net6785));
 sky130_fd_sc_hd__buf_1 wire6786 (.A(net6787),
    .X(net6786));
 sky130_fd_sc_hd__clkbuf_1 wire6787 (.A(\cordic0.vec[1][17] ),
    .X(net6787));
 sky130_fd_sc_hd__buf_1 fanout6788 (.A(net6806),
    .X(net6788));
 sky130_fd_sc_hd__clkbuf_2 wire6789 (.A(net6788),
    .X(net6789));
 sky130_fd_sc_hd__clkbuf_1 wire6790 (.A(net6791),
    .X(net6790));
 sky130_fd_sc_hd__buf_1 wire6791 (.A(net6788),
    .X(net6791));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout6792 (.A(net6797),
    .X(net6792));
 sky130_fd_sc_hd__buf_1 wire6793 (.A(net6792),
    .X(net6793));
 sky130_fd_sc_hd__buf_1 wire6794 (.A(net6792),
    .X(net6794));
 sky130_fd_sc_hd__buf_1 fanout6795 (.A(net6802),
    .X(net6795));
 sky130_fd_sc_hd__clkbuf_4 wire6796 (.A(net6795),
    .X(net6796));
 sky130_fd_sc_hd__buf_1 fanout6797 (.A(net6805),
    .X(net6797));
 sky130_fd_sc_hd__buf_1 max_length6798 (.A(net6799),
    .X(net6798));
 sky130_fd_sc_hd__buf_1 wire6799 (.A(net6801),
    .X(net6799));
 sky130_fd_sc_hd__clkbuf_1 wire6800 (.A(net6801),
    .X(net6800));
 sky130_fd_sc_hd__buf_1 wire6801 (.A(net6797),
    .X(net6801));
 sky130_fd_sc_hd__clkbuf_1 max_length6802 (.A(net6797),
    .X(net6802));
 sky130_fd_sc_hd__clkbuf_1 fanout6803 (.A(\cordic0.vec[1][16] ),
    .X(net6803));
 sky130_fd_sc_hd__buf_1 wire6804 (.A(net6806),
    .X(net6804));
 sky130_fd_sc_hd__clkbuf_1 wire6805 (.A(net6803),
    .X(net6805));
 sky130_fd_sc_hd__buf_1 max_length6806 (.A(net6803),
    .X(net6806));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout6807 (.A(net6821),
    .X(net6807));
 sky130_fd_sc_hd__buf_1 max_length6808 (.A(net6809),
    .X(net6808));
 sky130_fd_sc_hd__clkbuf_2 wire6809 (.A(net6807),
    .X(net6809));
 sky130_fd_sc_hd__buf_1 wire6810 (.A(net6811),
    .X(net6810));
 sky130_fd_sc_hd__clkbuf_2 wire6811 (.A(net6807),
    .X(net6811));
 sky130_fd_sc_hd__buf_1 fanout6812 (.A(net6816),
    .X(net6812));
 sky130_fd_sc_hd__buf_1 wire6813 (.A(net6814),
    .X(net6813));
 sky130_fd_sc_hd__buf_1 wire6814 (.A(net6812),
    .X(net6814));
 sky130_fd_sc_hd__buf_1 fanout6815 (.A(net6822),
    .X(net6815));
 sky130_fd_sc_hd__buf_1 max_length6816 (.A(net6817),
    .X(net6816));
 sky130_fd_sc_hd__clkbuf_2 max_length6817 (.A(net6818),
    .X(net6817));
 sky130_fd_sc_hd__buf_1 wire6818 (.A(net6815),
    .X(net6818));
 sky130_fd_sc_hd__buf_1 fanout6819 (.A(\cordic0.vec[1][15] ),
    .X(net6819));
 sky130_fd_sc_hd__clkbuf_1 max_length6820 (.A(net6821),
    .X(net6820));
 sky130_fd_sc_hd__buf_1 wire6821 (.A(net6822),
    .X(net6821));
 sky130_fd_sc_hd__buf_1 wire6822 (.A(net6819),
    .X(net6822));
 sky130_fd_sc_hd__clkbuf_1 max_length6823 (.A(net6824),
    .X(net6823));
 sky130_fd_sc_hd__buf_1 wire6824 (.A(net6819),
    .X(net6824));
 sky130_fd_sc_hd__clkbuf_2 fanout6825 (.A(net6835),
    .X(net6825));
 sky130_fd_sc_hd__buf_1 max_length6826 (.A(net6827),
    .X(net6826));
 sky130_fd_sc_hd__buf_1 wire6827 (.A(net6825),
    .X(net6827));
 sky130_fd_sc_hd__clkbuf_2 fanout6828 (.A(net6832),
    .X(net6828));
 sky130_fd_sc_hd__buf_1 max_length6829 (.A(net6830),
    .X(net6829));
 sky130_fd_sc_hd__clkbuf_2 max_length6830 (.A(net6828),
    .X(net6830));
 sky130_fd_sc_hd__buf_1 fanout6831 (.A(net6834),
    .X(net6831));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6832 (.A(net6833),
    .X(net6832));
 sky130_fd_sc_hd__clkbuf_2 max_length6833 (.A(net6831),
    .X(net6833));
 sky130_fd_sc_hd__buf_1 fanout6834 (.A(net6849),
    .X(net6834));
 sky130_fd_sc_hd__clkbuf_1 wire6835 (.A(net6836),
    .X(net6835));
 sky130_fd_sc_hd__buf_1 wire6836 (.A(net6838),
    .X(net6836));
 sky130_fd_sc_hd__buf_1 wire6837 (.A(net6838),
    .X(net6837));
 sky130_fd_sc_hd__buf_1 wire6838 (.A(net6834),
    .X(net6838));
 sky130_fd_sc_hd__buf_1 fanout6839 (.A(net6843),
    .X(net6839));
 sky130_fd_sc_hd__buf_1 wire6840 (.A(net6841),
    .X(net6840));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6841 (.A(net6839),
    .X(net6841));
 sky130_fd_sc_hd__clkbuf_2 wire6842 (.A(net6839),
    .X(net6842));
 sky130_fd_sc_hd__clkbuf_1 fanout6843 (.A(\cordic0.vec[1][14] ),
    .X(net6843));
 sky130_fd_sc_hd__buf_1 wire6844 (.A(net6846),
    .X(net6844));
 sky130_fd_sc_hd__buf_1 wire6845 (.A(net6846),
    .X(net6845));
 sky130_fd_sc_hd__buf_1 wire6846 (.A(net6847),
    .X(net6846));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6847 (.A(net6848),
    .X(net6847));
 sky130_fd_sc_hd__clkbuf_1 wire6848 (.A(net6849),
    .X(net6848));
 sky130_fd_sc_hd__buf_1 wire6849 (.A(net6843),
    .X(net6849));
 sky130_fd_sc_hd__clkbuf_2 fanout6850 (.A(\cordic0.vec[1][13] ),
    .X(net6850));
 sky130_fd_sc_hd__buf_1 wire6851 (.A(net6852),
    .X(net6851));
 sky130_fd_sc_hd__clkbuf_2 wire6852 (.A(net6850),
    .X(net6852));
 sky130_fd_sc_hd__buf_1 wire6853 (.A(net6850),
    .X(net6853));
 sky130_fd_sc_hd__buf_1 fanout6854 (.A(net6869),
    .X(net6854));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6855 (.A(net6854),
    .X(net6855));
 sky130_fd_sc_hd__buf_1 wire6856 (.A(net6854),
    .X(net6856));
 sky130_fd_sc_hd__buf_1 max_length6857 (.A(net6854),
    .X(net6857));
 sky130_fd_sc_hd__buf_1 fanout6858 (.A(net6861),
    .X(net6858));
 sky130_fd_sc_hd__buf_1 wire6859 (.A(net6858),
    .X(net6859));
 sky130_fd_sc_hd__clkbuf_2 wire6860 (.A(net6858),
    .X(net6860));
 sky130_fd_sc_hd__clkbuf_1 fanout6861 (.A(net6866),
    .X(net6861));
 sky130_fd_sc_hd__buf_1 wire6862 (.A(net6863),
    .X(net6862));
 sky130_fd_sc_hd__buf_1 wire6863 (.A(net6864),
    .X(net6863));
 sky130_fd_sc_hd__buf_1 wire6864 (.A(net6865),
    .X(net6864));
 sky130_fd_sc_hd__clkbuf_1 max_length6865 (.A(net6861),
    .X(net6865));
 sky130_fd_sc_hd__clkbuf_1 fanout6866 (.A(net6870),
    .X(net6866));
 sky130_fd_sc_hd__clkbuf_2 max_length6867 (.A(net6868),
    .X(net6867));
 sky130_fd_sc_hd__buf_1 wire6868 (.A(net6869),
    .X(net6868));
 sky130_fd_sc_hd__buf_1 wire6869 (.A(net6866),
    .X(net6869));
 sky130_fd_sc_hd__clkbuf_1 wire6870 (.A(\cordic0.vec[1][13] ),
    .X(net6870));
 sky130_fd_sc_hd__clkbuf_1 max_length6871 (.A(\cordic0.vec[1][13] ),
    .X(net6871));
 sky130_fd_sc_hd__buf_2 fanout6872 (.A(net6886),
    .X(net6872));
 sky130_fd_sc_hd__buf_1 wire6873 (.A(net6874),
    .X(net6873));
 sky130_fd_sc_hd__buf_1 wire6874 (.A(net6872),
    .X(net6874));
 sky130_fd_sc_hd__clkbuf_2 wire6875 (.A(net6872),
    .X(net6875));
 sky130_fd_sc_hd__clkbuf_2 fanout6876 (.A(net6878),
    .X(net6876));
 sky130_fd_sc_hd__buf_2 wire6877 (.A(net6876),
    .X(net6877));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout6878 (.A(net6880),
    .X(net6878));
 sky130_fd_sc_hd__clkbuf_1 fanout6879 (.A(net6883),
    .X(net6879));
 sky130_fd_sc_hd__clkbuf_1 max_length6880 (.A(net6882),
    .X(net6880));
 sky130_fd_sc_hd__buf_1 max_length6881 (.A(net6882),
    .X(net6881));
 sky130_fd_sc_hd__buf_1 wire6882 (.A(net6879),
    .X(net6882));
 sky130_fd_sc_hd__clkbuf_1 fanout6883 (.A(net6888),
    .X(net6883));
 sky130_fd_sc_hd__clkbuf_1 max_length6884 (.A(net6885),
    .X(net6884));
 sky130_fd_sc_hd__buf_1 wire6885 (.A(net6886),
    .X(net6885));
 sky130_fd_sc_hd__buf_1 wire6886 (.A(net6883),
    .X(net6886));
 sky130_fd_sc_hd__buf_1 fanout6887 (.A(\cordic0.vec[1][12] ),
    .X(net6887));
 sky130_fd_sc_hd__clkbuf_1 wire6888 (.A(net6889),
    .X(net6888));
 sky130_fd_sc_hd__clkbuf_1 max_length6889 (.A(net6887),
    .X(net6889));
 sky130_fd_sc_hd__buf_1 wire6890 (.A(net6891),
    .X(net6890));
 sky130_fd_sc_hd__clkbuf_2 max_length6891 (.A(net6887),
    .X(net6891));
 sky130_fd_sc_hd__buf_2 fanout6892 (.A(net6899),
    .X(net6892));
 sky130_fd_sc_hd__buf_1 wire6893 (.A(net6894),
    .X(net6893));
 sky130_fd_sc_hd__buf_1 max_length6894 (.A(net6892),
    .X(net6894));
 sky130_fd_sc_hd__buf_1 fanout6895 (.A(net6902),
    .X(net6895));
 sky130_fd_sc_hd__buf_1 wire6896 (.A(net6897),
    .X(net6896));
 sky130_fd_sc_hd__clkbuf_2 wire6897 (.A(net6900),
    .X(net6897));
 sky130_fd_sc_hd__clkbuf_1 wire6898 (.A(net6900),
    .X(net6898));
 sky130_fd_sc_hd__clkbuf_1 max_length6899 (.A(net6900),
    .X(net6899));
 sky130_fd_sc_hd__clkbuf_2 max_length6900 (.A(net6895),
    .X(net6900));
 sky130_fd_sc_hd__clkbuf_2 fanout6901 (.A(net6905),
    .X(net6901));
 sky130_fd_sc_hd__clkbuf_1 wire6902 (.A(net6903),
    .X(net6902));
 sky130_fd_sc_hd__buf_1 wire6903 (.A(net6901),
    .X(net6903));
 sky130_fd_sc_hd__buf_1 wire6904 (.A(net6901),
    .X(net6904));
 sky130_fd_sc_hd__buf_1 fanout6905 (.A(\cordic0.vec[1][11] ),
    .X(net6905));
 sky130_fd_sc_hd__clkbuf_1 wire6906 (.A(net6907),
    .X(net6906));
 sky130_fd_sc_hd__clkbuf_1 wire6907 (.A(net6908),
    .X(net6907));
 sky130_fd_sc_hd__buf_2 wire6908 (.A(net6910),
    .X(net6908));
 sky130_fd_sc_hd__buf_1 wire6909 (.A(net6910),
    .X(net6909));
 sky130_fd_sc_hd__buf_1 wire6910 (.A(net6911),
    .X(net6910));
 sky130_fd_sc_hd__buf_1 wire6911 (.A(net6912),
    .X(net6911));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6912 (.A(net6913),
    .X(net6912));
 sky130_fd_sc_hd__clkbuf_1 wire6913 (.A(net6905),
    .X(net6913));
 sky130_fd_sc_hd__clkbuf_2 fanout6914 (.A(\cordic0.vec[1][10] ),
    .X(net6914));
 sky130_fd_sc_hd__buf_1 max_length6915 (.A(net6916),
    .X(net6915));
 sky130_fd_sc_hd__buf_1 wire6916 (.A(net6914),
    .X(net6916));
 sky130_fd_sc_hd__buf_1 wire6917 (.A(net6914),
    .X(net6917));
 sky130_fd_sc_hd__clkbuf_1 max_length6918 (.A(net6914),
    .X(net6918));
 sky130_fd_sc_hd__clkbuf_2 fanout6919 (.A(net6929),
    .X(net6919));
 sky130_fd_sc_hd__buf_1 wire6920 (.A(net6921),
    .X(net6920));
 sky130_fd_sc_hd__buf_1 wire6921 (.A(net6919),
    .X(net6921));
 sky130_fd_sc_hd__clkbuf_1 wire6922 (.A(net6919),
    .X(net6922));
 sky130_fd_sc_hd__clkbuf_1 fanout6923 (.A(net6931),
    .X(net6923));
 sky130_fd_sc_hd__buf_1 wire6924 (.A(net6926),
    .X(net6924));
 sky130_fd_sc_hd__buf_1 wire6925 (.A(net6927),
    .X(net6925));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length6926 (.A(net6927),
    .X(net6926));
 sky130_fd_sc_hd__buf_1 wire6927 (.A(net6928),
    .X(net6927));
 sky130_fd_sc_hd__clkbuf_1 max_length6928 (.A(net6929),
    .X(net6928));
 sky130_fd_sc_hd__buf_1 wire6929 (.A(net6930),
    .X(net6929));
 sky130_fd_sc_hd__clkbuf_1 max_length6930 (.A(net6923),
    .X(net6930));
 sky130_fd_sc_hd__clkbuf_1 wire6931 (.A(\cordic0.vec[1][10] ),
    .X(net6931));
 sky130_fd_sc_hd__clkbuf_2 fanout6932 (.A(net6936),
    .X(net6932));
 sky130_fd_sc_hd__buf_1 max_length6933 (.A(net6934),
    .X(net6933));
 sky130_fd_sc_hd__buf_1 wire6934 (.A(net6932),
    .X(net6934));
 sky130_fd_sc_hd__clkbuf_1 max_length6935 (.A(net6932),
    .X(net6935));
 sky130_fd_sc_hd__buf_1 fanout6936 (.A(net6939),
    .X(net6936));
 sky130_fd_sc_hd__clkbuf_1 max_length6937 (.A(net6938),
    .X(net6937));
 sky130_fd_sc_hd__buf_1 wire6938 (.A(net6936),
    .X(net6938));
 sky130_fd_sc_hd__clkbuf_1 fanout6939 (.A(\cordic0.vec[1][9] ),
    .X(net6939));
 sky130_fd_sc_hd__buf_1 wire6940 (.A(net6941),
    .X(net6940));
 sky130_fd_sc_hd__buf_1 wire6941 (.A(net6944),
    .X(net6941));
 sky130_fd_sc_hd__clkbuf_1 wire6942 (.A(net6943),
    .X(net6942));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6943 (.A(net6944),
    .X(net6943));
 sky130_fd_sc_hd__buf_1 wire6944 (.A(net6939),
    .X(net6944));
 sky130_fd_sc_hd__buf_1 fanout6945 (.A(net6958),
    .X(net6945));
 sky130_fd_sc_hd__buf_1 wire6946 (.A(net6951),
    .X(net6946));
 sky130_fd_sc_hd__clkbuf_1 max_length6947 (.A(net6948),
    .X(net6947));
 sky130_fd_sc_hd__clkbuf_2 wire6948 (.A(net6951),
    .X(net6948));
 sky130_fd_sc_hd__clkbuf_1 wire6949 (.A(net6950),
    .X(net6949));
 sky130_fd_sc_hd__clkbuf_1 max_length6950 (.A(net6951),
    .X(net6950));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6951 (.A(net6945),
    .X(net6951));
 sky130_fd_sc_hd__clkbuf_1 fanout6952 (.A(net6960),
    .X(net6952));
 sky130_fd_sc_hd__clkbuf_1 wire6953 (.A(net6957),
    .X(net6953));
 sky130_fd_sc_hd__clkbuf_1 wire6954 (.A(net6955),
    .X(net6954));
 sky130_fd_sc_hd__clkbuf_2 wire6955 (.A(net6956),
    .X(net6955));
 sky130_fd_sc_hd__buf_1 wire6956 (.A(net6957),
    .X(net6956));
 sky130_fd_sc_hd__buf_1 max_length6957 (.A(net6952),
    .X(net6957));
 sky130_fd_sc_hd__clkbuf_1 wire6958 (.A(net6959),
    .X(net6958));
 sky130_fd_sc_hd__clkbuf_1 max_length6959 (.A(net6960),
    .X(net6959));
 sky130_fd_sc_hd__buf_1 wire6960 (.A(\cordic0.vec[1][9] ),
    .X(net6960));
 sky130_fd_sc_hd__buf_1 fanout6961 (.A(\cordic0.vec[1][8] ),
    .X(net6961));
 sky130_fd_sc_hd__buf_1 wire6962 (.A(net6961),
    .X(net6962));
 sky130_fd_sc_hd__buf_1 wire6963 (.A(net6964),
    .X(net6963));
 sky130_fd_sc_hd__buf_1 wire6964 (.A(net6965),
    .X(net6964));
 sky130_fd_sc_hd__buf_1 wire6965 (.A(net6969),
    .X(net6965));
 sky130_fd_sc_hd__buf_1 wire6966 (.A(net6968),
    .X(net6966));
 sky130_fd_sc_hd__clkbuf_1 max_length6967 (.A(net6968),
    .X(net6967));
 sky130_fd_sc_hd__buf_1 wire6968 (.A(net6961),
    .X(net6968));
 sky130_fd_sc_hd__clkbuf_1 max_length6969 (.A(net6961),
    .X(net6969));
 sky130_fd_sc_hd__clkbuf_2 fanout6970 (.A(net6980),
    .X(net6970));
 sky130_fd_sc_hd__clkbuf_1 wire6971 (.A(net6972),
    .X(net6971));
 sky130_fd_sc_hd__buf_1 wire6972 (.A(net6970),
    .X(net6972));
 sky130_fd_sc_hd__buf_1 fanout6973 (.A(net6979),
    .X(net6973));
 sky130_fd_sc_hd__clkbuf_2 wire6974 (.A(net6978),
    .X(net6974));
 sky130_fd_sc_hd__buf_1 wire6975 (.A(net6976),
    .X(net6975));
 sky130_fd_sc_hd__clkbuf_2 wire6976 (.A(net6977),
    .X(net6976));
 sky130_fd_sc_hd__clkbuf_1 wire6977 (.A(net6973),
    .X(net6977));
 sky130_fd_sc_hd__buf_1 max_length6978 (.A(net6973),
    .X(net6978));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6979 (.A(net6980),
    .X(net6979));
 sky130_fd_sc_hd__buf_1 wire6980 (.A(\cordic0.vec[1][8] ),
    .X(net6980));
 sky130_fd_sc_hd__clkbuf_2 fanout6981 (.A(net6992),
    .X(net6981));
 sky130_fd_sc_hd__buf_1 wire6982 (.A(net6984),
    .X(net6982));
 sky130_fd_sc_hd__buf_1 wire6983 (.A(net6981),
    .X(net6983));
 sky130_fd_sc_hd__buf_1 max_length6984 (.A(net6981),
    .X(net6984));
 sky130_fd_sc_hd__clkbuf_1 fanout6985 (.A(\cordic0.vec[1][7] ),
    .X(net6985));
 sky130_fd_sc_hd__clkbuf_1 wire6986 (.A(net6987),
    .X(net6986));
 sky130_fd_sc_hd__clkbuf_1 wire6987 (.A(net6989),
    .X(net6987));
 sky130_fd_sc_hd__clkbuf_1 max_length6988 (.A(net6989),
    .X(net6988));
 sky130_fd_sc_hd__buf_2 wire6989 (.A(net6992),
    .X(net6989));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire6990 (.A(net6991),
    .X(net6990));
 sky130_fd_sc_hd__clkbuf_1 wire6991 (.A(net6992),
    .X(net6991));
 sky130_fd_sc_hd__buf_1 wire6992 (.A(net6985),
    .X(net6992));
 sky130_fd_sc_hd__clkbuf_1 fanout6993 (.A(net7001),
    .X(net6993));
 sky130_fd_sc_hd__clkbuf_1 max_length6994 (.A(net6995),
    .X(net6994));
 sky130_fd_sc_hd__buf_1 wire6995 (.A(net6996),
    .X(net6995));
 sky130_fd_sc_hd__clkbuf_4 wire6996 (.A(net6993),
    .X(net6996));
 sky130_fd_sc_hd__buf_1 wire6997 (.A(net6993),
    .X(net6997));
 sky130_fd_sc_hd__clkbuf_2 fanout6998 (.A(net7002),
    .X(net6998));
 sky130_fd_sc_hd__clkbuf_1 wire6999 (.A(net6998),
    .X(net6999));
 sky130_fd_sc_hd__buf_1 wire7000 (.A(net6998),
    .X(net7000));
 sky130_fd_sc_hd__clkbuf_1 wire7001 (.A(net7002),
    .X(net7001));
 sky130_fd_sc_hd__buf_1 wire7002 (.A(net7003),
    .X(net7002));
 sky130_fd_sc_hd__clkbuf_1 wire7003 (.A(\cordic0.vec[1][7] ),
    .X(net7003));
 sky130_fd_sc_hd__clkbuf_2 fanout7004 (.A(\cordic0.vec[1][6] ),
    .X(net7004));
 sky130_fd_sc_hd__buf_1 wire7005 (.A(net7006),
    .X(net7005));
 sky130_fd_sc_hd__buf_1 wire7006 (.A(net7007),
    .X(net7006));
 sky130_fd_sc_hd__buf_1 wire7007 (.A(net7004),
    .X(net7007));
 sky130_fd_sc_hd__buf_1 fanout7008 (.A(net7026),
    .X(net7008));
 sky130_fd_sc_hd__clkbuf_1 wire7009 (.A(net7011),
    .X(net7009));
 sky130_fd_sc_hd__buf_1 wire7010 (.A(net7011),
    .X(net7010));
 sky130_fd_sc_hd__buf_1 wire7011 (.A(net7008),
    .X(net7011));
 sky130_fd_sc_hd__clkbuf_2 fanout7012 (.A(net7018),
    .X(net7012));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7013 (.A(net7012),
    .X(net7013));
 sky130_fd_sc_hd__buf_1 wire7014 (.A(net7012),
    .X(net7014));
 sky130_fd_sc_hd__clkbuf_1 fanout7015 (.A(net7023),
    .X(net7015));
 sky130_fd_sc_hd__buf_1 wire7016 (.A(net7017),
    .X(net7016));
 sky130_fd_sc_hd__buf_1 wire7017 (.A(net7015),
    .X(net7017));
 sky130_fd_sc_hd__clkbuf_1 fanout7018 (.A(net7024),
    .X(net7018));
 sky130_fd_sc_hd__buf_1 wire7019 (.A(net7021),
    .X(net7019));
 sky130_fd_sc_hd__buf_1 wire7020 (.A(net7022),
    .X(net7020));
 sky130_fd_sc_hd__buf_1 max_length7021 (.A(net7022),
    .X(net7021));
 sky130_fd_sc_hd__clkbuf_2 max_length7022 (.A(net7023),
    .X(net7022));
 sky130_fd_sc_hd__buf_1 wire7023 (.A(net7018),
    .X(net7023));
 sky130_fd_sc_hd__clkbuf_1 wire7024 (.A(net7025),
    .X(net7024));
 sky130_fd_sc_hd__clkbuf_1 wire7025 (.A(net7026),
    .X(net7025));
 sky130_fd_sc_hd__buf_1 max_length7026 (.A(\cordic0.vec[1][6] ),
    .X(net7026));
 sky130_fd_sc_hd__buf_2 fanout7027 (.A(net7031),
    .X(net7027));
 sky130_fd_sc_hd__buf_1 wire7028 (.A(net7029),
    .X(net7028));
 sky130_fd_sc_hd__buf_1 max_length7029 (.A(net7027),
    .X(net7029));
 sky130_fd_sc_hd__buf_1 fanout7030 (.A(net7037),
    .X(net7030));
 sky130_fd_sc_hd__buf_1 wire7031 (.A(net7033),
    .X(net7031));
 sky130_fd_sc_hd__buf_2 wire7032 (.A(net7030),
    .X(net7032));
 sky130_fd_sc_hd__buf_1 max_length7033 (.A(net7030),
    .X(net7033));
 sky130_fd_sc_hd__clkbuf_1 fanout7034 (.A(net7049),
    .X(net7034));
 sky130_fd_sc_hd__buf_1 wire7035 (.A(net7038),
    .X(net7035));
 sky130_fd_sc_hd__clkbuf_1 max_length7036 (.A(net7037),
    .X(net7036));
 sky130_fd_sc_hd__buf_1 wire7037 (.A(net7038),
    .X(net7037));
 sky130_fd_sc_hd__clkbuf_2 wire7038 (.A(net7034),
    .X(net7038));
 sky130_fd_sc_hd__clkbuf_2 fanout7039 (.A(\cordic0.vec[1][5] ),
    .X(net7039));
 sky130_fd_sc_hd__buf_1 wire7040 (.A(net7041),
    .X(net7040));
 sky130_fd_sc_hd__buf_1 wire7041 (.A(net7039),
    .X(net7041));
 sky130_fd_sc_hd__buf_1 wire7042 (.A(net7039),
    .X(net7042));
 sky130_fd_sc_hd__buf_1 fanout7043 (.A(net7047),
    .X(net7043));
 sky130_fd_sc_hd__clkbuf_1 wire7044 (.A(net7045),
    .X(net7044));
 sky130_fd_sc_hd__buf_1 wire7045 (.A(net7043),
    .X(net7045));
 sky130_fd_sc_hd__buf_1 wire7046 (.A(net7043),
    .X(net7046));
 sky130_fd_sc_hd__clkbuf_1 wire7047 (.A(net7048),
    .X(net7047));
 sky130_fd_sc_hd__clkbuf_1 wire7048 (.A(net7049),
    .X(net7048));
 sky130_fd_sc_hd__buf_1 max_length7049 (.A(\cordic0.vec[1][5] ),
    .X(net7049));
 sky130_fd_sc_hd__buf_1 fanout7050 (.A(net7055),
    .X(net7050));
 sky130_fd_sc_hd__buf_1 wire7051 (.A(net7052),
    .X(net7051));
 sky130_fd_sc_hd__buf_2 wire7052 (.A(net7050),
    .X(net7052));
 sky130_fd_sc_hd__buf_1 fanout7053 (.A(net7073),
    .X(net7053));
 sky130_fd_sc_hd__clkbuf_1 wire7054 (.A(net7055),
    .X(net7054));
 sky130_fd_sc_hd__buf_1 wire7055 (.A(net7057),
    .X(net7055));
 sky130_fd_sc_hd__buf_1 wire7056 (.A(net7057),
    .X(net7056));
 sky130_fd_sc_hd__clkbuf_2 max_length7057 (.A(net7053),
    .X(net7057));
 sky130_fd_sc_hd__clkbuf_1 fanout7058 (.A(net7062),
    .X(net7058));
 sky130_fd_sc_hd__clkbuf_1 max_length7059 (.A(net7060),
    .X(net7059));
 sky130_fd_sc_hd__buf_1 wire7060 (.A(net7061),
    .X(net7060));
 sky130_fd_sc_hd__clkbuf_2 wire7061 (.A(net7058),
    .X(net7061));
 sky130_fd_sc_hd__buf_1 fanout7062 (.A(net7067),
    .X(net7062));
 sky130_fd_sc_hd__buf_1 wire7063 (.A(net7064),
    .X(net7063));
 sky130_fd_sc_hd__buf_1 wire7064 (.A(net7065),
    .X(net7064));
 sky130_fd_sc_hd__buf_1 wire7065 (.A(net7062),
    .X(net7065));
 sky130_fd_sc_hd__buf_1 fanout7066 (.A(net7077),
    .X(net7066));
 sky130_fd_sc_hd__buf_1 max_length7067 (.A(net7066),
    .X(net7067));
 sky130_fd_sc_hd__clkbuf_1 wire7068 (.A(net7069),
    .X(net7068));
 sky130_fd_sc_hd__buf_1 wire7069 (.A(net7072),
    .X(net7069));
 sky130_fd_sc_hd__clkbuf_1 max_length7070 (.A(net7071),
    .X(net7070));
 sky130_fd_sc_hd__clkbuf_2 max_length7071 (.A(net7072),
    .X(net7071));
 sky130_fd_sc_hd__buf_1 wire7072 (.A(net7066),
    .X(net7072));
 sky130_fd_sc_hd__clkbuf_1 fanout7073 (.A(\cordic0.vec[1][4] ),
    .X(net7073));
 sky130_fd_sc_hd__clkbuf_1 wire7074 (.A(net7079),
    .X(net7074));
 sky130_fd_sc_hd__clkbuf_1 wire7075 (.A(net7077),
    .X(net7075));
 sky130_fd_sc_hd__buf_1 wire7076 (.A(net7077),
    .X(net7076));
 sky130_fd_sc_hd__buf_1 wire7077 (.A(net7078),
    .X(net7077));
 sky130_fd_sc_hd__buf_1 wire7078 (.A(net7079),
    .X(net7078));
 sky130_fd_sc_hd__buf_1 wire7079 (.A(net7073),
    .X(net7079));
 sky130_fd_sc_hd__buf_1 fanout7080 (.A(\cordic0.vec[1][3] ),
    .X(net7080));
 sky130_fd_sc_hd__buf_1 wire7081 (.A(net7083),
    .X(net7081));
 sky130_fd_sc_hd__buf_1 wire7082 (.A(net7083),
    .X(net7082));
 sky130_fd_sc_hd__clkbuf_2 wire7083 (.A(net7084),
    .X(net7083));
 sky130_fd_sc_hd__clkbuf_1 wire7084 (.A(net7085),
    .X(net7084));
 sky130_fd_sc_hd__clkbuf_1 wire7085 (.A(net7080),
    .X(net7085));
 sky130_fd_sc_hd__buf_1 fanout7086 (.A(net7102),
    .X(net7086));
 sky130_fd_sc_hd__clkbuf_1 wire7087 (.A(net7088),
    .X(net7087));
 sky130_fd_sc_hd__buf_1 wire7088 (.A(net7086),
    .X(net7088));
 sky130_fd_sc_hd__buf_1 fanout7089 (.A(net7093),
    .X(net7089));
 sky130_fd_sc_hd__buf_1 max_length7090 (.A(net7091),
    .X(net7090));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7091 (.A(net7089),
    .X(net7091));
 sky130_fd_sc_hd__clkbuf_2 fanout7092 (.A(net7093),
    .X(net7092));
 sky130_fd_sc_hd__buf_1 fanout7093 (.A(net7097),
    .X(net7093));
 sky130_fd_sc_hd__buf_1 wire7094 (.A(net7095),
    .X(net7094));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7095 (.A(net7093),
    .X(net7095));
 sky130_fd_sc_hd__clkbuf_2 fanout7096 (.A(net7100),
    .X(net7096));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7097 (.A(net7096),
    .X(net7097));
 sky130_fd_sc_hd__buf_1 max_length7098 (.A(net7099),
    .X(net7098));
 sky130_fd_sc_hd__buf_1 wire7099 (.A(net7096),
    .X(net7099));
 sky130_fd_sc_hd__clkbuf_1 wire7100 (.A(net7101),
    .X(net7100));
 sky130_fd_sc_hd__clkbuf_1 wire7101 (.A(net7102),
    .X(net7101));
 sky130_fd_sc_hd__buf_1 wire7102 (.A(\cordic0.vec[1][3] ),
    .X(net7102));
 sky130_fd_sc_hd__buf_1 fanout7103 (.A(net7109),
    .X(net7103));
 sky130_fd_sc_hd__buf_1 max_length7104 (.A(net7103),
    .X(net7104));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7105 (.A(net7103),
    .X(net7105));
 sky130_fd_sc_hd__buf_1 fanout7106 (.A(net7117),
    .X(net7106));
 sky130_fd_sc_hd__clkbuf_2 wire7107 (.A(net7108),
    .X(net7107));
 sky130_fd_sc_hd__clkbuf_2 max_length7108 (.A(net7109),
    .X(net7108));
 sky130_fd_sc_hd__buf_1 wire7109 (.A(net7106),
    .X(net7109));
 sky130_fd_sc_hd__buf_1 fanout7110 (.A(net7114),
    .X(net7110));
 sky130_fd_sc_hd__buf_1 max_length7111 (.A(net7112),
    .X(net7111));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7112 (.A(net7110),
    .X(net7112));
 sky130_fd_sc_hd__buf_1 wire7113 (.A(net7110),
    .X(net7113));
 sky130_fd_sc_hd__buf_1 fanout7114 (.A(\cordic0.vec[1][2] ),
    .X(net7114));
 sky130_fd_sc_hd__buf_1 wire7115 (.A(net7116),
    .X(net7115));
 sky130_fd_sc_hd__buf_1 wire7116 (.A(net7117),
    .X(net7116));
 sky130_fd_sc_hd__buf_1 wire7117 (.A(net7114),
    .X(net7117));
 sky130_fd_sc_hd__buf_1 fanout7118 (.A(net7127),
    .X(net7118));
 sky130_fd_sc_hd__buf_1 max_length7119 (.A(net7121),
    .X(net7119));
 sky130_fd_sc_hd__buf_1 max_length7120 (.A(net7121),
    .X(net7120));
 sky130_fd_sc_hd__buf_1 max_length7121 (.A(net7118),
    .X(net7121));
 sky130_fd_sc_hd__clkbuf_1 fanout7122 (.A(net7126),
    .X(net7122));
 sky130_fd_sc_hd__buf_1 wire7123 (.A(net7124),
    .X(net7123));
 sky130_fd_sc_hd__buf_2 wire7124 (.A(net7122),
    .X(net7124));
 sky130_fd_sc_hd__buf_1 fanout7125 (.A(\cordic0.vec[1][1] ),
    .X(net7125));
 sky130_fd_sc_hd__buf_1 wire7126 (.A(net7128),
    .X(net7126));
 sky130_fd_sc_hd__clkbuf_1 max_length7127 (.A(net7128),
    .X(net7127));
 sky130_fd_sc_hd__buf_1 wire7128 (.A(net7125),
    .X(net7128));
 sky130_fd_sc_hd__buf_1 wire7129 (.A(net7125),
    .X(net7129));
 sky130_fd_sc_hd__clkbuf_1 max_length7130 (.A(\cordic0.vec[1][1] ),
    .X(net7130));
 sky130_fd_sc_hd__clkbuf_1 fanout7131 (.A(net7137),
    .X(net7131));
 sky130_fd_sc_hd__buf_1 wire7132 (.A(net7133),
    .X(net7132));
 sky130_fd_sc_hd__clkbuf_4 wire7133 (.A(net7131),
    .X(net7133));
 sky130_fd_sc_hd__buf_1 fanout7134 (.A(net7143),
    .X(net7134));
 sky130_fd_sc_hd__buf_1 max_length7135 (.A(net7136),
    .X(net7135));
 sky130_fd_sc_hd__buf_1 wire7136 (.A(net7137),
    .X(net7136));
 sky130_fd_sc_hd__buf_1 wire7137 (.A(net7134),
    .X(net7137));
 sky130_fd_sc_hd__buf_1 wire7138 (.A(net7134),
    .X(net7138));
 sky130_fd_sc_hd__buf_1 fanout7139 (.A(net7145),
    .X(net7139));
 sky130_fd_sc_hd__buf_1 wire7140 (.A(net7139),
    .X(net7140));
 sky130_fd_sc_hd__buf_1 wire7141 (.A(net7142),
    .X(net7141));
 sky130_fd_sc_hd__clkbuf_2 wire7142 (.A(net7139),
    .X(net7142));
 sky130_fd_sc_hd__buf_1 fanout7143 (.A(\cordic0.vec[1][0] ),
    .X(net7143));
 sky130_fd_sc_hd__buf_1 wire7144 (.A(net7145),
    .X(net7144));
 sky130_fd_sc_hd__buf_1 wire7145 (.A(net7146),
    .X(net7145));
 sky130_fd_sc_hd__buf_1 wire7146 (.A(net7143),
    .X(net7146));
 sky130_fd_sc_hd__buf_1 max_length7147 (.A(net7143),
    .X(net7147));
 sky130_fd_sc_hd__clkbuf_2 wire7148 (.A(\matmul0.sin[13] ),
    .X(net7148));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7149 (.A(net7150),
    .X(net7149));
 sky130_fd_sc_hd__clkbuf_1 max_length7150 (.A(\matmul0.sin[9] ),
    .X(net7150));
 sky130_fd_sc_hd__buf_1 wire7151 (.A(\matmul0.sin[8] ),
    .X(net7151));
 sky130_fd_sc_hd__clkbuf_2 wire7152 (.A(\matmul0.sin[7] ),
    .X(net7152));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7153 (.A(net7154),
    .X(net7153));
 sky130_fd_sc_hd__clkbuf_1 max_length7154 (.A(\matmul0.sin[6] ),
    .X(net7154));
 sky130_fd_sc_hd__buf_1 wire7155 (.A(\matmul0.sin[5] ),
    .X(net7155));
 sky130_fd_sc_hd__buf_1 wire7156 (.A(net7157),
    .X(net7156));
 sky130_fd_sc_hd__clkbuf_1 max_length7157 (.A(\matmul0.sin[3] ),
    .X(net7157));
 sky130_fd_sc_hd__clkbuf_2 wire7158 (.A(net7159),
    .X(net7158));
 sky130_fd_sc_hd__buf_1 wire7159 (.A(\matmul0.sin[2] ),
    .X(net7159));
 sky130_fd_sc_hd__clkbuf_2 wire7160 (.A(net7161),
    .X(net7160));
 sky130_fd_sc_hd__buf_1 wire7161 (.A(\matmul0.sin[1] ),
    .X(net7161));
 sky130_fd_sc_hd__clkbuf_1 wire7162 (.A(net7163),
    .X(net7162));
 sky130_fd_sc_hd__buf_1 wire7163 (.A(net7164),
    .X(net7163));
 sky130_fd_sc_hd__buf_1 wire7164 (.A(net7165),
    .X(net7164));
 sky130_fd_sc_hd__clkbuf_1 wire7165 (.A(\matmul0.sin[0] ),
    .X(net7165));
 sky130_fd_sc_hd__buf_1 wire7166 (.A(\matmul0.cos[13] ),
    .X(net7166));
 sky130_fd_sc_hd__buf_1 wire7167 (.A(\matmul0.cos[12] ),
    .X(net7167));
 sky130_fd_sc_hd__buf_1 wire7168 (.A(\matmul0.cos[11] ),
    .X(net7168));
 sky130_fd_sc_hd__buf_1 wire7169 (.A(\matmul0.cos[10] ),
    .X(net7169));
 sky130_fd_sc_hd__buf_1 wire7170 (.A(net7171),
    .X(net7170));
 sky130_fd_sc_hd__clkbuf_1 wire7171 (.A(\matmul0.cos[9] ),
    .X(net7171));
 sky130_fd_sc_hd__buf_1 wire7172 (.A(net7173),
    .X(net7172));
 sky130_fd_sc_hd__clkbuf_1 wire7173 (.A(net7174),
    .X(net7173));
 sky130_fd_sc_hd__clkbuf_1 wire7174 (.A(\matmul0.cos[8] ),
    .X(net7174));
 sky130_fd_sc_hd__clkbuf_1 wire7175 (.A(net7176),
    .X(net7175));
 sky130_fd_sc_hd__clkbuf_1 wire7176 (.A(net7177),
    .X(net7176));
 sky130_fd_sc_hd__clkbuf_1 wire7177 (.A(\matmul0.cos[7] ),
    .X(net7177));
 sky130_fd_sc_hd__clkbuf_1 wire7178 (.A(net7179),
    .X(net7178));
 sky130_fd_sc_hd__clkbuf_1 wire7179 (.A(\matmul0.cos[5] ),
    .X(net7179));
 sky130_fd_sc_hd__clkbuf_1 max_length7180 (.A(\matmul0.cos[4] ),
    .X(net7180));
 sky130_fd_sc_hd__buf_1 wire7181 (.A(\matmul0.cos[2] ),
    .X(net7181));
 sky130_fd_sc_hd__buf_1 wire7182 (.A(\matmul0.cos[1] ),
    .X(net7182));
 sky130_fd_sc_hd__clkbuf_1 wire7183 (.A(\matmul0.a[0] ),
    .X(net7183));
 sky130_fd_sc_hd__clkbuf_1 max_length7184 (.A(\matmul0.b[8] ),
    .X(net7184));
 sky130_fd_sc_hd__clkbuf_1 wire7185 (.A(\matmul0.b[7] ),
    .X(net7185));
 sky130_fd_sc_hd__clkbuf_1 wire7186 (.A(\matmul0.b[4] ),
    .X(net7186));
 sky130_fd_sc_hd__clkbuf_1 wire7187 (.A(\matmul0.b[3] ),
    .X(net7187));
 sky130_fd_sc_hd__clkbuf_1 wire7188 (.A(net7189),
    .X(net7188));
 sky130_fd_sc_hd__clkbuf_1 wire7189 (.A(\matmul0.b[2] ),
    .X(net7189));
 sky130_fd_sc_hd__clkbuf_1 wire7190 (.A(net7191),
    .X(net7190));
 sky130_fd_sc_hd__clkbuf_1 max_length7191 (.A(\matmul0.b[1] ),
    .X(net7191));
 sky130_fd_sc_hd__buf_1 wire7192 (.A(net7193),
    .X(net7192));
 sky130_fd_sc_hd__clkbuf_1 wire7193 (.A(net7194),
    .X(net7193));
 sky130_fd_sc_hd__clkbuf_1 wire7194 (.A(net7195),
    .X(net7194));
 sky130_fd_sc_hd__clkbuf_1 wire7195 (.A(net7196),
    .X(net7195));
 sky130_fd_sc_hd__clkbuf_1 wire7196 (.A(net7197),
    .X(net7196));
 sky130_fd_sc_hd__clkbuf_1 wire7197 (.A(\matmul0.alpha_pass[15] ),
    .X(net7197));
 sky130_fd_sc_hd__clkbuf_1 wire7198 (.A(net7201),
    .X(net7198));
 sky130_fd_sc_hd__buf_1 wire7199 (.A(net7200),
    .X(net7199));
 sky130_fd_sc_hd__clkbuf_1 wire7200 (.A(net7202),
    .X(net7200));
 sky130_fd_sc_hd__clkbuf_1 max_length7201 (.A(net7202),
    .X(net7201));
 sky130_fd_sc_hd__buf_1 wire7202 (.A(\matmul0.alpha_pass[15] ),
    .X(net7202));
 sky130_fd_sc_hd__buf_1 wire7203 (.A(net7204),
    .X(net7203));
 sky130_fd_sc_hd__clkbuf_1 wire7204 (.A(net7205),
    .X(net7204));
 sky130_fd_sc_hd__clkbuf_1 wire7205 (.A(net7206),
    .X(net7205));
 sky130_fd_sc_hd__clkbuf_1 wire7206 (.A(net7207),
    .X(net7206));
 sky130_fd_sc_hd__clkbuf_1 wire7207 (.A(net7213),
    .X(net7207));
 sky130_fd_sc_hd__clkbuf_1 wire7208 (.A(net7209),
    .X(net7208));
 sky130_fd_sc_hd__buf_1 wire7209 (.A(net7211),
    .X(net7209));
 sky130_fd_sc_hd__clkbuf_1 wire7210 (.A(net7212),
    .X(net7210));
 sky130_fd_sc_hd__clkbuf_1 max_length7211 (.A(net7212),
    .X(net7211));
 sky130_fd_sc_hd__buf_1 wire7212 (.A(net7213),
    .X(net7212));
 sky130_fd_sc_hd__buf_1 wire7213 (.A(\matmul0.alpha_pass[14] ),
    .X(net7213));
 sky130_fd_sc_hd__clkbuf_2 wire7214 (.A(net7215),
    .X(net7214));
 sky130_fd_sc_hd__buf_1 wire7215 (.A(net7216),
    .X(net7215));
 sky130_fd_sc_hd__clkbuf_1 wire7216 (.A(net7217),
    .X(net7216));
 sky130_fd_sc_hd__clkbuf_1 wire7217 (.A(\matmul0.alpha_pass[13] ),
    .X(net7217));
 sky130_fd_sc_hd__buf_1 wire7218 (.A(net7219),
    .X(net7218));
 sky130_fd_sc_hd__clkbuf_1 wire7219 (.A(net7220),
    .X(net7219));
 sky130_fd_sc_hd__clkbuf_1 wire7220 (.A(net7221),
    .X(net7220));
 sky130_fd_sc_hd__clkbuf_1 wire7221 (.A(net7222),
    .X(net7221));
 sky130_fd_sc_hd__clkbuf_1 wire7222 (.A(net7223),
    .X(net7222));
 sky130_fd_sc_hd__clkbuf_1 wire7223 (.A(net7224),
    .X(net7223));
 sky130_fd_sc_hd__buf_1 max_length7224 (.A(\matmul0.alpha_pass[13] ),
    .X(net7224));
 sky130_fd_sc_hd__clkbuf_1 wire7225 (.A(net7226),
    .X(net7225));
 sky130_fd_sc_hd__clkbuf_1 wire7226 (.A(\matmul0.alpha_pass[12] ),
    .X(net7226));
 sky130_fd_sc_hd__buf_1 wire7227 (.A(net7228),
    .X(net7227));
 sky130_fd_sc_hd__clkbuf_1 wire7228 (.A(net7229),
    .X(net7228));
 sky130_fd_sc_hd__clkbuf_1 wire7229 (.A(net7230),
    .X(net7229));
 sky130_fd_sc_hd__clkbuf_1 wire7230 (.A(net7231),
    .X(net7230));
 sky130_fd_sc_hd__clkbuf_1 wire7231 (.A(net7236),
    .X(net7231));
 sky130_fd_sc_hd__clkbuf_1 wire7232 (.A(net7233),
    .X(net7232));
 sky130_fd_sc_hd__buf_1 wire7233 (.A(net7234),
    .X(net7233));
 sky130_fd_sc_hd__buf_1 wire7234 (.A(net7235),
    .X(net7234));
 sky130_fd_sc_hd__clkbuf_1 wire7235 (.A(net7236),
    .X(net7235));
 sky130_fd_sc_hd__buf_1 wire7236 (.A(\matmul0.alpha_pass[12] ),
    .X(net7236));
 sky130_fd_sc_hd__clkbuf_2 wire7237 (.A(net7238),
    .X(net7237));
 sky130_fd_sc_hd__clkbuf_1 wire7238 (.A(net7239),
    .X(net7238));
 sky130_fd_sc_hd__clkbuf_1 wire7239 (.A(net7240),
    .X(net7239));
 sky130_fd_sc_hd__clkbuf_1 wire7240 (.A(net7241),
    .X(net7240));
 sky130_fd_sc_hd__clkbuf_1 wire7241 (.A(net7242),
    .X(net7241));
 sky130_fd_sc_hd__clkbuf_1 wire7242 (.A(net7243),
    .X(net7242));
 sky130_fd_sc_hd__clkbuf_1 wire7243 (.A(net7248),
    .X(net7243));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7244 (.A(net7245),
    .X(net7244));
 sky130_fd_sc_hd__clkbuf_1 max_length7245 (.A(net7246),
    .X(net7245));
 sky130_fd_sc_hd__buf_1 wire7246 (.A(net7247),
    .X(net7246));
 sky130_fd_sc_hd__clkbuf_1 max_length7247 (.A(net7248),
    .X(net7247));
 sky130_fd_sc_hd__buf_1 wire7248 (.A(\matmul0.alpha_pass[11] ),
    .X(net7248));
 sky130_fd_sc_hd__clkbuf_1 fanout7249 (.A(net7262),
    .X(net7249));
 sky130_fd_sc_hd__clkbuf_2 wire7250 (.A(net7251),
    .X(net7250));
 sky130_fd_sc_hd__clkbuf_1 wire7251 (.A(net7252),
    .X(net7251));
 sky130_fd_sc_hd__clkbuf_1 wire7252 (.A(net7253),
    .X(net7252));
 sky130_fd_sc_hd__clkbuf_1 wire7253 (.A(net7254),
    .X(net7253));
 sky130_fd_sc_hd__clkbuf_1 wire7254 (.A(net7255),
    .X(net7254));
 sky130_fd_sc_hd__clkbuf_1 wire7255 (.A(net7259),
    .X(net7255));
 sky130_fd_sc_hd__clkbuf_1 wire7256 (.A(net7258),
    .X(net7256));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7257 (.A(net7258),
    .X(net7257));
 sky130_fd_sc_hd__buf_1 wire7258 (.A(net7249),
    .X(net7258));
 sky130_fd_sc_hd__buf_1 max_length7259 (.A(net7249),
    .X(net7259));
 sky130_fd_sc_hd__buf_1 wire7260 (.A(net7261),
    .X(net7260));
 sky130_fd_sc_hd__clkbuf_1 wire7261 (.A(net7262),
    .X(net7261));
 sky130_fd_sc_hd__buf_1 wire7262 (.A(net7263),
    .X(net7262));
 sky130_fd_sc_hd__clkbuf_1 wire7263 (.A(\matmul0.alpha_pass[10] ),
    .X(net7263));
 sky130_fd_sc_hd__clkbuf_2 wire7264 (.A(net7270),
    .X(net7264));
 sky130_fd_sc_hd__buf_1 wire7265 (.A(net7266),
    .X(net7265));
 sky130_fd_sc_hd__clkbuf_1 wire7266 (.A(net7267),
    .X(net7266));
 sky130_fd_sc_hd__clkbuf_1 wire7267 (.A(net7268),
    .X(net7267));
 sky130_fd_sc_hd__clkbuf_1 wire7268 (.A(net7269),
    .X(net7268));
 sky130_fd_sc_hd__clkbuf_1 wire7269 (.A(net7270),
    .X(net7269));
 sky130_fd_sc_hd__buf_1 wire7270 (.A(net7271),
    .X(net7270));
 sky130_fd_sc_hd__buf_1 wire7271 (.A(net7274),
    .X(net7271));
 sky130_fd_sc_hd__clkbuf_1 wire7272 (.A(net7273),
    .X(net7272));
 sky130_fd_sc_hd__clkbuf_1 max_length7273 (.A(net7274),
    .X(net7273));
 sky130_fd_sc_hd__buf_1 max_length7274 (.A(\matmul0.alpha_pass[9] ),
    .X(net7274));
 sky130_fd_sc_hd__clkbuf_1 wire7275 (.A(net7276),
    .X(net7275));
 sky130_fd_sc_hd__clkbuf_1 wire7276 (.A(net7277),
    .X(net7276));
 sky130_fd_sc_hd__clkbuf_1 wire7277 (.A(\matmul0.alpha_pass[8] ),
    .X(net7277));
 sky130_fd_sc_hd__clkbuf_2 wire7278 (.A(net7279),
    .X(net7278));
 sky130_fd_sc_hd__buf_1 max_length7279 (.A(net7280),
    .X(net7279));
 sky130_fd_sc_hd__buf_1 wire7280 (.A(net7281),
    .X(net7280));
 sky130_fd_sc_hd__buf_1 wire7281 (.A(\matmul0.alpha_pass[8] ),
    .X(net7281));
 sky130_fd_sc_hd__buf_1 wire7282 (.A(net7283),
    .X(net7282));
 sky130_fd_sc_hd__buf_1 wire7283 (.A(net7284),
    .X(net7283));
 sky130_fd_sc_hd__buf_1 wire7284 (.A(net7285),
    .X(net7284));
 sky130_fd_sc_hd__clkbuf_1 wire7285 (.A(net7286),
    .X(net7285));
 sky130_fd_sc_hd__clkbuf_1 wire7286 (.A(\matmul0.alpha_pass[7] ),
    .X(net7286));
 sky130_fd_sc_hd__buf_1 wire7287 (.A(net7288),
    .X(net7287));
 sky130_fd_sc_hd__clkbuf_1 wire7288 (.A(net7289),
    .X(net7288));
 sky130_fd_sc_hd__clkbuf_1 wire7289 (.A(net7290),
    .X(net7289));
 sky130_fd_sc_hd__clkbuf_1 wire7290 (.A(net7291),
    .X(net7290));
 sky130_fd_sc_hd__buf_1 wire7291 (.A(net7292),
    .X(net7291));
 sky130_fd_sc_hd__clkbuf_1 wire7292 (.A(net7293),
    .X(net7292));
 sky130_fd_sc_hd__clkbuf_1 wire7293 (.A(\matmul0.alpha_pass[7] ),
    .X(net7293));
 sky130_fd_sc_hd__buf_1 wire7294 (.A(net7295),
    .X(net7294));
 sky130_fd_sc_hd__clkbuf_1 wire7295 (.A(net7296),
    .X(net7295));
 sky130_fd_sc_hd__clkbuf_1 wire7296 (.A(net7297),
    .X(net7296));
 sky130_fd_sc_hd__clkbuf_1 wire7297 (.A(net7298),
    .X(net7297));
 sky130_fd_sc_hd__clkbuf_1 wire7298 (.A(net7299),
    .X(net7298));
 sky130_fd_sc_hd__buf_1 wire7299 (.A(net7300),
    .X(net7299));
 sky130_fd_sc_hd__clkbuf_1 wire7300 (.A(net7301),
    .X(net7300));
 sky130_fd_sc_hd__clkbuf_1 wire7301 (.A(\matmul0.alpha_pass[6] ),
    .X(net7301));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7302 (.A(net7303),
    .X(net7302));
 sky130_fd_sc_hd__buf_1 wire7303 (.A(net7304),
    .X(net7303));
 sky130_fd_sc_hd__clkbuf_1 wire7304 (.A(net7305),
    .X(net7304));
 sky130_fd_sc_hd__clkbuf_1 max_length7305 (.A(\matmul0.alpha_pass[6] ),
    .X(net7305));
 sky130_fd_sc_hd__buf_1 wire7306 (.A(net7307),
    .X(net7306));
 sky130_fd_sc_hd__clkbuf_1 wire7307 (.A(net7308),
    .X(net7307));
 sky130_fd_sc_hd__clkbuf_1 wire7308 (.A(net7309),
    .X(net7308));
 sky130_fd_sc_hd__buf_1 wire7309 (.A(net7310),
    .X(net7309));
 sky130_fd_sc_hd__clkbuf_1 wire7310 (.A(net7311),
    .X(net7310));
 sky130_fd_sc_hd__clkbuf_1 wire7311 (.A(net7312),
    .X(net7311));
 sky130_fd_sc_hd__clkbuf_1 wire7312 (.A(net7316),
    .X(net7312));
 sky130_fd_sc_hd__clkbuf_2 wire7313 (.A(net7314),
    .X(net7313));
 sky130_fd_sc_hd__buf_1 wire7314 (.A(net7315),
    .X(net7314));
 sky130_fd_sc_hd__clkbuf_1 wire7315 (.A(\matmul0.alpha_pass[5] ),
    .X(net7315));
 sky130_fd_sc_hd__clkbuf_1 max_length7316 (.A(\matmul0.alpha_pass[5] ),
    .X(net7316));
 sky130_fd_sc_hd__buf_1 wire7317 (.A(net7318),
    .X(net7317));
 sky130_fd_sc_hd__clkbuf_1 wire7318 (.A(net7319),
    .X(net7318));
 sky130_fd_sc_hd__clkbuf_1 wire7319 (.A(net7320),
    .X(net7319));
 sky130_fd_sc_hd__buf_1 wire7320 (.A(net7321),
    .X(net7320));
 sky130_fd_sc_hd__clkbuf_1 wire7321 (.A(net7322),
    .X(net7321));
 sky130_fd_sc_hd__clkbuf_1 wire7322 (.A(net7323),
    .X(net7322));
 sky130_fd_sc_hd__clkbuf_1 wire7323 (.A(net7328),
    .X(net7323));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7324 (.A(net7325),
    .X(net7324));
 sky130_fd_sc_hd__buf_1 wire7325 (.A(net7326),
    .X(net7325));
 sky130_fd_sc_hd__clkbuf_1 wire7326 (.A(net7327),
    .X(net7326));
 sky130_fd_sc_hd__clkbuf_1 wire7327 (.A(\matmul0.alpha_pass[4] ),
    .X(net7327));
 sky130_fd_sc_hd__clkbuf_1 max_length7328 (.A(\matmul0.alpha_pass[4] ),
    .X(net7328));
 sky130_fd_sc_hd__buf_1 wire7329 (.A(net7330),
    .X(net7329));
 sky130_fd_sc_hd__clkbuf_1 wire7330 (.A(net7331),
    .X(net7330));
 sky130_fd_sc_hd__clkbuf_1 wire7331 (.A(net7332),
    .X(net7331));
 sky130_fd_sc_hd__buf_1 wire7332 (.A(net7333),
    .X(net7332));
 sky130_fd_sc_hd__clkbuf_1 wire7333 (.A(net7334),
    .X(net7333));
 sky130_fd_sc_hd__clkbuf_1 wire7334 (.A(net7335),
    .X(net7334));
 sky130_fd_sc_hd__clkbuf_1 wire7335 (.A(\matmul0.alpha_pass[3] ),
    .X(net7335));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7336 (.A(net7337),
    .X(net7336));
 sky130_fd_sc_hd__buf_1 wire7337 (.A(net7338),
    .X(net7337));
 sky130_fd_sc_hd__clkbuf_1 wire7338 (.A(net7339),
    .X(net7338));
 sky130_fd_sc_hd__clkbuf_1 wire7339 (.A(\matmul0.alpha_pass[3] ),
    .X(net7339));
 sky130_fd_sc_hd__buf_1 wire7340 (.A(net7341),
    .X(net7340));
 sky130_fd_sc_hd__buf_1 wire7341 (.A(net7342),
    .X(net7341));
 sky130_fd_sc_hd__clkbuf_1 wire7342 (.A(net7351),
    .X(net7342));
 sky130_fd_sc_hd__buf_1 wire7343 (.A(net7344),
    .X(net7343));
 sky130_fd_sc_hd__clkbuf_1 wire7344 (.A(net7345),
    .X(net7344));
 sky130_fd_sc_hd__clkbuf_1 wire7345 (.A(net7346),
    .X(net7345));
 sky130_fd_sc_hd__buf_1 wire7346 (.A(net7347),
    .X(net7346));
 sky130_fd_sc_hd__clkbuf_1 wire7347 (.A(net7348),
    .X(net7347));
 sky130_fd_sc_hd__clkbuf_1 wire7348 (.A(net7349),
    .X(net7348));
 sky130_fd_sc_hd__clkbuf_1 wire7349 (.A(net7350),
    .X(net7349));
 sky130_fd_sc_hd__clkbuf_1 wire7350 (.A(net7351),
    .X(net7350));
 sky130_fd_sc_hd__buf_1 wire7351 (.A(\matmul0.alpha_pass[2] ),
    .X(net7351));
 sky130_fd_sc_hd__clkbuf_1 max_length7352 (.A(net7353),
    .X(net7352));
 sky130_fd_sc_hd__buf_1 wire7353 (.A(net7354),
    .X(net7353));
 sky130_fd_sc_hd__clkbuf_1 wire7354 (.A(net7355),
    .X(net7354));
 sky130_fd_sc_hd__clkbuf_1 max_length7355 (.A(net7356),
    .X(net7355));
 sky130_fd_sc_hd__buf_1 wire7356 (.A(net7357),
    .X(net7356));
 sky130_fd_sc_hd__clkbuf_1 wire7357 (.A(net7358),
    .X(net7357));
 sky130_fd_sc_hd__clkbuf_1 wire7358 (.A(net7359),
    .X(net7358));
 sky130_fd_sc_hd__clkbuf_1 wire7359 (.A(net7360),
    .X(net7359));
 sky130_fd_sc_hd__clkbuf_1 wire7360 (.A(\matmul0.alpha_pass[1] ),
    .X(net7360));
 sky130_fd_sc_hd__buf_1 max_length7361 (.A(net7362),
    .X(net7361));
 sky130_fd_sc_hd__buf_1 wire7362 (.A(net7363),
    .X(net7362));
 sky130_fd_sc_hd__clkbuf_1 wire7363 (.A(\matmul0.alpha_pass[1] ),
    .X(net7363));
 sky130_fd_sc_hd__buf_1 wire7364 (.A(net7365),
    .X(net7364));
 sky130_fd_sc_hd__buf_1 wire7365 (.A(net7366),
    .X(net7365));
 sky130_fd_sc_hd__clkbuf_1 wire7366 (.A(net7367),
    .X(net7366));
 sky130_fd_sc_hd__clkbuf_1 wire7367 (.A(net7374),
    .X(net7367));
 sky130_fd_sc_hd__buf_1 wire7368 (.A(net7369),
    .X(net7368));
 sky130_fd_sc_hd__buf_1 wire7369 (.A(net7370),
    .X(net7369));
 sky130_fd_sc_hd__clkbuf_1 wire7370 (.A(net7371),
    .X(net7370));
 sky130_fd_sc_hd__clkbuf_1 wire7371 (.A(net7372),
    .X(net7371));
 sky130_fd_sc_hd__clkbuf_1 wire7372 (.A(net7373),
    .X(net7372));
 sky130_fd_sc_hd__buf_1 wire7373 (.A(\matmul0.alpha_pass[0] ),
    .X(net7373));
 sky130_fd_sc_hd__clkbuf_1 max_length7374 (.A(\matmul0.alpha_pass[0] ),
    .X(net7374));
 sky130_fd_sc_hd__buf_1 max_length7375 (.A(\matmul0.matmul_stage_inst.mult2[13] ),
    .X(net7375));
 sky130_fd_sc_hd__buf_1 wire7376 (.A(net7377),
    .X(net7376));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length7377 (.A(\svm0.delta[0] ),
    .X(net7377));
 sky130_fd_sc_hd__buf_1 wire7378 (.A(net7379),
    .X(net7378));
 sky130_fd_sc_hd__clkbuf_1 max_length7379 (.A(\matmul0.matmul_stage_inst.f[15] ),
    .X(net7379));
 sky130_fd_sc_hd__clkbuf_1 wire7380 (.A(\matmul0.matmul_stage_inst.f[14] ),
    .X(net7380));
 sky130_fd_sc_hd__clkbuf_1 wire7381 (.A(\matmul0.matmul_stage_inst.f[12] ),
    .X(net7381));
 sky130_fd_sc_hd__buf_1 max_length7382 (.A(\matmul0.matmul_stage_inst.f[11] ),
    .X(net7382));
 sky130_fd_sc_hd__clkbuf_1 max_length7383 (.A(\matmul0.matmul_stage_inst.f[10] ),
    .X(net7383));
 sky130_fd_sc_hd__clkbuf_1 wire7384 (.A(\matmul0.matmul_stage_inst.f[6] ),
    .X(net7384));
 sky130_fd_sc_hd__clkbuf_1 wire7385 (.A(\matmul0.matmul_stage_inst.f[5] ),
    .X(net7385));
 sky130_fd_sc_hd__clkbuf_1 wire7386 (.A(net7387),
    .X(net7386));
 sky130_fd_sc_hd__clkbuf_1 wire7387 (.A(net7388),
    .X(net7387));
 sky130_fd_sc_hd__clkbuf_1 max_length7388 (.A(\matmul0.matmul_stage_inst.e[10] ),
    .X(net7388));
 sky130_fd_sc_hd__clkbuf_1 wire7389 (.A(net7390),
    .X(net7389));
 sky130_fd_sc_hd__clkbuf_1 max_length7390 (.A(\matmul0.matmul_stage_inst.e[9] ),
    .X(net7390));
 sky130_fd_sc_hd__clkbuf_1 wire7391 (.A(\matmul0.matmul_stage_inst.e[8] ),
    .X(net7391));
 sky130_fd_sc_hd__clkbuf_1 wire7392 (.A(net7393),
    .X(net7392));
 sky130_fd_sc_hd__clkbuf_1 wire7393 (.A(net7394),
    .X(net7393));
 sky130_fd_sc_hd__clkbuf_1 wire7394 (.A(net7395),
    .X(net7394));
 sky130_fd_sc_hd__clkbuf_1 max_length7395 (.A(\matmul0.matmul_stage_inst.e[4] ),
    .X(net7395));
 sky130_fd_sc_hd__clkbuf_1 wire7396 (.A(net7397),
    .X(net7396));
 sky130_fd_sc_hd__clkbuf_1 max_length7397 (.A(\matmul0.matmul_stage_inst.e[2] ),
    .X(net7397));
 sky130_fd_sc_hd__clkbuf_1 wire7398 (.A(net7399),
    .X(net7398));
 sky130_fd_sc_hd__clkbuf_1 wire7399 (.A(net7400),
    .X(net7399));
 sky130_fd_sc_hd__clkbuf_1 max_length7400 (.A(\matmul0.matmul_stage_inst.e[1] ),
    .X(net7400));
 sky130_fd_sc_hd__clkbuf_1 wire7401 (.A(net7402),
    .X(net7401));
 sky130_fd_sc_hd__clkbuf_1 wire7402 (.A(net7403),
    .X(net7402));
 sky130_fd_sc_hd__clkbuf_1 wire7403 (.A(\matmul0.matmul_stage_inst.a[14] ),
    .X(net7403));
 sky130_fd_sc_hd__clkbuf_1 wire7404 (.A(\matmul0.matmul_stage_inst.a[3] ),
    .X(net7404));
 sky130_fd_sc_hd__clkbuf_1 wire7405 (.A(\matmul0.matmul_stage_inst.c[11] ),
    .X(net7405));
 sky130_fd_sc_hd__clkbuf_1 wire7406 (.A(net7407),
    .X(net7406));
 sky130_fd_sc_hd__clkbuf_1 max_length7407 (.A(\matmul0.matmul_stage_inst.c[10] ),
    .X(net7407));
 sky130_fd_sc_hd__clkbuf_1 wire7408 (.A(net7409),
    .X(net7408));
 sky130_fd_sc_hd__clkbuf_1 max_length7409 (.A(\matmul0.matmul_stage_inst.c[9] ),
    .X(net7409));
 sky130_fd_sc_hd__clkbuf_1 wire7410 (.A(\matmul0.matmul_stage_inst.c[8] ),
    .X(net7410));
 sky130_fd_sc_hd__clkbuf_1 wire7411 (.A(net7412),
    .X(net7411));
 sky130_fd_sc_hd__clkbuf_1 wire7412 (.A(\matmul0.matmul_stage_inst.c[6] ),
    .X(net7412));
 sky130_fd_sc_hd__clkbuf_1 wire7413 (.A(\matmul0.matmul_stage_inst.c[5] ),
    .X(net7413));
 sky130_fd_sc_hd__clkbuf_1 wire7414 (.A(net7415),
    .X(net7414));
 sky130_fd_sc_hd__clkbuf_1 wire7415 (.A(net7416),
    .X(net7415));
 sky130_fd_sc_hd__clkbuf_1 wire7416 (.A(\matmul0.matmul_stage_inst.c[4] ),
    .X(net7416));
 sky130_fd_sc_hd__clkbuf_1 wire7417 (.A(\matmul0.matmul_stage_inst.c[2] ),
    .X(net7417));
 sky130_fd_sc_hd__clkbuf_1 wire7418 (.A(net7419),
    .X(net7418));
 sky130_fd_sc_hd__clkbuf_1 wire7419 (.A(\matmul0.matmul_stage_inst.c[1] ),
    .X(net7419));
 sky130_fd_sc_hd__clkbuf_1 wire7420 (.A(\matmul0.matmul_stage_inst.b[10] ),
    .X(net7420));
 sky130_fd_sc_hd__clkbuf_1 wire7421 (.A(net7422),
    .X(net7421));
 sky130_fd_sc_hd__clkbuf_1 max_length7422 (.A(\matmul0.matmul_stage_inst.b[9] ),
    .X(net7422));
 sky130_fd_sc_hd__clkbuf_1 wire7423 (.A(\matmul0.matmul_stage_inst.b[8] ),
    .X(net7423));
 sky130_fd_sc_hd__clkbuf_1 wire7424 (.A(\matmul0.matmul_stage_inst.b[7] ),
    .X(net7424));
 sky130_fd_sc_hd__clkbuf_1 wire7425 (.A(net7426),
    .X(net7425));
 sky130_fd_sc_hd__clkbuf_1 wire7426 (.A(\matmul0.matmul_stage_inst.b[6] ),
    .X(net7426));
 sky130_fd_sc_hd__clkbuf_1 wire7427 (.A(net7428),
    .X(net7427));
 sky130_fd_sc_hd__clkbuf_1 max_length7428 (.A(\matmul0.matmul_stage_inst.b[5] ),
    .X(net7428));
 sky130_fd_sc_hd__clkbuf_1 wire7429 (.A(net7430),
    .X(net7429));
 sky130_fd_sc_hd__clkbuf_1 wire7430 (.A(net7431),
    .X(net7430));
 sky130_fd_sc_hd__clkbuf_1 max_length7431 (.A(\matmul0.matmul_stage_inst.b[4] ),
    .X(net7431));
 sky130_fd_sc_hd__clkbuf_1 wire7432 (.A(net7433),
    .X(net7432));
 sky130_fd_sc_hd__buf_1 wire7433 (.A(\matmul0.matmul_stage_inst.b[2] ),
    .X(net7433));
 sky130_fd_sc_hd__clkbuf_1 wire7434 (.A(net7435),
    .X(net7434));
 sky130_fd_sc_hd__clkbuf_1 max_length7435 (.A(\matmul0.matmul_stage_inst.b[1] ),
    .X(net7435));
 sky130_fd_sc_hd__clkbuf_1 fanout7436 (.A(net7443),
    .X(net7436));
 sky130_fd_sc_hd__buf_1 wire7437 (.A(net7438),
    .X(net7437));
 sky130_fd_sc_hd__buf_1 max_length7438 (.A(net7439),
    .X(net7438));
 sky130_fd_sc_hd__buf_1 wire7439 (.A(net7436),
    .X(net7439));
 sky130_fd_sc_hd__buf_1 fanout7440 (.A(net7443),
    .X(net7440));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7441 (.A(net7442),
    .X(net7441));
 sky130_fd_sc_hd__buf_1 wire7442 (.A(net7440),
    .X(net7442));
 sky130_fd_sc_hd__buf_1 fanout7443 (.A(net7450),
    .X(net7443));
 sky130_fd_sc_hd__clkbuf_1 wire7444 (.A(net7447),
    .X(net7444));
 sky130_fd_sc_hd__clkbuf_1 max_length7445 (.A(net7446),
    .X(net7445));
 sky130_fd_sc_hd__buf_1 wire7446 (.A(net7443),
    .X(net7446));
 sky130_fd_sc_hd__clkbuf_1 max_length7447 (.A(net7443),
    .X(net7447));
 sky130_fd_sc_hd__buf_2 fanout7448 (.A(net7449),
    .X(net7448));
 sky130_fd_sc_hd__clkbuf_1 wire7449 (.A(net7452),
    .X(net7449));
 sky130_fd_sc_hd__clkbuf_1 wire7450 (.A(net7451),
    .X(net7450));
 sky130_fd_sc_hd__clkbuf_1 max_length7451 (.A(net7452),
    .X(net7451));
 sky130_fd_sc_hd__buf_1 wire7452 (.A(\matmul0.op[1] ),
    .X(net7452));
 sky130_fd_sc_hd__buf_1 fanout7453 (.A(net7460),
    .X(net7453));
 sky130_fd_sc_hd__clkbuf_2 wire7454 (.A(net7453),
    .X(net7454));
 sky130_fd_sc_hd__buf_1 fanout7455 (.A(net7460),
    .X(net7455));
 sky130_fd_sc_hd__buf_1 wire7456 (.A(net7457),
    .X(net7456));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7457 (.A(net7455),
    .X(net7457));
 sky130_fd_sc_hd__clkbuf_1 fanout7458 (.A(\matmul0.op[0] ),
    .X(net7458));
 sky130_fd_sc_hd__buf_1 max_length7459 (.A(net7460),
    .X(net7459));
 sky130_fd_sc_hd__buf_1 wire7460 (.A(net7461),
    .X(net7460));
 sky130_fd_sc_hd__clkbuf_1 wire7461 (.A(net7458),
    .X(net7461));
 sky130_fd_sc_hd__clkbuf_1 fanout7462 (.A(net7469),
    .X(net7462));
 sky130_fd_sc_hd__buf_1 wire7463 (.A(net7465),
    .X(net7463));
 sky130_fd_sc_hd__buf_1 max_length7464 (.A(net7465),
    .X(net7464));
 sky130_fd_sc_hd__clkbuf_2 wire7465 (.A(net7462),
    .X(net7465));
 sky130_fd_sc_hd__clkbuf_2 fanout7466 (.A(\pid_q.state[5] ),
    .X(net7466));
 sky130_fd_sc_hd__buf_1 wire7467 (.A(net7466),
    .X(net7467));
 sky130_fd_sc_hd__buf_1 wire7468 (.A(net7466),
    .X(net7468));
 sky130_fd_sc_hd__clkbuf_1 wire7469 (.A(\pid_q.state[5] ),
    .X(net7469));
 sky130_fd_sc_hd__buf_1 fanout7470 (.A(\pid_q.state[4] ),
    .X(net7470));
 sky130_fd_sc_hd__clkbuf_1 max_length7471 (.A(net7472),
    .X(net7471));
 sky130_fd_sc_hd__buf_1 wire7472 (.A(net7473),
    .X(net7472));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7473 (.A(net7474),
    .X(net7473));
 sky130_fd_sc_hd__clkbuf_1 wire7474 (.A(net7470),
    .X(net7474));
 sky130_fd_sc_hd__clkbuf_1 wire7475 (.A(net7476),
    .X(net7475));
 sky130_fd_sc_hd__clkbuf_1 wire7476 (.A(net7470),
    .X(net7476));
 sky130_fd_sc_hd__buf_1 wire7477 (.A(\pid_q.state[4] ),
    .X(net7477));
 sky130_fd_sc_hd__clkbuf_1 max_length7478 (.A(\pid_q.state[4] ),
    .X(net7478));
 sky130_fd_sc_hd__buf_1 fanout7479 (.A(net7487),
    .X(net7479));
 sky130_fd_sc_hd__buf_1 wire7480 (.A(net7482),
    .X(net7480));
 sky130_fd_sc_hd__buf_1 wire7481 (.A(net7482),
    .X(net7481));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7482 (.A(net7479),
    .X(net7482));
 sky130_fd_sc_hd__buf_1 fanout7483 (.A(\pid_q.state[3] ),
    .X(net7483));
 sky130_fd_sc_hd__clkbuf_1 wire7484 (.A(net7485),
    .X(net7484));
 sky130_fd_sc_hd__buf_1 wire7485 (.A(net7486),
    .X(net7485));
 sky130_fd_sc_hd__buf_1 wire7486 (.A(net7483),
    .X(net7486));
 sky130_fd_sc_hd__clkbuf_1 wire7487 (.A(net7488),
    .X(net7487));
 sky130_fd_sc_hd__buf_1 wire7488 (.A(net7489),
    .X(net7488));
 sky130_fd_sc_hd__buf_1 max_length7489 (.A(net7483),
    .X(net7489));
 sky130_fd_sc_hd__buf_1 wire7490 (.A(net7491),
    .X(net7490));
 sky130_fd_sc_hd__clkbuf_1 wire7491 (.A(net7492),
    .X(net7491));
 sky130_fd_sc_hd__clkbuf_1 wire7492 (.A(net7493),
    .X(net7492));
 sky130_fd_sc_hd__clkbuf_1 wire7493 (.A(net7494),
    .X(net7493));
 sky130_fd_sc_hd__clkbuf_1 wire7494 (.A(net7495),
    .X(net7494));
 sky130_fd_sc_hd__clkbuf_1 wire7495 (.A(\pid_q.state[3] ),
    .X(net7495));
 sky130_fd_sc_hd__buf_1 fanout7496 (.A(net7508),
    .X(net7496));
 sky130_fd_sc_hd__clkbuf_1 max_length7497 (.A(net7498),
    .X(net7497));
 sky130_fd_sc_hd__buf_1 wire7498 (.A(net7499),
    .X(net7498));
 sky130_fd_sc_hd__buf_1 wire7499 (.A(net7500),
    .X(net7499));
 sky130_fd_sc_hd__buf_1 wire7500 (.A(net7496),
    .X(net7500));
 sky130_fd_sc_hd__buf_1 fanout7501 (.A(net7507),
    .X(net7501));
 sky130_fd_sc_hd__clkbuf_1 wire7502 (.A(net7501),
    .X(net7502));
 sky130_fd_sc_hd__clkbuf_1 wire7503 (.A(net7504),
    .X(net7503));
 sky130_fd_sc_hd__buf_1 wire7504 (.A(net7505),
    .X(net7504));
 sky130_fd_sc_hd__buf_1 wire7505 (.A(net7506),
    .X(net7505));
 sky130_fd_sc_hd__buf_1 wire7506 (.A(net7501),
    .X(net7506));
 sky130_fd_sc_hd__buf_1 fanout7507 (.A(net7516),
    .X(net7507));
 sky130_fd_sc_hd__clkbuf_1 wire7508 (.A(net7509),
    .X(net7508));
 sky130_fd_sc_hd__clkbuf_1 wire7509 (.A(net7507),
    .X(net7509));
 sky130_fd_sc_hd__clkbuf_1 max_length7510 (.A(net7511),
    .X(net7510));
 sky130_fd_sc_hd__buf_1 wire7511 (.A(net7515),
    .X(net7511));
 sky130_fd_sc_hd__buf_1 wire7512 (.A(net7513),
    .X(net7512));
 sky130_fd_sc_hd__clkbuf_1 wire7513 (.A(net7514),
    .X(net7513));
 sky130_fd_sc_hd__clkbuf_1 wire7514 (.A(net7515),
    .X(net7514));
 sky130_fd_sc_hd__buf_1 wire7515 (.A(net7507),
    .X(net7515));
 sky130_fd_sc_hd__clkbuf_1 wire7516 (.A(net7517),
    .X(net7516));
 sky130_fd_sc_hd__clkbuf_1 wire7517 (.A(net7518),
    .X(net7517));
 sky130_fd_sc_hd__clkbuf_1 wire7518 (.A(net7519),
    .X(net7518));
 sky130_fd_sc_hd__clkbuf_1 wire7519 (.A(net7520),
    .X(net7519));
 sky130_fd_sc_hd__clkbuf_1 wire7520 (.A(\pid_q.state[2] ),
    .X(net7520));
 sky130_fd_sc_hd__buf_1 fanout7521 (.A(\pid_q.state[1] ),
    .X(net7521));
 sky130_fd_sc_hd__buf_1 wire7522 (.A(net7524),
    .X(net7522));
 sky130_fd_sc_hd__buf_1 wire7523 (.A(net7524),
    .X(net7523));
 sky130_fd_sc_hd__clkbuf_2 wire7524 (.A(net7521),
    .X(net7524));
 sky130_fd_sc_hd__clkbuf_1 fanout7525 (.A(net7528),
    .X(net7525));
 sky130_fd_sc_hd__buf_1 wire7526 (.A(net7527),
    .X(net7526));
 sky130_fd_sc_hd__buf_1 wire7527 (.A(net7525),
    .X(net7527));
 sky130_fd_sc_hd__clkbuf_1 wire7528 (.A(net7529),
    .X(net7528));
 sky130_fd_sc_hd__clkbuf_1 wire7529 (.A(\pid_q.state[1] ),
    .X(net7529));
 sky130_fd_sc_hd__clkbuf_1 max_length7530 (.A(net7531),
    .X(net7530));
 sky130_fd_sc_hd__clkbuf_2 wire7531 (.A(net7532),
    .X(net7531));
 sky130_fd_sc_hd__clkbuf_1 wire7532 (.A(net7533),
    .X(net7532));
 sky130_fd_sc_hd__clkbuf_1 wire7533 (.A(net7534),
    .X(net7533));
 sky130_fd_sc_hd__clkbuf_1 wire7534 (.A(\pid_d.iterate_enable ),
    .X(net7534));
 sky130_fd_sc_hd__clkbuf_1 wire7535 (.A(net7536),
    .X(net7535));
 sky130_fd_sc_hd__clkbuf_1 wire7536 (.A(net7537),
    .X(net7536));
 sky130_fd_sc_hd__clkbuf_1 wire7537 (.A(net7538),
    .X(net7537));
 sky130_fd_sc_hd__clkbuf_1 wire7538 (.A(net7539),
    .X(net7538));
 sky130_fd_sc_hd__clkbuf_1 wire7539 (.A(net7540),
    .X(net7539));
 sky130_fd_sc_hd__clkbuf_1 wire7540 (.A(net7541),
    .X(net7540));
 sky130_fd_sc_hd__clkbuf_1 wire7541 (.A(net7542),
    .X(net7541));
 sky130_fd_sc_hd__clkbuf_1 wire7542 (.A(net7543),
    .X(net7542));
 sky130_fd_sc_hd__clkbuf_1 wire7543 (.A(net7544),
    .X(net7543));
 sky130_fd_sc_hd__clkbuf_1 wire7544 (.A(net7545),
    .X(net7544));
 sky130_fd_sc_hd__clkbuf_1 wire7545 (.A(\cordic0.in_valid ),
    .X(net7545));
 sky130_fd_sc_hd__clkbuf_1 wire7546 (.A(net7547),
    .X(net7546));
 sky130_fd_sc_hd__clkbuf_1 wire7547 (.A(\svm0.vC[11] ),
    .X(net7547));
 sky130_fd_sc_hd__clkbuf_1 wire7548 (.A(net7549),
    .X(net7548));
 sky130_fd_sc_hd__clkbuf_1 wire7549 (.A(\svm0.vC[9] ),
    .X(net7549));
 sky130_fd_sc_hd__clkbuf_1 wire7550 (.A(\matmul0.op_in[1] ),
    .X(net7550));
 sky130_fd_sc_hd__clkbuf_1 wire7551 (.A(net7552),
    .X(net7551));
 sky130_fd_sc_hd__clkbuf_1 wire7552 (.A(\matmul0.op_in[0] ),
    .X(net7552));
 sky130_fd_sc_hd__clkbuf_1 wire7553 (.A(net7554),
    .X(net7553));
 sky130_fd_sc_hd__clkbuf_1 wire7554 (.A(net7555),
    .X(net7554));
 sky130_fd_sc_hd__clkbuf_1 wire7555 (.A(\matmul0.b_in[15] ),
    .X(net7555));
 sky130_fd_sc_hd__clkbuf_1 wire7556 (.A(net7557),
    .X(net7556));
 sky130_fd_sc_hd__clkbuf_1 wire7557 (.A(net7558),
    .X(net7557));
 sky130_fd_sc_hd__clkbuf_1 wire7558 (.A(\matmul0.b_in[14] ),
    .X(net7558));
 sky130_fd_sc_hd__clkbuf_1 wire7559 (.A(net7560),
    .X(net7559));
 sky130_fd_sc_hd__clkbuf_1 wire7560 (.A(\matmul0.b_in[13] ),
    .X(net7560));
 sky130_fd_sc_hd__clkbuf_1 wire7561 (.A(\matmul0.b_in[12] ),
    .X(net7561));
 sky130_fd_sc_hd__clkbuf_1 wire7562 (.A(net7563),
    .X(net7562));
 sky130_fd_sc_hd__clkbuf_1 max_length7563 (.A(\matmul0.b_in[11] ),
    .X(net7563));
 sky130_fd_sc_hd__clkbuf_1 wire7564 (.A(net7565),
    .X(net7564));
 sky130_fd_sc_hd__clkbuf_1 wire7565 (.A(\matmul0.b_in[10] ),
    .X(net7565));
 sky130_fd_sc_hd__clkbuf_1 wire7566 (.A(\matmul0.b_in[9] ),
    .X(net7566));
 sky130_fd_sc_hd__clkbuf_1 wire7567 (.A(\matmul0.b_in[7] ),
    .X(net7567));
 sky130_fd_sc_hd__clkbuf_1 wire7568 (.A(net7569),
    .X(net7568));
 sky130_fd_sc_hd__clkbuf_1 wire7569 (.A(net7570),
    .X(net7569));
 sky130_fd_sc_hd__clkbuf_1 wire7570 (.A(\matmul0.b_in[6] ),
    .X(net7570));
 sky130_fd_sc_hd__clkbuf_1 wire7571 (.A(net7572),
    .X(net7571));
 sky130_fd_sc_hd__clkbuf_1 wire7572 (.A(\matmul0.b_in[5] ),
    .X(net7572));
 sky130_fd_sc_hd__clkbuf_1 wire7573 (.A(\matmul0.b_in[3] ),
    .X(net7573));
 sky130_fd_sc_hd__clkbuf_1 wire7574 (.A(\matmul0.b_in[1] ),
    .X(net7574));
 sky130_fd_sc_hd__clkbuf_1 wire7575 (.A(net7576),
    .X(net7575));
 sky130_fd_sc_hd__clkbuf_1 max_length7576 (.A(\matmul0.b_in[0] ),
    .X(net7576));
 sky130_fd_sc_hd__clkbuf_1 wire7577 (.A(net7578),
    .X(net7577));
 sky130_fd_sc_hd__clkbuf_1 wire7578 (.A(net7579),
    .X(net7578));
 sky130_fd_sc_hd__clkbuf_1 wire7579 (.A(net7580),
    .X(net7579));
 sky130_fd_sc_hd__buf_1 wire7580 (.A(\matmul0.a_in[15] ),
    .X(net7580));
 sky130_fd_sc_hd__clkbuf_1 wire7581 (.A(net7582),
    .X(net7581));
 sky130_fd_sc_hd__clkbuf_1 wire7582 (.A(net7583),
    .X(net7582));
 sky130_fd_sc_hd__clkbuf_1 wire7583 (.A(net7584),
    .X(net7583));
 sky130_fd_sc_hd__buf_1 wire7584 (.A(\matmul0.a_in[14] ),
    .X(net7584));
 sky130_fd_sc_hd__clkbuf_1 wire7585 (.A(net7586),
    .X(net7585));
 sky130_fd_sc_hd__clkbuf_1 wire7586 (.A(net7587),
    .X(net7586));
 sky130_fd_sc_hd__clkbuf_1 wire7587 (.A(net7588),
    .X(net7587));
 sky130_fd_sc_hd__clkbuf_1 wire7588 (.A(\matmul0.a_in[13] ),
    .X(net7588));
 sky130_fd_sc_hd__clkbuf_1 wire7589 (.A(net7590),
    .X(net7589));
 sky130_fd_sc_hd__clkbuf_1 wire7590 (.A(net7591),
    .X(net7590));
 sky130_fd_sc_hd__clkbuf_1 wire7591 (.A(\matmul0.a_in[12] ),
    .X(net7591));
 sky130_fd_sc_hd__clkbuf_1 wire7592 (.A(net7593),
    .X(net7592));
 sky130_fd_sc_hd__clkbuf_1 wire7593 (.A(net7594),
    .X(net7593));
 sky130_fd_sc_hd__clkbuf_1 wire7594 (.A(\matmul0.a_in[11] ),
    .X(net7594));
 sky130_fd_sc_hd__clkbuf_1 wire7595 (.A(net7596),
    .X(net7595));
 sky130_fd_sc_hd__clkbuf_1 wire7596 (.A(net7597),
    .X(net7596));
 sky130_fd_sc_hd__clkbuf_1 wire7597 (.A(\matmul0.a_in[10] ),
    .X(net7597));
 sky130_fd_sc_hd__clkbuf_1 wire7598 (.A(net7599),
    .X(net7598));
 sky130_fd_sc_hd__clkbuf_1 wire7599 (.A(\matmul0.a_in[9] ),
    .X(net7599));
 sky130_fd_sc_hd__clkbuf_1 wire7600 (.A(\matmul0.a_in[8] ),
    .X(net7600));
 sky130_fd_sc_hd__clkbuf_1 fanout7601 (.A(net7611),
    .X(net7601));
 sky130_fd_sc_hd__buf_1 wire7602 (.A(net7603),
    .X(net7602));
 sky130_fd_sc_hd__buf_1 wire7603 (.A(net7604),
    .X(net7603));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7604 (.A(net7601),
    .X(net7604));
 sky130_fd_sc_hd__clkbuf_1 fanout7605 (.A(net7613),
    .X(net7605));
 sky130_fd_sc_hd__buf_1 wire7606 (.A(net7607),
    .X(net7606));
 sky130_fd_sc_hd__buf_1 wire7607 (.A(net7609),
    .X(net7607));
 sky130_fd_sc_hd__clkbuf_1 max_length7608 (.A(net7609),
    .X(net7608));
 sky130_fd_sc_hd__buf_1 wire7609 (.A(net7610),
    .X(net7609));
 sky130_fd_sc_hd__buf_1 wire7610 (.A(net7605),
    .X(net7610));
 sky130_fd_sc_hd__buf_1 fanout7611 (.A(net7620),
    .X(net7611));
 sky130_fd_sc_hd__clkbuf_1 wire7612 (.A(net7613),
    .X(net7612));
 sky130_fd_sc_hd__buf_1 wire7613 (.A(net7611),
    .X(net7613));
 sky130_fd_sc_hd__clkbuf_1 fanout7614 (.A(\svm0.periodTop[15] ),
    .X(net7614));
 sky130_fd_sc_hd__clkbuf_2 wire7615 (.A(net7616),
    .X(net7615));
 sky130_fd_sc_hd__buf_1 max_length7616 (.A(net7617),
    .X(net7616));
 sky130_fd_sc_hd__buf_1 wire7617 (.A(net7618),
    .X(net7617));
 sky130_fd_sc_hd__clkbuf_1 wire7618 (.A(net7619),
    .X(net7618));
 sky130_fd_sc_hd__buf_1 wire7619 (.A(net7614),
    .X(net7619));
 sky130_fd_sc_hd__clkbuf_1 wire7620 (.A(net7621),
    .X(net7620));
 sky130_fd_sc_hd__buf_1 wire7621 (.A(net7622),
    .X(net7621));
 sky130_fd_sc_hd__clkbuf_1 wire7622 (.A(net7623),
    .X(net7622));
 sky130_fd_sc_hd__clkbuf_1 wire7623 (.A(net7624),
    .X(net7623));
 sky130_fd_sc_hd__clkbuf_1 wire7624 (.A(\svm0.periodTop[15] ),
    .X(net7624));
 sky130_fd_sc_hd__buf_1 fanout7625 (.A(net7633),
    .X(net7625));
 sky130_fd_sc_hd__buf_1 wire7626 (.A(net7627),
    .X(net7626));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7627 (.A(net7625),
    .X(net7627));
 sky130_fd_sc_hd__clkbuf_1 fanout7628 (.A(net7633),
    .X(net7628));
 sky130_fd_sc_hd__buf_1 wire7629 (.A(net7631),
    .X(net7629));
 sky130_fd_sc_hd__buf_1 wire7630 (.A(net7631),
    .X(net7630));
 sky130_fd_sc_hd__buf_1 wire7631 (.A(net7632),
    .X(net7631));
 sky130_fd_sc_hd__buf_1 wire7632 (.A(net7628),
    .X(net7632));
 sky130_fd_sc_hd__clkbuf_2 fanout7633 (.A(net7635),
    .X(net7633));
 sky130_fd_sc_hd__clkbuf_1 fanout7634 (.A(\svm0.periodTop[14] ),
    .X(net7634));
 sky130_fd_sc_hd__clkbuf_1 max_length7635 (.A(net7636),
    .X(net7635));
 sky130_fd_sc_hd__clkbuf_1 wire7636 (.A(net7637),
    .X(net7636));
 sky130_fd_sc_hd__buf_1 max_length7637 (.A(net7638),
    .X(net7637));
 sky130_fd_sc_hd__buf_1 wire7638 (.A(net7639),
    .X(net7638));
 sky130_fd_sc_hd__clkbuf_1 wire7639 (.A(net7640),
    .X(net7639));
 sky130_fd_sc_hd__buf_1 wire7640 (.A(net7634),
    .X(net7640));
 sky130_fd_sc_hd__buf_1 fanout7641 (.A(net7648),
    .X(net7641));
 sky130_fd_sc_hd__buf_1 wire7642 (.A(net7641),
    .X(net7642));
 sky130_fd_sc_hd__buf_1 wire7643 (.A(net7644),
    .X(net7643));
 sky130_fd_sc_hd__clkbuf_1 wire7644 (.A(net7645),
    .X(net7644));
 sky130_fd_sc_hd__buf_1 wire7645 (.A(net7641),
    .X(net7645));
 sky130_fd_sc_hd__buf_1 fanout7646 (.A(net7651),
    .X(net7646));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7647 (.A(net7646),
    .X(net7647));
 sky130_fd_sc_hd__buf_1 wire7648 (.A(net7646),
    .X(net7648));
 sky130_fd_sc_hd__buf_1 fanout7649 (.A(\svm0.periodTop[13] ),
    .X(net7649));
 sky130_fd_sc_hd__buf_1 wire7650 (.A(net7649),
    .X(net7650));
 sky130_fd_sc_hd__clkbuf_1 wire7651 (.A(net7652),
    .X(net7651));
 sky130_fd_sc_hd__clkbuf_1 wire7652 (.A(net7653),
    .X(net7652));
 sky130_fd_sc_hd__buf_1 max_length7653 (.A(net7654),
    .X(net7653));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7654 (.A(net7655),
    .X(net7654));
 sky130_fd_sc_hd__buf_1 wire7655 (.A(net7656),
    .X(net7655));
 sky130_fd_sc_hd__clkbuf_1 wire7656 (.A(net7649),
    .X(net7656));
 sky130_fd_sc_hd__clkbuf_1 wire7657 (.A(net7658),
    .X(net7657));
 sky130_fd_sc_hd__clkbuf_1 wire7658 (.A(net7659),
    .X(net7658));
 sky130_fd_sc_hd__clkbuf_1 wire7659 (.A(\svm0.periodTop[13] ),
    .X(net7659));
 sky130_fd_sc_hd__clkbuf_1 fanout7660 (.A(net7665),
    .X(net7660));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7661 (.A(net7663),
    .X(net7661));
 sky130_fd_sc_hd__buf_1 max_length7662 (.A(net7663),
    .X(net7662));
 sky130_fd_sc_hd__buf_1 wire7663 (.A(net7664),
    .X(net7663));
 sky130_fd_sc_hd__buf_1 wire7664 (.A(net7660),
    .X(net7664));
 sky130_fd_sc_hd__buf_1 fanout7665 (.A(net7675),
    .X(net7665));
 sky130_fd_sc_hd__buf_1 wire7666 (.A(net7667),
    .X(net7666));
 sky130_fd_sc_hd__clkbuf_1 wire7667 (.A(net7668),
    .X(net7667));
 sky130_fd_sc_hd__clkbuf_1 wire7668 (.A(net7669),
    .X(net7668));
 sky130_fd_sc_hd__buf_1 wire7669 (.A(net7665),
    .X(net7669));
 sky130_fd_sc_hd__buf_1 fanout7670 (.A(\svm0.periodTop[12] ),
    .X(net7670));
 sky130_fd_sc_hd__buf_1 wire7671 (.A(net7673),
    .X(net7671));
 sky130_fd_sc_hd__buf_1 wire7672 (.A(net7674),
    .X(net7672));
 sky130_fd_sc_hd__clkbuf_1 max_length7673 (.A(net7674),
    .X(net7673));
 sky130_fd_sc_hd__buf_1 wire7674 (.A(net7670),
    .X(net7674));
 sky130_fd_sc_hd__buf_1 wire7675 (.A(net7676),
    .X(net7675));
 sky130_fd_sc_hd__clkbuf_1 wire7676 (.A(net7677),
    .X(net7676));
 sky130_fd_sc_hd__clkbuf_1 wire7677 (.A(net7678),
    .X(net7677));
 sky130_fd_sc_hd__clkbuf_1 wire7678 (.A(\svm0.periodTop[12] ),
    .X(net7678));
 sky130_fd_sc_hd__buf_1 fanout7679 (.A(net7695),
    .X(net7679));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7680 (.A(net7681),
    .X(net7680));
 sky130_fd_sc_hd__buf_1 wire7681 (.A(net7679),
    .X(net7681));
 sky130_fd_sc_hd__buf_1 wire7682 (.A(net7683),
    .X(net7682));
 sky130_fd_sc_hd__buf_1 max_length7683 (.A(net7679),
    .X(net7683));
 sky130_fd_sc_hd__buf_1 fanout7684 (.A(net7699),
    .X(net7684));
 sky130_fd_sc_hd__clkbuf_1 wire7685 (.A(net7684),
    .X(net7685));
 sky130_fd_sc_hd__clkbuf_1 wire7686 (.A(net7687),
    .X(net7686));
 sky130_fd_sc_hd__buf_1 wire7687 (.A(net7690),
    .X(net7687));
 sky130_fd_sc_hd__clkbuf_1 max_length7688 (.A(net7689),
    .X(net7688));
 sky130_fd_sc_hd__clkbuf_1 wire7689 (.A(net7690),
    .X(net7689));
 sky130_fd_sc_hd__buf_1 wire7690 (.A(net7684),
    .X(net7690));
 sky130_fd_sc_hd__clkbuf_1 fanout7691 (.A(\svm0.periodTop[11] ),
    .X(net7691));
 sky130_fd_sc_hd__clkbuf_1 wire7692 (.A(net7693),
    .X(net7692));
 sky130_fd_sc_hd__clkbuf_1 wire7693 (.A(net7694),
    .X(net7693));
 sky130_fd_sc_hd__clkbuf_1 wire7694 (.A(net7697),
    .X(net7694));
 sky130_fd_sc_hd__clkbuf_1 max_length7695 (.A(net7696),
    .X(net7695));
 sky130_fd_sc_hd__clkbuf_1 wire7696 (.A(net7697),
    .X(net7696));
 sky130_fd_sc_hd__buf_1 wire7697 (.A(net7698),
    .X(net7697));
 sky130_fd_sc_hd__buf_1 wire7698 (.A(net7699),
    .X(net7698));
 sky130_fd_sc_hd__buf_1 wire7699 (.A(net7691),
    .X(net7699));
 sky130_fd_sc_hd__clkbuf_1 fanout7700 (.A(net7708),
    .X(net7700));
 sky130_fd_sc_hd__clkbuf_1 max_length7701 (.A(net7702),
    .X(net7701));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7702 (.A(net7703),
    .X(net7702));
 sky130_fd_sc_hd__buf_1 wire7703 (.A(net7704),
    .X(net7703));
 sky130_fd_sc_hd__buf_1 wire7704 (.A(net7700),
    .X(net7704));
 sky130_fd_sc_hd__buf_1 fanout7705 (.A(net7712),
    .X(net7705));
 sky130_fd_sc_hd__buf_1 wire7706 (.A(net7707),
    .X(net7706));
 sky130_fd_sc_hd__clkbuf_1 wire7707 (.A(net7709),
    .X(net7707));
 sky130_fd_sc_hd__buf_1 wire7708 (.A(net7709),
    .X(net7708));
 sky130_fd_sc_hd__buf_1 wire7709 (.A(net7710),
    .X(net7709));
 sky130_fd_sc_hd__buf_1 wire7710 (.A(net7705),
    .X(net7710));
 sky130_fd_sc_hd__clkbuf_1 fanout7711 (.A(\svm0.periodTop[10] ),
    .X(net7711));
 sky130_fd_sc_hd__clkbuf_1 max_length7712 (.A(net7713),
    .X(net7712));
 sky130_fd_sc_hd__buf_1 wire7713 (.A(net7714),
    .X(net7713));
 sky130_fd_sc_hd__buf_1 wire7714 (.A(net7716),
    .X(net7714));
 sky130_fd_sc_hd__buf_1 wire7715 (.A(net7716),
    .X(net7715));
 sky130_fd_sc_hd__buf_1 wire7716 (.A(net7711),
    .X(net7716));
 sky130_fd_sc_hd__clkbuf_1 fanout7717 (.A(net7729),
    .X(net7717));
 sky130_fd_sc_hd__buf_1 wire7718 (.A(net7721),
    .X(net7718));
 sky130_fd_sc_hd__buf_1 wire7719 (.A(net7720),
    .X(net7719));
 sky130_fd_sc_hd__buf_1 max_length7720 (.A(net7721),
    .X(net7720));
 sky130_fd_sc_hd__buf_1 wire7721 (.A(net7717),
    .X(net7721));
 sky130_fd_sc_hd__buf_1 fanout7722 (.A(net7730),
    .X(net7722));
 sky130_fd_sc_hd__clkbuf_1 max_length7723 (.A(net7722),
    .X(net7723));
 sky130_fd_sc_hd__buf_1 fanout7724 (.A(\svm0.periodTop[9] ),
    .X(net7724));
 sky130_fd_sc_hd__clkbuf_1 wire7725 (.A(net7726),
    .X(net7725));
 sky130_fd_sc_hd__clkbuf_1 wire7726 (.A(net7727),
    .X(net7726));
 sky130_fd_sc_hd__buf_1 wire7727 (.A(net7728),
    .X(net7727));
 sky130_fd_sc_hd__buf_1 wire7728 (.A(net7733),
    .X(net7728));
 sky130_fd_sc_hd__clkbuf_1 wire7729 (.A(net7730),
    .X(net7729));
 sky130_fd_sc_hd__buf_1 wire7730 (.A(net7731),
    .X(net7730));
 sky130_fd_sc_hd__clkbuf_1 wire7731 (.A(net7732),
    .X(net7731));
 sky130_fd_sc_hd__clkbuf_1 max_length7732 (.A(net7733),
    .X(net7732));
 sky130_fd_sc_hd__buf_1 wire7733 (.A(net7724),
    .X(net7733));
 sky130_fd_sc_hd__buf_1 fanout7734 (.A(net7754),
    .X(net7734));
 sky130_fd_sc_hd__clkbuf_1 wire7735 (.A(net7736),
    .X(net7735));
 sky130_fd_sc_hd__buf_1 wire7736 (.A(net7737),
    .X(net7736));
 sky130_fd_sc_hd__buf_1 wire7737 (.A(net7738),
    .X(net7737));
 sky130_fd_sc_hd__buf_1 wire7738 (.A(net7739),
    .X(net7738));
 sky130_fd_sc_hd__clkbuf_1 wire7739 (.A(net7740),
    .X(net7739));
 sky130_fd_sc_hd__buf_1 wire7740 (.A(net7734),
    .X(net7740));
 sky130_fd_sc_hd__buf_1 fanout7741 (.A(net7750),
    .X(net7741));
 sky130_fd_sc_hd__buf_1 max_length7742 (.A(net7743),
    .X(net7742));
 sky130_fd_sc_hd__buf_1 wire7743 (.A(net7741),
    .X(net7743));
 sky130_fd_sc_hd__buf_1 wire7744 (.A(net7741),
    .X(net7744));
 sky130_fd_sc_hd__buf_1 fanout7745 (.A(net7752),
    .X(net7745));
 sky130_fd_sc_hd__buf_1 wire7746 (.A(net7747),
    .X(net7746));
 sky130_fd_sc_hd__buf_1 wire7747 (.A(net7745),
    .X(net7747));
 sky130_fd_sc_hd__clkbuf_1 wire7748 (.A(net7749),
    .X(net7748));
 sky130_fd_sc_hd__clkbuf_1 wire7749 (.A(net7753),
    .X(net7749));
 sky130_fd_sc_hd__clkbuf_1 wire7750 (.A(net7751),
    .X(net7750));
 sky130_fd_sc_hd__clkbuf_1 wire7751 (.A(net7752),
    .X(net7751));
 sky130_fd_sc_hd__buf_1 wire7752 (.A(net7753),
    .X(net7752));
 sky130_fd_sc_hd__buf_1 wire7753 (.A(net7754),
    .X(net7753));
 sky130_fd_sc_hd__buf_1 wire7754 (.A(\svm0.periodTop[8] ),
    .X(net7754));
 sky130_fd_sc_hd__clkbuf_1 fanout7755 (.A(net7774),
    .X(net7755));
 sky130_fd_sc_hd__clkbuf_1 wire7756 (.A(net7757),
    .X(net7756));
 sky130_fd_sc_hd__buf_1 wire7757 (.A(net7758),
    .X(net7757));
 sky130_fd_sc_hd__buf_1 wire7758 (.A(net7759),
    .X(net7758));
 sky130_fd_sc_hd__buf_1 wire7759 (.A(net7760),
    .X(net7759));
 sky130_fd_sc_hd__buf_1 wire7760 (.A(net7761),
    .X(net7760));
 sky130_fd_sc_hd__clkbuf_1 wire7761 (.A(net7762),
    .X(net7761));
 sky130_fd_sc_hd__clkbuf_1 max_length7762 (.A(net7755),
    .X(net7762));
 sky130_fd_sc_hd__clkbuf_1 fanout7763 (.A(net7772),
    .X(net7763));
 sky130_fd_sc_hd__clkbuf_1 max_length7764 (.A(net7765),
    .X(net7764));
 sky130_fd_sc_hd__buf_1 wire7765 (.A(net7766),
    .X(net7765));
 sky130_fd_sc_hd__buf_1 wire7766 (.A(net7767),
    .X(net7766));
 sky130_fd_sc_hd__clkbuf_1 wire7767 (.A(net7763),
    .X(net7767));
 sky130_fd_sc_hd__buf_1 max_length7768 (.A(net7763),
    .X(net7768));
 sky130_fd_sc_hd__clkbuf_2 fanout7769 (.A(net7774),
    .X(net7769));
 sky130_fd_sc_hd__buf_1 wire7770 (.A(net7769),
    .X(net7770));
 sky130_fd_sc_hd__buf_1 fanout7771 (.A(\svm0.periodTop[7] ),
    .X(net7771));
 sky130_fd_sc_hd__clkbuf_1 wire7772 (.A(net7773),
    .X(net7772));
 sky130_fd_sc_hd__clkbuf_1 wire7773 (.A(net7774),
    .X(net7773));
 sky130_fd_sc_hd__clkbuf_2 wire7774 (.A(net7775),
    .X(net7774));
 sky130_fd_sc_hd__clkbuf_1 wire7775 (.A(net7776),
    .X(net7775));
 sky130_fd_sc_hd__clkbuf_1 max_length7776 (.A(net7771),
    .X(net7776));
 sky130_fd_sc_hd__buf_1 fanout7777 (.A(net7797),
    .X(net7777));
 sky130_fd_sc_hd__buf_1 wire7778 (.A(net7779),
    .X(net7778));
 sky130_fd_sc_hd__buf_1 wire7779 (.A(net7783),
    .X(net7779));
 sky130_fd_sc_hd__clkbuf_1 wire7780 (.A(net7781),
    .X(net7780));
 sky130_fd_sc_hd__clkbuf_1 wire7781 (.A(net7782),
    .X(net7781));
 sky130_fd_sc_hd__clkbuf_1 max_length7782 (.A(net7783),
    .X(net7782));
 sky130_fd_sc_hd__buf_1 wire7783 (.A(net7785),
    .X(net7783));
 sky130_fd_sc_hd__buf_1 wire7784 (.A(net7777),
    .X(net7784));
 sky130_fd_sc_hd__buf_1 max_length7785 (.A(net7777),
    .X(net7785));
 sky130_fd_sc_hd__clkbuf_1 fanout7786 (.A(net7793),
    .X(net7786));
 sky130_fd_sc_hd__buf_1 wire7787 (.A(net7788),
    .X(net7787));
 sky130_fd_sc_hd__buf_1 wire7788 (.A(net7789),
    .X(net7788));
 sky130_fd_sc_hd__buf_1 wire7789 (.A(net7790),
    .X(net7789));
 sky130_fd_sc_hd__buf_1 wire7790 (.A(net7786),
    .X(net7790));
 sky130_fd_sc_hd__buf_1 fanout7791 (.A(\svm0.periodTop[6] ),
    .X(net7791));
 sky130_fd_sc_hd__buf_1 wire7792 (.A(net7793),
    .X(net7792));
 sky130_fd_sc_hd__buf_1 wire7793 (.A(net7794),
    .X(net7793));
 sky130_fd_sc_hd__clkbuf_1 wire7794 (.A(net7795),
    .X(net7794));
 sky130_fd_sc_hd__clkbuf_1 wire7795 (.A(net7796),
    .X(net7795));
 sky130_fd_sc_hd__clkbuf_1 wire7796 (.A(net7799),
    .X(net7796));
 sky130_fd_sc_hd__clkbuf_1 wire7797 (.A(net7798),
    .X(net7797));
 sky130_fd_sc_hd__clkbuf_1 wire7798 (.A(net7791),
    .X(net7798));
 sky130_fd_sc_hd__clkbuf_1 max_length7799 (.A(net7791),
    .X(net7799));
 sky130_fd_sc_hd__buf_1 fanout7800 (.A(net7813),
    .X(net7800));
 sky130_fd_sc_hd__clkbuf_1 max_length7801 (.A(net7802),
    .X(net7801));
 sky130_fd_sc_hd__buf_1 wire7802 (.A(net7803),
    .X(net7802));
 sky130_fd_sc_hd__buf_1 max_length7803 (.A(net7804),
    .X(net7803));
 sky130_fd_sc_hd__clkbuf_2 wire7804 (.A(net7800),
    .X(net7804));
 sky130_fd_sc_hd__clkbuf_1 fanout7805 (.A(net7814),
    .X(net7805));
 sky130_fd_sc_hd__buf_1 wire7806 (.A(net7807),
    .X(net7806));
 sky130_fd_sc_hd__buf_1 wire7807 (.A(net7811),
    .X(net7807));
 sky130_fd_sc_hd__clkbuf_1 wire7808 (.A(net7809),
    .X(net7808));
 sky130_fd_sc_hd__clkbuf_1 wire7809 (.A(net7810),
    .X(net7809));
 sky130_fd_sc_hd__buf_1 wire7810 (.A(net7811),
    .X(net7810));
 sky130_fd_sc_hd__buf_1 wire7811 (.A(net7805),
    .X(net7811));
 sky130_fd_sc_hd__buf_1 fanout7812 (.A(\svm0.periodTop[5] ),
    .X(net7812));
 sky130_fd_sc_hd__buf_1 wire7813 (.A(net7819),
    .X(net7813));
 sky130_fd_sc_hd__buf_1 wire7814 (.A(net7815),
    .X(net7814));
 sky130_fd_sc_hd__buf_1 wire7815 (.A(net7816),
    .X(net7815));
 sky130_fd_sc_hd__clkbuf_1 wire7816 (.A(net7817),
    .X(net7816));
 sky130_fd_sc_hd__clkbuf_1 wire7817 (.A(net7818),
    .X(net7817));
 sky130_fd_sc_hd__clkbuf_1 wire7818 (.A(net7812),
    .X(net7818));
 sky130_fd_sc_hd__buf_1 max_length7819 (.A(net7812),
    .X(net7819));
 sky130_fd_sc_hd__clkbuf_1 fanout7820 (.A(net7843),
    .X(net7820));
 sky130_fd_sc_hd__buf_1 wire7821 (.A(net7822),
    .X(net7821));
 sky130_fd_sc_hd__buf_1 wire7822 (.A(net7823),
    .X(net7822));
 sky130_fd_sc_hd__buf_1 wire7823 (.A(net7824),
    .X(net7823));
 sky130_fd_sc_hd__buf_1 wire7824 (.A(net7825),
    .X(net7824));
 sky130_fd_sc_hd__buf_1 wire7825 (.A(net7826),
    .X(net7825));
 sky130_fd_sc_hd__buf_1 wire7826 (.A(net7820),
    .X(net7826));
 sky130_fd_sc_hd__buf_1 fanout7827 (.A(net7837),
    .X(net7827));
 sky130_fd_sc_hd__buf_1 wire7828 (.A(net7829),
    .X(net7828));
 sky130_fd_sc_hd__clkbuf_1 wire7829 (.A(net7830),
    .X(net7829));
 sky130_fd_sc_hd__clkbuf_1 wire7830 (.A(net7833),
    .X(net7830));
 sky130_fd_sc_hd__buf_1 max_length7831 (.A(net7832),
    .X(net7831));
 sky130_fd_sc_hd__buf_1 wire7832 (.A(net7833),
    .X(net7832));
 sky130_fd_sc_hd__buf_1 wire7833 (.A(net7834),
    .X(net7833));
 sky130_fd_sc_hd__buf_1 wire7834 (.A(net7827),
    .X(net7834));
 sky130_fd_sc_hd__buf_1 fanout7835 (.A(\svm0.periodTop[4] ),
    .X(net7835));
 sky130_fd_sc_hd__buf_1 wire7836 (.A(net7843),
    .X(net7836));
 sky130_fd_sc_hd__clkbuf_1 wire7837 (.A(net7840),
    .X(net7837));
 sky130_fd_sc_hd__clkbuf_1 wire7838 (.A(net7839),
    .X(net7838));
 sky130_fd_sc_hd__clkbuf_1 max_length7839 (.A(net7840),
    .X(net7839));
 sky130_fd_sc_hd__buf_1 wire7840 (.A(net7841),
    .X(net7840));
 sky130_fd_sc_hd__clkbuf_1 wire7841 (.A(net7842),
    .X(net7841));
 sky130_fd_sc_hd__clkbuf_1 wire7842 (.A(net7835),
    .X(net7842));
 sky130_fd_sc_hd__clkbuf_1 max_length7843 (.A(net7835),
    .X(net7843));
 sky130_fd_sc_hd__clkbuf_1 fanout7844 (.A(net7857),
    .X(net7844));
 sky130_fd_sc_hd__clkbuf_1 wire7845 (.A(net7846),
    .X(net7845));
 sky130_fd_sc_hd__clkbuf_1 wire7846 (.A(net7848),
    .X(net7846));
 sky130_fd_sc_hd__buf_1 wire7847 (.A(net7848),
    .X(net7847));
 sky130_fd_sc_hd__buf_1 wire7848 (.A(net7849),
    .X(net7848));
 sky130_fd_sc_hd__buf_1 wire7849 (.A(net7850),
    .X(net7849));
 sky130_fd_sc_hd__buf_1 wire7850 (.A(net7844),
    .X(net7850));
 sky130_fd_sc_hd__clkbuf_1 fanout7851 (.A(net7856),
    .X(net7851));
 sky130_fd_sc_hd__clkbuf_1 wire7852 (.A(net7853),
    .X(net7852));
 sky130_fd_sc_hd__buf_1 wire7853 (.A(net7854),
    .X(net7853));
 sky130_fd_sc_hd__buf_1 wire7854 (.A(net7855),
    .X(net7854));
 sky130_fd_sc_hd__buf_1 wire7855 (.A(net7851),
    .X(net7855));
 sky130_fd_sc_hd__buf_1 fanout7856 (.A(\svm0.periodTop[3] ),
    .X(net7856));
 sky130_fd_sc_hd__clkbuf_1 wire7857 (.A(net7858),
    .X(net7857));
 sky130_fd_sc_hd__clkbuf_1 wire7858 (.A(net7859),
    .X(net7858));
 sky130_fd_sc_hd__clkbuf_1 wire7859 (.A(net7856),
    .X(net7859));
 sky130_fd_sc_hd__clkbuf_1 wire7860 (.A(net7861),
    .X(net7860));
 sky130_fd_sc_hd__clkbuf_1 wire7861 (.A(net7868),
    .X(net7861));
 sky130_fd_sc_hd__clkbuf_1 wire7862 (.A(net7863),
    .X(net7862));
 sky130_fd_sc_hd__clkbuf_1 wire7863 (.A(net7864),
    .X(net7863));
 sky130_fd_sc_hd__clkbuf_1 wire7864 (.A(net7865),
    .X(net7864));
 sky130_fd_sc_hd__buf_1 max_length7865 (.A(net7866),
    .X(net7865));
 sky130_fd_sc_hd__buf_1 wire7866 (.A(net7867),
    .X(net7866));
 sky130_fd_sc_hd__clkbuf_1 wire7867 (.A(net7868),
    .X(net7867));
 sky130_fd_sc_hd__buf_1 wire7868 (.A(net7856),
    .X(net7868));
 sky130_fd_sc_hd__clkbuf_1 wire7869 (.A(net7870),
    .X(net7869));
 sky130_fd_sc_hd__clkbuf_1 wire7870 (.A(net7871),
    .X(net7870));
 sky130_fd_sc_hd__clkbuf_1 wire7871 (.A(net7872),
    .X(net7871));
 sky130_fd_sc_hd__clkbuf_1 wire7872 (.A(\svm0.periodTop[3] ),
    .X(net7872));
 sky130_fd_sc_hd__clkbuf_1 fanout7873 (.A(net7885),
    .X(net7873));
 sky130_fd_sc_hd__buf_1 max_length7874 (.A(net7875),
    .X(net7874));
 sky130_fd_sc_hd__buf_1 wire7875 (.A(net7876),
    .X(net7875));
 sky130_fd_sc_hd__buf_1 wire7876 (.A(net7877),
    .X(net7876));
 sky130_fd_sc_hd__buf_1 wire7877 (.A(net7873),
    .X(net7877));
 sky130_fd_sc_hd__buf_1 fanout7878 (.A(net7884),
    .X(net7878));
 sky130_fd_sc_hd__clkbuf_1 wire7879 (.A(net7878),
    .X(net7879));
 sky130_fd_sc_hd__buf_1 fanout7880 (.A(net7899),
    .X(net7880));
 sky130_fd_sc_hd__buf_1 wire7881 (.A(net7882),
    .X(net7881));
 sky130_fd_sc_hd__buf_1 wire7882 (.A(net7883),
    .X(net7882));
 sky130_fd_sc_hd__buf_1 wire7883 (.A(net7880),
    .X(net7883));
 sky130_fd_sc_hd__clkbuf_1 max_length7884 (.A(net7885),
    .X(net7884));
 sky130_fd_sc_hd__buf_1 wire7885 (.A(net7886),
    .X(net7885));
 sky130_fd_sc_hd__clkbuf_1 wire7886 (.A(net7887),
    .X(net7886));
 sky130_fd_sc_hd__clkbuf_1 wire7887 (.A(net7880),
    .X(net7887));
 sky130_fd_sc_hd__buf_1 fanout7888 (.A(\svm0.periodTop[2] ),
    .X(net7888));
 sky130_fd_sc_hd__buf_1 wire7889 (.A(net7899),
    .X(net7889));
 sky130_fd_sc_hd__buf_1 wire7890 (.A(net7891),
    .X(net7890));
 sky130_fd_sc_hd__clkbuf_1 wire7891 (.A(net7892),
    .X(net7891));
 sky130_fd_sc_hd__clkbuf_1 wire7892 (.A(net7893),
    .X(net7892));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7893 (.A(net7894),
    .X(net7893));
 sky130_fd_sc_hd__clkbuf_1 wire7894 (.A(net7898),
    .X(net7894));
 sky130_fd_sc_hd__clkbuf_1 wire7895 (.A(net7896),
    .X(net7895));
 sky130_fd_sc_hd__clkbuf_1 wire7896 (.A(net7897),
    .X(net7896));
 sky130_fd_sc_hd__clkbuf_1 max_length7897 (.A(net7898),
    .X(net7897));
 sky130_fd_sc_hd__buf_1 wire7898 (.A(net7888),
    .X(net7898));
 sky130_fd_sc_hd__buf_1 max_length7899 (.A(net7888),
    .X(net7899));
 sky130_fd_sc_hd__clkbuf_1 wire7900 (.A(net7901),
    .X(net7900));
 sky130_fd_sc_hd__buf_1 wire7901 (.A(net7902),
    .X(net7901));
 sky130_fd_sc_hd__clkbuf_1 wire7902 (.A(net7903),
    .X(net7902));
 sky130_fd_sc_hd__clkbuf_1 wire7903 (.A(net7904),
    .X(net7903));
 sky130_fd_sc_hd__clkbuf_1 wire7904 (.A(\svm0.periodTop[2] ),
    .X(net7904));
 sky130_fd_sc_hd__buf_1 fanout7905 (.A(net7925),
    .X(net7905));
 sky130_fd_sc_hd__buf_1 wire7906 (.A(net7907),
    .X(net7906));
 sky130_fd_sc_hd__buf_1 wire7907 (.A(net7908),
    .X(net7907));
 sky130_fd_sc_hd__buf_1 wire7908 (.A(net7909),
    .X(net7908));
 sky130_fd_sc_hd__buf_1 wire7909 (.A(net7910),
    .X(net7909));
 sky130_fd_sc_hd__clkbuf_1 wire7910 (.A(net7905),
    .X(net7910));
 sky130_fd_sc_hd__clkbuf_1 wire7911 (.A(net7912),
    .X(net7911));
 sky130_fd_sc_hd__clkbuf_1 wire7912 (.A(net7913),
    .X(net7912));
 sky130_fd_sc_hd__clkbuf_1 wire7913 (.A(net7905),
    .X(net7913));
 sky130_fd_sc_hd__buf_1 fanout7914 (.A(net7918),
    .X(net7914));
 sky130_fd_sc_hd__clkbuf_1 wire7915 (.A(net7916),
    .X(net7915));
 sky130_fd_sc_hd__buf_1 max_length7916 (.A(net7917),
    .X(net7916));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7917 (.A(net7914),
    .X(net7917));
 sky130_fd_sc_hd__buf_1 fanout7918 (.A(net7929),
    .X(net7918));
 sky130_fd_sc_hd__buf_1 wire7919 (.A(net7920),
    .X(net7919));
 sky130_fd_sc_hd__clkbuf_1 wire7920 (.A(net7921),
    .X(net7920));
 sky130_fd_sc_hd__buf_1 wire7921 (.A(net7922),
    .X(net7921));
 sky130_fd_sc_hd__clkbuf_1 wire7922 (.A(net7924),
    .X(net7922));
 sky130_fd_sc_hd__buf_1 wire7923 (.A(net7925),
    .X(net7923));
 sky130_fd_sc_hd__clkbuf_1 max_length7924 (.A(net7925),
    .X(net7924));
 sky130_fd_sc_hd__buf_1 wire7925 (.A(net7918),
    .X(net7925));
 sky130_fd_sc_hd__clkbuf_1 wire7926 (.A(net7927),
    .X(net7926));
 sky130_fd_sc_hd__clkbuf_1 wire7927 (.A(net7928),
    .X(net7927));
 sky130_fd_sc_hd__clkbuf_1 wire7928 (.A(net7929),
    .X(net7928));
 sky130_fd_sc_hd__buf_1 wire7929 (.A(\svm0.periodTop[1] ),
    .X(net7929));
 sky130_fd_sc_hd__clkbuf_1 fanout7930 (.A(net7936),
    .X(net7930));
 sky130_fd_sc_hd__buf_1 wire7931 (.A(net7932),
    .X(net7931));
 sky130_fd_sc_hd__buf_1 wire7932 (.A(net7933),
    .X(net7932));
 sky130_fd_sc_hd__clkbuf_2 wire7933 (.A(net7930),
    .X(net7933));
 sky130_fd_sc_hd__clkbuf_1 fanout7934 (.A(net7942),
    .X(net7934));
 sky130_fd_sc_hd__clkbuf_1 max_length7935 (.A(net7936),
    .X(net7935));
 sky130_fd_sc_hd__buf_1 wire7936 (.A(net7937),
    .X(net7936));
 sky130_fd_sc_hd__clkbuf_1 wire7937 (.A(net7938),
    .X(net7937));
 sky130_fd_sc_hd__clkbuf_1 wire7938 (.A(net7941),
    .X(net7938));
 sky130_fd_sc_hd__clkbuf_1 wire7939 (.A(net7940),
    .X(net7939));
 sky130_fd_sc_hd__buf_1 wire7940 (.A(net7941),
    .X(net7940));
 sky130_fd_sc_hd__buf_1 wire7941 (.A(net7934),
    .X(net7941));
 sky130_fd_sc_hd__clkbuf_1 fanout7942 (.A(\svm0.periodTop[0] ),
    .X(net7942));
 sky130_fd_sc_hd__buf_1 wire7943 (.A(net7944),
    .X(net7943));
 sky130_fd_sc_hd__clkbuf_1 wire7944 (.A(net7945),
    .X(net7944));
 sky130_fd_sc_hd__clkbuf_1 wire7945 (.A(net7946),
    .X(net7945));
 sky130_fd_sc_hd__buf_1 wire7946 (.A(net7947),
    .X(net7946));
 sky130_fd_sc_hd__buf_1 wire7947 (.A(net7948),
    .X(net7947));
 sky130_fd_sc_hd__buf_1 wire7948 (.A(net7942),
    .X(net7948));
 sky130_fd_sc_hd__buf_1 wire7949 (.A(net7950),
    .X(net7949));
 sky130_fd_sc_hd__clkbuf_1 wire7950 (.A(net7951),
    .X(net7950));
 sky130_fd_sc_hd__clkbuf_1 wire7951 (.A(net7952),
    .X(net7951));
 sky130_fd_sc_hd__clkbuf_1 wire7952 (.A(net7953),
    .X(net7952));
 sky130_fd_sc_hd__clkbuf_1 wire7953 (.A(net7954),
    .X(net7953));
 sky130_fd_sc_hd__buf_1 wire7954 (.A(\pid_q.target[15] ),
    .X(net7954));
 sky130_fd_sc_hd__clkbuf_2 wire7955 (.A(net7956),
    .X(net7955));
 sky130_fd_sc_hd__clkbuf_1 wire7956 (.A(net7957),
    .X(net7956));
 sky130_fd_sc_hd__clkbuf_1 wire7957 (.A(net7958),
    .X(net7957));
 sky130_fd_sc_hd__clkbuf_1 wire7958 (.A(net7959),
    .X(net7958));
 sky130_fd_sc_hd__clkbuf_1 wire7959 (.A(net7960),
    .X(net7959));
 sky130_fd_sc_hd__clkbuf_1 wire7960 (.A(\pid_q.target[14] ),
    .X(net7960));
 sky130_fd_sc_hd__clkbuf_2 wire7961 (.A(net7962),
    .X(net7961));
 sky130_fd_sc_hd__clkbuf_1 wire7962 (.A(net7963),
    .X(net7962));
 sky130_fd_sc_hd__clkbuf_1 wire7963 (.A(net7964),
    .X(net7963));
 sky130_fd_sc_hd__clkbuf_1 wire7964 (.A(net7965),
    .X(net7964));
 sky130_fd_sc_hd__clkbuf_1 wire7965 (.A(net7966),
    .X(net7965));
 sky130_fd_sc_hd__clkbuf_1 wire7966 (.A(\pid_q.target[13] ),
    .X(net7966));
 sky130_fd_sc_hd__buf_1 wire7967 (.A(net7968),
    .X(net7967));
 sky130_fd_sc_hd__clkbuf_1 wire7968 (.A(net7969),
    .X(net7968));
 sky130_fd_sc_hd__clkbuf_1 wire7969 (.A(net7970),
    .X(net7969));
 sky130_fd_sc_hd__clkbuf_1 wire7970 (.A(net7971),
    .X(net7970));
 sky130_fd_sc_hd__clkbuf_1 wire7971 (.A(net7972),
    .X(net7971));
 sky130_fd_sc_hd__clkbuf_1 wire7972 (.A(net7973),
    .X(net7972));
 sky130_fd_sc_hd__buf_1 wire7973 (.A(\pid_q.target[12] ),
    .X(net7973));
 sky130_fd_sc_hd__buf_1 wire7974 (.A(net7975),
    .X(net7974));
 sky130_fd_sc_hd__clkbuf_1 wire7975 (.A(net7976),
    .X(net7975));
 sky130_fd_sc_hd__clkbuf_1 wire7976 (.A(net7977),
    .X(net7976));
 sky130_fd_sc_hd__clkbuf_1 wire7977 (.A(net7978),
    .X(net7977));
 sky130_fd_sc_hd__clkbuf_1 wire7978 (.A(net7979),
    .X(net7978));
 sky130_fd_sc_hd__clkbuf_1 wire7979 (.A(\pid_q.target[11] ),
    .X(net7979));
 sky130_fd_sc_hd__clkbuf_2 wire7980 (.A(net7981),
    .X(net7980));
 sky130_fd_sc_hd__clkbuf_1 wire7981 (.A(net7982),
    .X(net7981));
 sky130_fd_sc_hd__clkbuf_1 wire7982 (.A(net7983),
    .X(net7982));
 sky130_fd_sc_hd__clkbuf_1 wire7983 (.A(net7984),
    .X(net7983));
 sky130_fd_sc_hd__clkbuf_1 wire7984 (.A(\pid_q.target[10] ),
    .X(net7984));
 sky130_fd_sc_hd__clkbuf_2 wire7985 (.A(net7986),
    .X(net7985));
 sky130_fd_sc_hd__clkbuf_1 wire7986 (.A(net7987),
    .X(net7986));
 sky130_fd_sc_hd__clkbuf_1 wire7987 (.A(net7988),
    .X(net7987));
 sky130_fd_sc_hd__clkbuf_1 wire7988 (.A(net7989),
    .X(net7988));
 sky130_fd_sc_hd__clkbuf_1 wire7989 (.A(\pid_q.target[9] ),
    .X(net7989));
 sky130_fd_sc_hd__clkbuf_2 wire7990 (.A(net7991),
    .X(net7990));
 sky130_fd_sc_hd__clkbuf_1 wire7991 (.A(net7992),
    .X(net7991));
 sky130_fd_sc_hd__clkbuf_1 wire7992 (.A(net7993),
    .X(net7992));
 sky130_fd_sc_hd__clkbuf_1 wire7993 (.A(net7994),
    .X(net7993));
 sky130_fd_sc_hd__clkbuf_1 wire7994 (.A(net7995),
    .X(net7994));
 sky130_fd_sc_hd__clkbuf_1 max_length7995 (.A(\pid_q.target[8] ),
    .X(net7995));
 sky130_fd_sc_hd__clkbuf_2 wire7996 (.A(net7997),
    .X(net7996));
 sky130_fd_sc_hd__clkbuf_1 wire7997 (.A(net7998),
    .X(net7997));
 sky130_fd_sc_hd__clkbuf_1 wire7998 (.A(net7999),
    .X(net7998));
 sky130_fd_sc_hd__clkbuf_1 wire7999 (.A(net8000),
    .X(net7999));
 sky130_fd_sc_hd__clkbuf_1 wire8000 (.A(net8001),
    .X(net8000));
 sky130_fd_sc_hd__clkbuf_1 max_length8001 (.A(\pid_q.target[7] ),
    .X(net8001));
 sky130_fd_sc_hd__clkbuf_2 wire8002 (.A(net8003),
    .X(net8002));
 sky130_fd_sc_hd__clkbuf_1 wire8003 (.A(net8004),
    .X(net8003));
 sky130_fd_sc_hd__clkbuf_1 wire8004 (.A(net8005),
    .X(net8004));
 sky130_fd_sc_hd__clkbuf_1 wire8005 (.A(net8006),
    .X(net8005));
 sky130_fd_sc_hd__clkbuf_1 wire8006 (.A(\pid_q.target[6] ),
    .X(net8006));
 sky130_fd_sc_hd__buf_1 wire8007 (.A(net8008),
    .X(net8007));
 sky130_fd_sc_hd__clkbuf_1 wire8008 (.A(net8009),
    .X(net8008));
 sky130_fd_sc_hd__clkbuf_1 wire8009 (.A(net8010),
    .X(net8009));
 sky130_fd_sc_hd__clkbuf_1 wire8010 (.A(net8011),
    .X(net8010));
 sky130_fd_sc_hd__clkbuf_1 max_length8011 (.A(\pid_q.target[5] ),
    .X(net8011));
 sky130_fd_sc_hd__clkbuf_2 wire8012 (.A(net8013),
    .X(net8012));
 sky130_fd_sc_hd__clkbuf_1 wire8013 (.A(net8014),
    .X(net8013));
 sky130_fd_sc_hd__clkbuf_1 wire8014 (.A(net8015),
    .X(net8014));
 sky130_fd_sc_hd__clkbuf_1 wire8015 (.A(net8016),
    .X(net8015));
 sky130_fd_sc_hd__clkbuf_1 max_length8016 (.A(\pid_q.target[4] ),
    .X(net8016));
 sky130_fd_sc_hd__clkbuf_2 wire8017 (.A(net8018),
    .X(net8017));
 sky130_fd_sc_hd__clkbuf_1 wire8018 (.A(net8019),
    .X(net8018));
 sky130_fd_sc_hd__clkbuf_1 wire8019 (.A(net8020),
    .X(net8019));
 sky130_fd_sc_hd__clkbuf_1 wire8020 (.A(net8021),
    .X(net8020));
 sky130_fd_sc_hd__clkbuf_1 wire8021 (.A(\pid_q.target[3] ),
    .X(net8021));
 sky130_fd_sc_hd__buf_1 wire8022 (.A(net8023),
    .X(net8022));
 sky130_fd_sc_hd__buf_1 wire8023 (.A(net8024),
    .X(net8023));
 sky130_fd_sc_hd__clkbuf_1 wire8024 (.A(net8025),
    .X(net8024));
 sky130_fd_sc_hd__clkbuf_1 wire8025 (.A(net8026),
    .X(net8025));
 sky130_fd_sc_hd__clkbuf_1 wire8026 (.A(net8027),
    .X(net8026));
 sky130_fd_sc_hd__clkbuf_1 max_length8027 (.A(\pid_q.target[2] ),
    .X(net8027));
 sky130_fd_sc_hd__clkbuf_2 wire8028 (.A(net8029),
    .X(net8028));
 sky130_fd_sc_hd__clkbuf_1 wire8029 (.A(net8030),
    .X(net8029));
 sky130_fd_sc_hd__clkbuf_1 wire8030 (.A(net8031),
    .X(net8030));
 sky130_fd_sc_hd__clkbuf_1 wire8031 (.A(net8032),
    .X(net8031));
 sky130_fd_sc_hd__clkbuf_1 wire8032 (.A(net8033),
    .X(net8032));
 sky130_fd_sc_hd__clkbuf_1 wire8033 (.A(\pid_q.target[1] ),
    .X(net8033));
 sky130_fd_sc_hd__buf_1 wire8034 (.A(net8035),
    .X(net8034));
 sky130_fd_sc_hd__clkbuf_1 wire8035 (.A(net8036),
    .X(net8035));
 sky130_fd_sc_hd__clkbuf_1 wire8036 (.A(net8037),
    .X(net8036));
 sky130_fd_sc_hd__clkbuf_1 wire8037 (.A(net8038),
    .X(net8037));
 sky130_fd_sc_hd__clkbuf_1 wire8038 (.A(net8039),
    .X(net8038));
 sky130_fd_sc_hd__clkbuf_1 wire8039 (.A(net8040),
    .X(net8039));
 sky130_fd_sc_hd__clkbuf_1 max_length8040 (.A(\pid_q.target[0] ),
    .X(net8040));
 sky130_fd_sc_hd__clkbuf_1 fanout8041 (.A(net8046),
    .X(net8041));
 sky130_fd_sc_hd__clkbuf_1 wire8042 (.A(net8045),
    .X(net8042));
 sky130_fd_sc_hd__buf_1 wire8043 (.A(net8044),
    .X(net8043));
 sky130_fd_sc_hd__clkbuf_2 wire8044 (.A(net8045),
    .X(net8044));
 sky130_fd_sc_hd__buf_1 wire8045 (.A(net8041),
    .X(net8045));
 sky130_fd_sc_hd__clkbuf_1 fanout8046 (.A(net8065),
    .X(net8046));
 sky130_fd_sc_hd__clkbuf_1 max_length8047 (.A(net8048),
    .X(net8047));
 sky130_fd_sc_hd__buf_1 wire8048 (.A(net8049),
    .X(net8048));
 sky130_fd_sc_hd__buf_1 wire8049 (.A(net8050),
    .X(net8049));
 sky130_fd_sc_hd__buf_1 wire8050 (.A(net8051),
    .X(net8050));
 sky130_fd_sc_hd__clkbuf_1 wire8051 (.A(net8052),
    .X(net8051));
 sky130_fd_sc_hd__buf_1 wire8052 (.A(net8053),
    .X(net8052));
 sky130_fd_sc_hd__buf_1 wire8053 (.A(net8046),
    .X(net8053));
 sky130_fd_sc_hd__buf_1 fanout8054 (.A(net8064),
    .X(net8054));
 sky130_fd_sc_hd__buf_1 wire8055 (.A(net8056),
    .X(net8055));
 sky130_fd_sc_hd__buf_1 wire8056 (.A(net8057),
    .X(net8056));
 sky130_fd_sc_hd__clkbuf_2 wire8057 (.A(net8054),
    .X(net8057));
 sky130_fd_sc_hd__buf_1 fanout8058 (.A(net8074),
    .X(net8058));
 sky130_fd_sc_hd__clkbuf_1 wire8059 (.A(net8061),
    .X(net8059));
 sky130_fd_sc_hd__buf_1 wire8060 (.A(net8061),
    .X(net8060));
 sky130_fd_sc_hd__buf_1 wire8061 (.A(net8058),
    .X(net8061));
 sky130_fd_sc_hd__buf_1 wire8062 (.A(net8063),
    .X(net8062));
 sky130_fd_sc_hd__clkbuf_1 wire8063 (.A(net8058),
    .X(net8063));
 sky130_fd_sc_hd__buf_1 fanout8064 (.A(\cordic0.state[0] ),
    .X(net8064));
 sky130_fd_sc_hd__clkbuf_1 wire8065 (.A(net8066),
    .X(net8065));
 sky130_fd_sc_hd__clkbuf_1 wire8066 (.A(net8067),
    .X(net8066));
 sky130_fd_sc_hd__clkbuf_1 wire8067 (.A(net8068),
    .X(net8067));
 sky130_fd_sc_hd__clkbuf_1 wire8068 (.A(net8064),
    .X(net8068));
 sky130_fd_sc_hd__buf_1 wire8069 (.A(net8070),
    .X(net8069));
 sky130_fd_sc_hd__clkbuf_1 wire8070 (.A(net8071),
    .X(net8070));
 sky130_fd_sc_hd__clkbuf_1 wire8071 (.A(net8072),
    .X(net8071));
 sky130_fd_sc_hd__clkbuf_1 wire8072 (.A(net8073),
    .X(net8072));
 sky130_fd_sc_hd__clkbuf_1 max_length8073 (.A(net8074),
    .X(net8073));
 sky130_fd_sc_hd__buf_1 wire8074 (.A(net8064),
    .X(net8074));
 sky130_fd_sc_hd__clkbuf_1 wire8075 (.A(net8076),
    .X(net8075));
 sky130_fd_sc_hd__clkbuf_1 wire8076 (.A(net8077),
    .X(net8076));
 sky130_fd_sc_hd__clkbuf_1 wire8077 (.A(net8078),
    .X(net8077));
 sky130_fd_sc_hd__clkbuf_1 wire8078 (.A(net8079),
    .X(net8078));
 sky130_fd_sc_hd__clkbuf_1 wire8079 (.A(net8080),
    .X(net8079));
 sky130_fd_sc_hd__clkbuf_1 wire8080 (.A(net8081),
    .X(net8080));
 sky130_fd_sc_hd__clkbuf_1 wire8081 (.A(net8082),
    .X(net8081));
 sky130_fd_sc_hd__clkbuf_1 wire8082 (.A(net8083),
    .X(net8082));
 sky130_fd_sc_hd__clkbuf_1 wire8083 (.A(net152),
    .X(net8083));
 sky130_fd_sc_hd__clkbuf_1 wire8084 (.A(net8085),
    .X(net8084));
 sky130_fd_sc_hd__clkbuf_1 wire8085 (.A(_02657_),
    .X(net8085));
 sky130_fd_sc_hd__clkbuf_1 wire8086 (.A(net8087),
    .X(net8086));
 sky130_fd_sc_hd__clkbuf_1 wire8087 (.A(net8088),
    .X(net8087));
 sky130_fd_sc_hd__clkbuf_1 wire8088 (.A(net8089),
    .X(net8088));
 sky130_fd_sc_hd__clkbuf_1 wire8089 (.A(net8090),
    .X(net8089));
 sky130_fd_sc_hd__clkbuf_1 wire8090 (.A(net8091),
    .X(net8090));
 sky130_fd_sc_hd__clkbuf_1 wire8091 (.A(net99),
    .X(net8091));
 sky130_fd_sc_hd__clkbuf_1 wire8092 (.A(net8093),
    .X(net8092));
 sky130_fd_sc_hd__clkbuf_1 wire8093 (.A(net8094),
    .X(net8093));
 sky130_fd_sc_hd__clkbuf_1 wire8094 (.A(net8095),
    .X(net8094));
 sky130_fd_sc_hd__clkbuf_1 wire8095 (.A(net98),
    .X(net8095));
 sky130_fd_sc_hd__clkbuf_1 wire8096 (.A(net8097),
    .X(net8096));
 sky130_fd_sc_hd__clkbuf_1 wire8097 (.A(net96),
    .X(net8097));
 sky130_fd_sc_hd__clkbuf_1 wire8098 (.A(net95),
    .X(net8098));
 sky130_fd_sc_hd__clkbuf_1 wire8099 (.A(net91),
    .X(net8099));
 sky130_fd_sc_hd__buf_1 wire8100 (.A(net9),
    .X(net8100));
 sky130_fd_sc_hd__clkbuf_1 wire8101 (.A(net89),
    .X(net8101));
 sky130_fd_sc_hd__clkbuf_1 wire8102 (.A(net88),
    .X(net8102));
 sky130_fd_sc_hd__clkbuf_1 wire8103 (.A(net8104),
    .X(net8103));
 sky130_fd_sc_hd__clkbuf_1 wire8104 (.A(net87),
    .X(net8104));
 sky130_fd_sc_hd__clkbuf_1 wire8105 (.A(net85),
    .X(net8105));
 sky130_fd_sc_hd__clkbuf_1 wire8106 (.A(net83),
    .X(net8106));
 sky130_fd_sc_hd__clkbuf_1 wire8107 (.A(net82),
    .X(net8107));
 sky130_fd_sc_hd__buf_1 wire8108 (.A(net8109),
    .X(net8108));
 sky130_fd_sc_hd__clkbuf_1 wire8109 (.A(net8110),
    .X(net8109));
 sky130_fd_sc_hd__clkbuf_1 wire8110 (.A(net8111),
    .X(net8110));
 sky130_fd_sc_hd__clkbuf_1 wire8111 (.A(net8112),
    .X(net8111));
 sky130_fd_sc_hd__clkbuf_1 wire8112 (.A(net8113),
    .X(net8112));
 sky130_fd_sc_hd__clkbuf_1 wire8113 (.A(net8114),
    .X(net8113));
 sky130_fd_sc_hd__clkbuf_1 wire8114 (.A(net8115),
    .X(net8114));
 sky130_fd_sc_hd__clkbuf_1 wire8115 (.A(net8116),
    .X(net8115));
 sky130_fd_sc_hd__clkbuf_1 wire8116 (.A(net8117),
    .X(net8116));
 sky130_fd_sc_hd__clkbuf_1 wire8117 (.A(net81),
    .X(net8117));
 sky130_fd_sc_hd__clkbuf_1 wire8118 (.A(net74),
    .X(net8118));
 sky130_fd_sc_hd__buf_1 wire8119 (.A(net7),
    .X(net8119));
 sky130_fd_sc_hd__clkbuf_2 fanout8120 (.A(net6),
    .X(net8120));
 sky130_fd_sc_hd__clkbuf_2 max_length8121 (.A(net8120),
    .X(net8121));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout8122 (.A(net6),
    .X(net8122));
 sky130_fd_sc_hd__clkbuf_1 wire8123 (.A(net8124),
    .X(net8123));
 sky130_fd_sc_hd__clkbuf_1 wire8124 (.A(net8125),
    .X(net8124));
 sky130_fd_sc_hd__clkbuf_1 wire8125 (.A(net8126),
    .X(net8125));
 sky130_fd_sc_hd__clkbuf_1 wire8126 (.A(net48),
    .X(net8126));
 sky130_fd_sc_hd__clkbuf_1 wire8127 (.A(net8128),
    .X(net8127));
 sky130_fd_sc_hd__clkbuf_1 wire8128 (.A(net8129),
    .X(net8128));
 sky130_fd_sc_hd__clkbuf_1 wire8129 (.A(net8130),
    .X(net8129));
 sky130_fd_sc_hd__clkbuf_1 wire8130 (.A(net8131),
    .X(net8130));
 sky130_fd_sc_hd__clkbuf_1 wire8131 (.A(net47),
    .X(net8131));
 sky130_fd_sc_hd__clkbuf_1 wire8132 (.A(net8133),
    .X(net8132));
 sky130_fd_sc_hd__clkbuf_1 wire8133 (.A(net8134),
    .X(net8133));
 sky130_fd_sc_hd__clkbuf_1 wire8134 (.A(net8135),
    .X(net8134));
 sky130_fd_sc_hd__clkbuf_1 wire8135 (.A(net46),
    .X(net8135));
 sky130_fd_sc_hd__clkbuf_1 wire8136 (.A(net8137),
    .X(net8136));
 sky130_fd_sc_hd__clkbuf_1 wire8137 (.A(net8138),
    .X(net8137));
 sky130_fd_sc_hd__clkbuf_1 wire8138 (.A(net8139),
    .X(net8138));
 sky130_fd_sc_hd__clkbuf_1 wire8139 (.A(net8140),
    .X(net8139));
 sky130_fd_sc_hd__clkbuf_1 wire8140 (.A(net45),
    .X(net8140));
 sky130_fd_sc_hd__clkbuf_1 wire8141 (.A(net8142),
    .X(net8141));
 sky130_fd_sc_hd__clkbuf_1 wire8142 (.A(net8143),
    .X(net8142));
 sky130_fd_sc_hd__clkbuf_1 wire8143 (.A(net8144),
    .X(net8143));
 sky130_fd_sc_hd__clkbuf_1 wire8144 (.A(net8145),
    .X(net8144));
 sky130_fd_sc_hd__clkbuf_1 wire8145 (.A(net44),
    .X(net8145));
 sky130_fd_sc_hd__clkbuf_1 wire8146 (.A(net8147),
    .X(net8146));
 sky130_fd_sc_hd__clkbuf_1 wire8147 (.A(net8148),
    .X(net8147));
 sky130_fd_sc_hd__clkbuf_1 wire8148 (.A(net8149),
    .X(net8148));
 sky130_fd_sc_hd__clkbuf_1 wire8149 (.A(net8150),
    .X(net8149));
 sky130_fd_sc_hd__clkbuf_1 wire8150 (.A(net43),
    .X(net8150));
 sky130_fd_sc_hd__clkbuf_1 wire8151 (.A(net8152),
    .X(net8151));
 sky130_fd_sc_hd__clkbuf_1 wire8152 (.A(net8153),
    .X(net8152));
 sky130_fd_sc_hd__clkbuf_1 wire8153 (.A(net8154),
    .X(net8153));
 sky130_fd_sc_hd__clkbuf_1 wire8154 (.A(net8155),
    .X(net8154));
 sky130_fd_sc_hd__clkbuf_1 wire8155 (.A(net8156),
    .X(net8155));
 sky130_fd_sc_hd__clkbuf_1 wire8156 (.A(net42),
    .X(net8156));
 sky130_fd_sc_hd__clkbuf_1 wire8157 (.A(net8158),
    .X(net8157));
 sky130_fd_sc_hd__clkbuf_1 wire8158 (.A(net8159),
    .X(net8158));
 sky130_fd_sc_hd__clkbuf_1 wire8159 (.A(net8160),
    .X(net8159));
 sky130_fd_sc_hd__clkbuf_1 wire8160 (.A(net8161),
    .X(net8160));
 sky130_fd_sc_hd__clkbuf_1 wire8161 (.A(net8162),
    .X(net8161));
 sky130_fd_sc_hd__clkbuf_1 wire8162 (.A(net41),
    .X(net8162));
 sky130_fd_sc_hd__clkbuf_1 wire8163 (.A(net8164),
    .X(net8163));
 sky130_fd_sc_hd__clkbuf_1 wire8164 (.A(net8165),
    .X(net8164));
 sky130_fd_sc_hd__clkbuf_1 wire8165 (.A(net8166),
    .X(net8165));
 sky130_fd_sc_hd__clkbuf_1 wire8166 (.A(net8167),
    .X(net8166));
 sky130_fd_sc_hd__clkbuf_1 wire8167 (.A(net40),
    .X(net8167));
 sky130_fd_sc_hd__clkbuf_1 wire8168 (.A(net8169),
    .X(net8168));
 sky130_fd_sc_hd__clkbuf_1 wire8169 (.A(net8170),
    .X(net8169));
 sky130_fd_sc_hd__clkbuf_1 wire8170 (.A(net8171),
    .X(net8170));
 sky130_fd_sc_hd__clkbuf_1 wire8171 (.A(net8172),
    .X(net8171));
 sky130_fd_sc_hd__clkbuf_1 wire8172 (.A(net8173),
    .X(net8172));
 sky130_fd_sc_hd__clkbuf_1 wire8173 (.A(net39),
    .X(net8173));
 sky130_fd_sc_hd__clkbuf_1 wire8174 (.A(net8175),
    .X(net8174));
 sky130_fd_sc_hd__clkbuf_1 wire8175 (.A(net8176),
    .X(net8175));
 sky130_fd_sc_hd__clkbuf_1 wire8176 (.A(net8177),
    .X(net8176));
 sky130_fd_sc_hd__clkbuf_1 wire8177 (.A(net8178),
    .X(net8177));
 sky130_fd_sc_hd__clkbuf_1 wire8178 (.A(net8179),
    .X(net8178));
 sky130_fd_sc_hd__clkbuf_1 wire8179 (.A(net38),
    .X(net8179));
 sky130_fd_sc_hd__clkbuf_1 wire8180 (.A(net8181),
    .X(net8180));
 sky130_fd_sc_hd__clkbuf_1 wire8181 (.A(net8182),
    .X(net8181));
 sky130_fd_sc_hd__clkbuf_1 wire8182 (.A(net8183),
    .X(net8182));
 sky130_fd_sc_hd__clkbuf_1 wire8183 (.A(net8184),
    .X(net8183));
 sky130_fd_sc_hd__clkbuf_1 wire8184 (.A(net8185),
    .X(net8184));
 sky130_fd_sc_hd__clkbuf_1 wire8185 (.A(net37),
    .X(net8185));
 sky130_fd_sc_hd__clkbuf_1 wire8186 (.A(net8187),
    .X(net8186));
 sky130_fd_sc_hd__clkbuf_1 wire8187 (.A(net8188),
    .X(net8187));
 sky130_fd_sc_hd__clkbuf_1 wire8188 (.A(net8189),
    .X(net8188));
 sky130_fd_sc_hd__clkbuf_1 wire8189 (.A(net36),
    .X(net8189));
 sky130_fd_sc_hd__clkbuf_1 wire8190 (.A(net8191),
    .X(net8190));
 sky130_fd_sc_hd__clkbuf_1 wire8191 (.A(net8192),
    .X(net8191));
 sky130_fd_sc_hd__clkbuf_1 wire8192 (.A(net8193),
    .X(net8192));
 sky130_fd_sc_hd__clkbuf_1 wire8193 (.A(net35),
    .X(net8193));
 sky130_fd_sc_hd__clkbuf_1 wire8194 (.A(net8195),
    .X(net8194));
 sky130_fd_sc_hd__clkbuf_1 wire8195 (.A(net8196),
    .X(net8195));
 sky130_fd_sc_hd__clkbuf_1 wire8196 (.A(net8197),
    .X(net8196));
 sky130_fd_sc_hd__clkbuf_1 wire8197 (.A(net34),
    .X(net8197));
 sky130_fd_sc_hd__clkbuf_1 wire8198 (.A(net8199),
    .X(net8198));
 sky130_fd_sc_hd__clkbuf_1 wire8199 (.A(net8200),
    .X(net8199));
 sky130_fd_sc_hd__clkbuf_1 wire8200 (.A(net8201),
    .X(net8200));
 sky130_fd_sc_hd__clkbuf_1 wire8201 (.A(net8202),
    .X(net8201));
 sky130_fd_sc_hd__clkbuf_1 wire8202 (.A(net8203),
    .X(net8202));
 sky130_fd_sc_hd__clkbuf_1 wire8203 (.A(net33),
    .X(net8203));
 sky130_fd_sc_hd__clkbuf_1 wire8204 (.A(net8205),
    .X(net8204));
 sky130_fd_sc_hd__clkbuf_1 wire8205 (.A(net8206),
    .X(net8205));
 sky130_fd_sc_hd__clkbuf_1 wire8206 (.A(net8207),
    .X(net8206));
 sky130_fd_sc_hd__clkbuf_1 wire8207 (.A(net8208),
    .X(net8207));
 sky130_fd_sc_hd__clkbuf_1 wire8208 (.A(net8209),
    .X(net8208));
 sky130_fd_sc_hd__clkbuf_1 wire8209 (.A(net32),
    .X(net8209));
 sky130_fd_sc_hd__clkbuf_1 wire8210 (.A(net8211),
    .X(net8210));
 sky130_fd_sc_hd__clkbuf_1 wire8211 (.A(net8212),
    .X(net8211));
 sky130_fd_sc_hd__clkbuf_1 wire8212 (.A(net8213),
    .X(net8212));
 sky130_fd_sc_hd__clkbuf_1 wire8213 (.A(net8214),
    .X(net8213));
 sky130_fd_sc_hd__clkbuf_1 wire8214 (.A(net8215),
    .X(net8214));
 sky130_fd_sc_hd__clkbuf_1 wire8215 (.A(net8216),
    .X(net8215));
 sky130_fd_sc_hd__clkbuf_1 wire8216 (.A(net31),
    .X(net8216));
 sky130_fd_sc_hd__clkbuf_1 wire8217 (.A(net8218),
    .X(net8217));
 sky130_fd_sc_hd__clkbuf_1 wire8218 (.A(net8219),
    .X(net8218));
 sky130_fd_sc_hd__clkbuf_1 wire8219 (.A(net8220),
    .X(net8219));
 sky130_fd_sc_hd__clkbuf_1 wire8220 (.A(net8221),
    .X(net8220));
 sky130_fd_sc_hd__clkbuf_1 wire8221 (.A(net8222),
    .X(net8221));
 sky130_fd_sc_hd__clkbuf_1 wire8222 (.A(net8223),
    .X(net8222));
 sky130_fd_sc_hd__clkbuf_1 wire8223 (.A(net8224),
    .X(net8223));
 sky130_fd_sc_hd__clkbuf_1 wire8224 (.A(net30),
    .X(net8224));
 sky130_fd_sc_hd__clkbuf_1 wire8225 (.A(net8226),
    .X(net8225));
 sky130_fd_sc_hd__clkbuf_1 wire8226 (.A(net8227),
    .X(net8226));
 sky130_fd_sc_hd__clkbuf_1 wire8227 (.A(net8228),
    .X(net8227));
 sky130_fd_sc_hd__clkbuf_1 wire8228 (.A(net8229),
    .X(net8228));
 sky130_fd_sc_hd__clkbuf_1 wire8229 (.A(net8230),
    .X(net8229));
 sky130_fd_sc_hd__clkbuf_1 wire8230 (.A(net8231),
    .X(net8230));
 sky130_fd_sc_hd__clkbuf_1 wire8231 (.A(net8232),
    .X(net8231));
 sky130_fd_sc_hd__clkbuf_1 wire8232 (.A(net29),
    .X(net8232));
 sky130_fd_sc_hd__clkbuf_1 wire8233 (.A(net8234),
    .X(net8233));
 sky130_fd_sc_hd__clkbuf_1 wire8234 (.A(net8235),
    .X(net8234));
 sky130_fd_sc_hd__clkbuf_1 wire8235 (.A(net8236),
    .X(net8235));
 sky130_fd_sc_hd__clkbuf_1 wire8236 (.A(net8237),
    .X(net8236));
 sky130_fd_sc_hd__clkbuf_1 wire8237 (.A(net8238),
    .X(net8237));
 sky130_fd_sc_hd__clkbuf_1 wire8238 (.A(net8239),
    .X(net8238));
 sky130_fd_sc_hd__clkbuf_1 wire8239 (.A(net8240),
    .X(net8239));
 sky130_fd_sc_hd__clkbuf_1 wire8240 (.A(net8241),
    .X(net8240));
 sky130_fd_sc_hd__clkbuf_1 wire8241 (.A(net8242),
    .X(net8241));
 sky130_fd_sc_hd__clkbuf_1 wire8242 (.A(net28),
    .X(net8242));
 sky130_fd_sc_hd__clkbuf_1 wire8243 (.A(net8244),
    .X(net8243));
 sky130_fd_sc_hd__clkbuf_1 wire8244 (.A(net8245),
    .X(net8244));
 sky130_fd_sc_hd__clkbuf_1 wire8245 (.A(net8246),
    .X(net8245));
 sky130_fd_sc_hd__clkbuf_1 wire8246 (.A(net8247),
    .X(net8246));
 sky130_fd_sc_hd__clkbuf_1 wire8247 (.A(net8248),
    .X(net8247));
 sky130_fd_sc_hd__clkbuf_1 wire8248 (.A(net8249),
    .X(net8248));
 sky130_fd_sc_hd__clkbuf_1 wire8249 (.A(net8250),
    .X(net8249));
 sky130_fd_sc_hd__clkbuf_1 wire8250 (.A(net8251),
    .X(net8250));
 sky130_fd_sc_hd__clkbuf_1 wire8251 (.A(net8252),
    .X(net8251));
 sky130_fd_sc_hd__clkbuf_1 wire8252 (.A(net27),
    .X(net8252));
 sky130_fd_sc_hd__clkbuf_1 wire8253 (.A(net8254),
    .X(net8253));
 sky130_fd_sc_hd__clkbuf_1 wire8254 (.A(net8255),
    .X(net8254));
 sky130_fd_sc_hd__clkbuf_1 wire8255 (.A(net8256),
    .X(net8255));
 sky130_fd_sc_hd__clkbuf_1 wire8256 (.A(net8257),
    .X(net8256));
 sky130_fd_sc_hd__clkbuf_1 wire8257 (.A(net8258),
    .X(net8257));
 sky130_fd_sc_hd__clkbuf_1 wire8258 (.A(net8259),
    .X(net8258));
 sky130_fd_sc_hd__clkbuf_1 wire8259 (.A(net8260),
    .X(net8259));
 sky130_fd_sc_hd__clkbuf_1 wire8260 (.A(net8261),
    .X(net8260));
 sky130_fd_sc_hd__clkbuf_1 wire8261 (.A(net26),
    .X(net8261));
 sky130_fd_sc_hd__clkbuf_1 wire8262 (.A(net8263),
    .X(net8262));
 sky130_fd_sc_hd__clkbuf_1 wire8263 (.A(net8264),
    .X(net8263));
 sky130_fd_sc_hd__clkbuf_1 wire8264 (.A(net8265),
    .X(net8264));
 sky130_fd_sc_hd__clkbuf_1 wire8265 (.A(net8266),
    .X(net8265));
 sky130_fd_sc_hd__clkbuf_1 wire8266 (.A(net8267),
    .X(net8266));
 sky130_fd_sc_hd__clkbuf_1 wire8267 (.A(net8268),
    .X(net8267));
 sky130_fd_sc_hd__clkbuf_1 wire8268 (.A(net8269),
    .X(net8268));
 sky130_fd_sc_hd__clkbuf_1 wire8269 (.A(net8270),
    .X(net8269));
 sky130_fd_sc_hd__clkbuf_1 wire8270 (.A(net25),
    .X(net8270));
 sky130_fd_sc_hd__clkbuf_1 wire8271 (.A(net8272),
    .X(net8271));
 sky130_fd_sc_hd__clkbuf_1 wire8272 (.A(net8273),
    .X(net8272));
 sky130_fd_sc_hd__clkbuf_1 wire8273 (.A(net8274),
    .X(net8273));
 sky130_fd_sc_hd__clkbuf_1 wire8274 (.A(net8275),
    .X(net8274));
 sky130_fd_sc_hd__clkbuf_1 wire8275 (.A(net8276),
    .X(net8275));
 sky130_fd_sc_hd__clkbuf_1 wire8276 (.A(net8277),
    .X(net8276));
 sky130_fd_sc_hd__clkbuf_1 wire8277 (.A(net8278),
    .X(net8277));
 sky130_fd_sc_hd__clkbuf_1 wire8278 (.A(net8279),
    .X(net8278));
 sky130_fd_sc_hd__clkbuf_1 wire8279 (.A(net24),
    .X(net8279));
 sky130_fd_sc_hd__clkbuf_1 wire8280 (.A(net8281),
    .X(net8280));
 sky130_fd_sc_hd__clkbuf_1 wire8281 (.A(net8282),
    .X(net8281));
 sky130_fd_sc_hd__clkbuf_1 wire8282 (.A(net8283),
    .X(net8282));
 sky130_fd_sc_hd__clkbuf_1 wire8283 (.A(net8284),
    .X(net8283));
 sky130_fd_sc_hd__clkbuf_1 wire8284 (.A(net23),
    .X(net8284));
 sky130_fd_sc_hd__clkbuf_1 wire8285 (.A(net8286),
    .X(net8285));
 sky130_fd_sc_hd__clkbuf_1 wire8286 (.A(net8287),
    .X(net8286));
 sky130_fd_sc_hd__clkbuf_1 wire8287 (.A(net8288),
    .X(net8287));
 sky130_fd_sc_hd__clkbuf_1 wire8288 (.A(net8289),
    .X(net8288));
 sky130_fd_sc_hd__clkbuf_1 wire8289 (.A(net22),
    .X(net8289));
 sky130_fd_sc_hd__clkbuf_1 wire8290 (.A(net8291),
    .X(net8290));
 sky130_fd_sc_hd__clkbuf_1 wire8291 (.A(net8292),
    .X(net8291));
 sky130_fd_sc_hd__clkbuf_1 wire8292 (.A(net8293),
    .X(net8292));
 sky130_fd_sc_hd__clkbuf_1 wire8293 (.A(net8294),
    .X(net8293));
 sky130_fd_sc_hd__clkbuf_1 wire8294 (.A(net21),
    .X(net8294));
 sky130_fd_sc_hd__clkbuf_1 wire8295 (.A(net8296),
    .X(net8295));
 sky130_fd_sc_hd__clkbuf_1 wire8296 (.A(net8297),
    .X(net8296));
 sky130_fd_sc_hd__clkbuf_1 wire8297 (.A(net8298),
    .X(net8297));
 sky130_fd_sc_hd__clkbuf_1 wire8298 (.A(net8299),
    .X(net8298));
 sky130_fd_sc_hd__clkbuf_1 wire8299 (.A(net20),
    .X(net8299));
 sky130_fd_sc_hd__clkbuf_1 wire8300 (.A(net8301),
    .X(net8300));
 sky130_fd_sc_hd__clkbuf_1 wire8301 (.A(net8302),
    .X(net8301));
 sky130_fd_sc_hd__clkbuf_1 wire8302 (.A(net8303),
    .X(net8302));
 sky130_fd_sc_hd__clkbuf_1 wire8303 (.A(net8304),
    .X(net8303));
 sky130_fd_sc_hd__clkbuf_1 wire8304 (.A(net19),
    .X(net8304));
 sky130_fd_sc_hd__clkbuf_1 wire8305 (.A(net8306),
    .X(net8305));
 sky130_fd_sc_hd__clkbuf_1 wire8306 (.A(net8307),
    .X(net8306));
 sky130_fd_sc_hd__clkbuf_1 wire8307 (.A(net8308),
    .X(net8307));
 sky130_fd_sc_hd__clkbuf_1 wire8308 (.A(net8309),
    .X(net8308));
 sky130_fd_sc_hd__clkbuf_1 wire8309 (.A(net8310),
    .X(net8309));
 sky130_fd_sc_hd__clkbuf_1 wire8310 (.A(net8311),
    .X(net8310));
 sky130_fd_sc_hd__clkbuf_1 wire8311 (.A(net18),
    .X(net8311));
 sky130_fd_sc_hd__clkbuf_1 wire8312 (.A(net8313),
    .X(net8312));
 sky130_fd_sc_hd__clkbuf_1 wire8313 (.A(net8314),
    .X(net8313));
 sky130_fd_sc_hd__clkbuf_1 wire8314 (.A(net8315),
    .X(net8314));
 sky130_fd_sc_hd__clkbuf_1 wire8315 (.A(net8316),
    .X(net8315));
 sky130_fd_sc_hd__clkbuf_1 wire8316 (.A(net8317),
    .X(net8316));
 sky130_fd_sc_hd__clkbuf_1 wire8317 (.A(net8318),
    .X(net8317));
 sky130_fd_sc_hd__clkbuf_1 wire8318 (.A(net17),
    .X(net8318));
 sky130_fd_sc_hd__clkbuf_1 wire8319 (.A(net8320),
    .X(net8319));
 sky130_fd_sc_hd__clkbuf_1 wire8320 (.A(net8321),
    .X(net8320));
 sky130_fd_sc_hd__clkbuf_1 wire8321 (.A(net8322),
    .X(net8321));
 sky130_fd_sc_hd__clkbuf_1 wire8322 (.A(net8323),
    .X(net8322));
 sky130_fd_sc_hd__clkbuf_1 wire8323 (.A(net8324),
    .X(net8323));
 sky130_fd_sc_hd__clkbuf_1 wire8324 (.A(net8325),
    .X(net8324));
 sky130_fd_sc_hd__clkbuf_1 wire8325 (.A(net8326),
    .X(net8325));
 sky130_fd_sc_hd__clkbuf_1 wire8326 (.A(net8327),
    .X(net8326));
 sky130_fd_sc_hd__clkbuf_1 wire8327 (.A(net148),
    .X(net8327));
 sky130_fd_sc_hd__clkbuf_1 fanout8328 (.A(net8339),
    .X(net8328));
 sky130_fd_sc_hd__buf_1 wire8329 (.A(net8331),
    .X(net8329));
 sky130_fd_sc_hd__clkbuf_1 wire8330 (.A(net8331),
    .X(net8330));
 sky130_fd_sc_hd__buf_1 wire8331 (.A(net8332),
    .X(net8331));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8332 (.A(net8328),
    .X(net8332));
 sky130_fd_sc_hd__clkbuf_1 wire8333 (.A(net8328),
    .X(net8333));
 sky130_fd_sc_hd__buf_1 fanout8334 (.A(net8339),
    .X(net8334));
 sky130_fd_sc_hd__buf_1 max_length8335 (.A(net8336),
    .X(net8335));
 sky130_fd_sc_hd__buf_1 wire8336 (.A(net8337),
    .X(net8336));
 sky130_fd_sc_hd__buf_1 wire8337 (.A(net8334),
    .X(net8337));
 sky130_fd_sc_hd__buf_1 fanout8338 (.A(net8538),
    .X(net8338));
 sky130_fd_sc_hd__buf_1 wire8339 (.A(net8340),
    .X(net8339));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8340 (.A(net8338),
    .X(net8340));
 sky130_fd_sc_hd__buf_1 max_length8341 (.A(net8342),
    .X(net8341));
 sky130_fd_sc_hd__buf_1 max_length8342 (.A(net8338),
    .X(net8342));
 sky130_fd_sc_hd__buf_1 fanout8343 (.A(net8348),
    .X(net8343));
 sky130_fd_sc_hd__buf_1 wire8344 (.A(net8345),
    .X(net8344));
 sky130_fd_sc_hd__buf_1 max_length8345 (.A(net8346),
    .X(net8345));
 sky130_fd_sc_hd__buf_1 wire8346 (.A(net8343),
    .X(net8346));
 sky130_fd_sc_hd__buf_1 max_length8347 (.A(net8343),
    .X(net8347));
 sky130_fd_sc_hd__buf_1 fanout8348 (.A(net8370),
    .X(net8348));
 sky130_fd_sc_hd__buf_1 wire8349 (.A(net8352),
    .X(net8349));
 sky130_fd_sc_hd__buf_1 wire8350 (.A(net8351),
    .X(net8350));
 sky130_fd_sc_hd__buf_1 max_length8351 (.A(net8352),
    .X(net8351));
 sky130_fd_sc_hd__buf_1 wire8352 (.A(net8348),
    .X(net8352));
 sky130_fd_sc_hd__buf_1 fanout8353 (.A(net8360),
    .X(net8353));
 sky130_fd_sc_hd__buf_1 wire8354 (.A(net8356),
    .X(net8354));
 sky130_fd_sc_hd__buf_1 max_length8355 (.A(net8356),
    .X(net8355));
 sky130_fd_sc_hd__clkbuf_2 max_length8356 (.A(net8353),
    .X(net8356));
 sky130_fd_sc_hd__buf_1 fanout8357 (.A(net8361),
    .X(net8357));
 sky130_fd_sc_hd__buf_1 wire8358 (.A(net8357),
    .X(net8358));
 sky130_fd_sc_hd__clkbuf_1 fanout8359 (.A(net8374),
    .X(net8359));
 sky130_fd_sc_hd__clkbuf_1 wire8360 (.A(net8361),
    .X(net8360));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8361 (.A(net8359),
    .X(net8361));
 sky130_fd_sc_hd__buf_1 fanout8362 (.A(net8369),
    .X(net8362));
 sky130_fd_sc_hd__clkbuf_1 wire8363 (.A(net8364),
    .X(net8363));
 sky130_fd_sc_hd__buf_1 wire8364 (.A(net8365),
    .X(net8364));
 sky130_fd_sc_hd__buf_1 wire8365 (.A(net8366),
    .X(net8365));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8366 (.A(net8367),
    .X(net8366));
 sky130_fd_sc_hd__buf_1 wire8367 (.A(net8368),
    .X(net8367));
 sky130_fd_sc_hd__buf_1 wire8368 (.A(net8362),
    .X(net8368));
 sky130_fd_sc_hd__buf_1 fanout8369 (.A(net8540),
    .X(net8369));
 sky130_fd_sc_hd__clkbuf_1 wire8370 (.A(net8371),
    .X(net8370));
 sky130_fd_sc_hd__clkbuf_1 wire8371 (.A(net8372),
    .X(net8371));
 sky130_fd_sc_hd__clkbuf_1 wire8372 (.A(net8373),
    .X(net8372));
 sky130_fd_sc_hd__clkbuf_1 wire8373 (.A(net8369),
    .X(net8373));
 sky130_fd_sc_hd__clkbuf_1 wire8374 (.A(net8375),
    .X(net8374));
 sky130_fd_sc_hd__buf_1 wire8375 (.A(net8376),
    .X(net8375));
 sky130_fd_sc_hd__buf_1 wire8376 (.A(net8377),
    .X(net8376));
 sky130_fd_sc_hd__clkbuf_1 wire8377 (.A(net8378),
    .X(net8377));
 sky130_fd_sc_hd__clkbuf_1 wire8378 (.A(net8379),
    .X(net8378));
 sky130_fd_sc_hd__clkbuf_1 max_length8379 (.A(net8369),
    .X(net8379));
 sky130_fd_sc_hd__buf_1 fanout8380 (.A(net8386),
    .X(net8380));
 sky130_fd_sc_hd__buf_1 max_length8381 (.A(net8382),
    .X(net8381));
 sky130_fd_sc_hd__clkbuf_2 wire8382 (.A(net8380),
    .X(net8382));
 sky130_fd_sc_hd__clkbuf_2 fanout8383 (.A(net8386),
    .X(net8383));
 sky130_fd_sc_hd__buf_1 wire8384 (.A(net8383),
    .X(net8384));
 sky130_fd_sc_hd__buf_1 fanout8385 (.A(net8393),
    .X(net8385));
 sky130_fd_sc_hd__buf_1 wire8386 (.A(net8385),
    .X(net8386));
 sky130_fd_sc_hd__buf_1 wire8387 (.A(net8385),
    .X(net8387));
 sky130_fd_sc_hd__clkbuf_1 fanout8388 (.A(net8415),
    .X(net8388));
 sky130_fd_sc_hd__buf_1 wire8389 (.A(net8390),
    .X(net8389));
 sky130_fd_sc_hd__clkbuf_2 wire8390 (.A(net8391),
    .X(net8390));
 sky130_fd_sc_hd__clkbuf_1 wire8391 (.A(net8392),
    .X(net8391));
 sky130_fd_sc_hd__clkbuf_1 wire8392 (.A(net8393),
    .X(net8392));
 sky130_fd_sc_hd__buf_1 wire8393 (.A(net8388),
    .X(net8393));
 sky130_fd_sc_hd__buf_1 fanout8394 (.A(net8414),
    .X(net8394));
 sky130_fd_sc_hd__clkbuf_2 wire8395 (.A(net8394),
    .X(net8395));
 sky130_fd_sc_hd__buf_1 wire8396 (.A(net8397),
    .X(net8396));
 sky130_fd_sc_hd__buf_1 max_length8397 (.A(net8394),
    .X(net8397));
 sky130_fd_sc_hd__clkbuf_2 fanout8398 (.A(net8411),
    .X(net8398));
 sky130_fd_sc_hd__buf_1 wire8399 (.A(net8400),
    .X(net8399));
 sky130_fd_sc_hd__buf_1 wire8400 (.A(net8398),
    .X(net8400));
 sky130_fd_sc_hd__buf_1 fanout8401 (.A(net8408),
    .X(net8401));
 sky130_fd_sc_hd__buf_1 wire8402 (.A(net8403),
    .X(net8402));
 sky130_fd_sc_hd__clkbuf_2 wire8403 (.A(net8404),
    .X(net8403));
 sky130_fd_sc_hd__clkbuf_2 wire8404 (.A(net8401),
    .X(net8404));
 sky130_fd_sc_hd__clkbuf_2 fanout8405 (.A(net8410),
    .X(net8405));
 sky130_fd_sc_hd__buf_1 max_length8406 (.A(net8407),
    .X(net8406));
 sky130_fd_sc_hd__buf_1 wire8407 (.A(net8405),
    .X(net8407));
 sky130_fd_sc_hd__clkbuf_1 max_length8408 (.A(net8405),
    .X(net8408));
 sky130_fd_sc_hd__clkbuf_2 max_length8409 (.A(net8405),
    .X(net8409));
 sky130_fd_sc_hd__clkbuf_1 fanout8410 (.A(net8418),
    .X(net8410));
 sky130_fd_sc_hd__clkbuf_1 wire8411 (.A(net8412),
    .X(net8411));
 sky130_fd_sc_hd__buf_1 wire8412 (.A(net8413),
    .X(net8412));
 sky130_fd_sc_hd__buf_1 wire8413 (.A(net8410),
    .X(net8413));
 sky130_fd_sc_hd__buf_1 fanout8414 (.A(net8537),
    .X(net8414));
 sky130_fd_sc_hd__clkbuf_1 wire8415 (.A(net8416),
    .X(net8415));
 sky130_fd_sc_hd__clkbuf_1 wire8416 (.A(net8417),
    .X(net8416));
 sky130_fd_sc_hd__clkbuf_1 max_length8417 (.A(net8418),
    .X(net8417));
 sky130_fd_sc_hd__buf_1 wire8418 (.A(net8419),
    .X(net8418));
 sky130_fd_sc_hd__buf_1 wire8419 (.A(net8414),
    .X(net8419));
 sky130_fd_sc_hd__clkbuf_2 fanout8420 (.A(net8424),
    .X(net8420));
 sky130_fd_sc_hd__buf_1 wire8421 (.A(net8422),
    .X(net8421));
 sky130_fd_sc_hd__clkbuf_2 wire8422 (.A(net8420),
    .X(net8422));
 sky130_fd_sc_hd__buf_1 fanout8423 (.A(net8521),
    .X(net8423));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8424 (.A(net8425),
    .X(net8424));
 sky130_fd_sc_hd__clkbuf_2 max_length8425 (.A(net8423),
    .X(net8425));
 sky130_fd_sc_hd__buf_1 fanout8426 (.A(net8432),
    .X(net8426));
 sky130_fd_sc_hd__clkbuf_2 max_length8427 (.A(net8428),
    .X(net8427));
 sky130_fd_sc_hd__clkbuf_2 wire8428 (.A(net8426),
    .X(net8428));
 sky130_fd_sc_hd__clkbuf_2 fanout8429 (.A(net8434),
    .X(net8429));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8430 (.A(net8429),
    .X(net8430));
 sky130_fd_sc_hd__clkbuf_2 wire8431 (.A(net8429),
    .X(net8431));
 sky130_fd_sc_hd__buf_1 fanout8432 (.A(net8522),
    .X(net8432));
 sky130_fd_sc_hd__clkbuf_1 max_length8433 (.A(net8434),
    .X(net8433));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8434 (.A(net8432),
    .X(net8434));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout8435 (.A(net8438),
    .X(net8435));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8436 (.A(net8437),
    .X(net8436));
 sky130_fd_sc_hd__buf_1 wire8437 (.A(net8435),
    .X(net8437));
 sky130_fd_sc_hd__buf_1 fanout8438 (.A(net8441),
    .X(net8438));
 sky130_fd_sc_hd__clkbuf_2 wire8439 (.A(net8440),
    .X(net8439));
 sky130_fd_sc_hd__buf_1 wire8440 (.A(net8438),
    .X(net8440));
 sky130_fd_sc_hd__clkbuf_1 fanout8441 (.A(net8519),
    .X(net8441));
 sky130_fd_sc_hd__buf_1 wire8442 (.A(net8444),
    .X(net8442));
 sky130_fd_sc_hd__buf_1 max_length8443 (.A(net8444),
    .X(net8443));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8444 (.A(net8441),
    .X(net8444));
 sky130_fd_sc_hd__buf_1 fanout8445 (.A(net8480),
    .X(net8445));
 sky130_fd_sc_hd__clkbuf_1 wire8446 (.A(net8449),
    .X(net8446));
 sky130_fd_sc_hd__buf_1 wire8447 (.A(net8448),
    .X(net8447));
 sky130_fd_sc_hd__buf_1 wire8448 (.A(net8449),
    .X(net8448));
 sky130_fd_sc_hd__buf_1 wire8449 (.A(net8445),
    .X(net8449));
 sky130_fd_sc_hd__clkbuf_2 fanout8450 (.A(net8456),
    .X(net8450));
 sky130_fd_sc_hd__buf_1 wire8451 (.A(net8450),
    .X(net8451));
 sky130_fd_sc_hd__clkbuf_2 max_length8452 (.A(net8450),
    .X(net8452));
 sky130_fd_sc_hd__buf_1 fanout8453 (.A(net8479),
    .X(net8453));
 sky130_fd_sc_hd__buf_1 wire8454 (.A(net8456),
    .X(net8454));
 sky130_fd_sc_hd__clkbuf_2 max_length8455 (.A(net8456),
    .X(net8455));
 sky130_fd_sc_hd__buf_1 wire8456 (.A(net8453),
    .X(net8456));
 sky130_fd_sc_hd__clkbuf_2 fanout8457 (.A(net8459),
    .X(net8457));
 sky130_fd_sc_hd__clkbuf_2 wire8458 (.A(net8457),
    .X(net8458));
 sky130_fd_sc_hd__clkbuf_2 fanout8459 (.A(net8484),
    .X(net8459));
 sky130_fd_sc_hd__buf_1 wire8460 (.A(net8461),
    .X(net8460));
 sky130_fd_sc_hd__clkbuf_2 max_length8461 (.A(net8459),
    .X(net8461));
 sky130_fd_sc_hd__clkbuf_2 fanout8462 (.A(net8483),
    .X(net8462));
 sky130_fd_sc_hd__buf_1 wire8463 (.A(net8462),
    .X(net8463));
 sky130_fd_sc_hd__clkbuf_2 wire8464 (.A(net8462),
    .X(net8464));
 sky130_fd_sc_hd__clkbuf_1 fanout8465 (.A(net8483),
    .X(net8465));
 sky130_fd_sc_hd__clkbuf_2 max_length8466 (.A(net8467),
    .X(net8466));
 sky130_fd_sc_hd__buf_1 wire8467 (.A(net8465),
    .X(net8467));
 sky130_fd_sc_hd__clkbuf_2 fanout8468 (.A(net8475),
    .X(net8468));
 sky130_fd_sc_hd__clkbuf_2 wire8469 (.A(net8468),
    .X(net8469));
 sky130_fd_sc_hd__buf_1 wire8470 (.A(net8468),
    .X(net8470));
 sky130_fd_sc_hd__buf_1 fanout8471 (.A(net8476),
    .X(net8471));
 sky130_fd_sc_hd__buf_1 wire8472 (.A(net8471),
    .X(net8472));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8473 (.A(net8474),
    .X(net8473));
 sky130_fd_sc_hd__buf_1 max_length8474 (.A(net8471),
    .X(net8474));
 sky130_fd_sc_hd__clkbuf_1 fanout8475 (.A(net8486),
    .X(net8475));
 sky130_fd_sc_hd__buf_1 wire8476 (.A(net8477),
    .X(net8476));
 sky130_fd_sc_hd__clkbuf_2 max_length8477 (.A(net8478),
    .X(net8477));
 sky130_fd_sc_hd__buf_1 wire8478 (.A(net8475),
    .X(net8478));
 sky130_fd_sc_hd__buf_1 fanout8479 (.A(net8529),
    .X(net8479));
 sky130_fd_sc_hd__clkbuf_1 wire8480 (.A(net8481),
    .X(net8480));
 sky130_fd_sc_hd__clkbuf_1 wire8481 (.A(net8482),
    .X(net8481));
 sky130_fd_sc_hd__clkbuf_1 wire8482 (.A(net8479),
    .X(net8482));
 sky130_fd_sc_hd__buf_1 wire8483 (.A(net8485),
    .X(net8483));
 sky130_fd_sc_hd__buf_1 max_length8484 (.A(net8485),
    .X(net8484));
 sky130_fd_sc_hd__clkbuf_1 wire8485 (.A(net8486),
    .X(net8485));
 sky130_fd_sc_hd__buf_1 wire8486 (.A(net8487),
    .X(net8486));
 sky130_fd_sc_hd__clkbuf_1 max_length8487 (.A(net8479),
    .X(net8487));
 sky130_fd_sc_hd__buf_1 fanout8488 (.A(net8494),
    .X(net8488));
 sky130_fd_sc_hd__buf_1 wire8489 (.A(net8488),
    .X(net8489));
 sky130_fd_sc_hd__buf_1 wire8490 (.A(net8491),
    .X(net8490));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8491 (.A(net8488),
    .X(net8491));
 sky130_fd_sc_hd__clkbuf_1 fanout8492 (.A(net8509),
    .X(net8492));
 sky130_fd_sc_hd__buf_1 wire8493 (.A(net8494),
    .X(net8493));
 sky130_fd_sc_hd__buf_1 wire8494 (.A(net8492),
    .X(net8494));
 sky130_fd_sc_hd__buf_1 fanout8495 (.A(net8504),
    .X(net8495));
 sky130_fd_sc_hd__clkbuf_2 max_length8496 (.A(net8497),
    .X(net8496));
 sky130_fd_sc_hd__buf_1 wire8497 (.A(net8498),
    .X(net8497));
 sky130_fd_sc_hd__clkbuf_2 max_length8498 (.A(net8495),
    .X(net8498));
 sky130_fd_sc_hd__buf_1 fanout8499 (.A(net8501),
    .X(net8499));
 sky130_fd_sc_hd__clkbuf_2 wire8500 (.A(net8499),
    .X(net8500));
 sky130_fd_sc_hd__clkbuf_1 fanout8501 (.A(net8505),
    .X(net8501));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8502 (.A(net8503),
    .X(net8502));
 sky130_fd_sc_hd__clkbuf_2 wire8503 (.A(net8504),
    .X(net8503));
 sky130_fd_sc_hd__buf_1 wire8504 (.A(net8501),
    .X(net8504));
 sky130_fd_sc_hd__buf_1 fanout8505 (.A(net8517),
    .X(net8505));
 sky130_fd_sc_hd__buf_1 wire8506 (.A(net8507),
    .X(net8506));
 sky130_fd_sc_hd__clkbuf_2 wire8507 (.A(net8508),
    .X(net8507));
 sky130_fd_sc_hd__buf_1 wire8508 (.A(net8509),
    .X(net8508));
 sky130_fd_sc_hd__buf_1 wire8509 (.A(net8505),
    .X(net8509));
 sky130_fd_sc_hd__buf_1 fanout8510 (.A(net8525),
    .X(net8510));
 sky130_fd_sc_hd__clkbuf_2 wire8511 (.A(net8512),
    .X(net8511));
 sky130_fd_sc_hd__clkbuf_1 wire8512 (.A(net8517),
    .X(net8512));
 sky130_fd_sc_hd__clkbuf_1 wire8513 (.A(net8514),
    .X(net8513));
 sky130_fd_sc_hd__clkbuf_1 wire8514 (.A(net8515),
    .X(net8514));
 sky130_fd_sc_hd__clkbuf_1 wire8515 (.A(net8516),
    .X(net8515));
 sky130_fd_sc_hd__clkbuf_1 wire8516 (.A(net8510),
    .X(net8516));
 sky130_fd_sc_hd__buf_1 max_length8517 (.A(net8510),
    .X(net8517));
 sky130_fd_sc_hd__buf_1 fanout8518 (.A(net8530),
    .X(net8518));
 sky130_fd_sc_hd__clkbuf_1 wire8519 (.A(net8520),
    .X(net8519));
 sky130_fd_sc_hd__clkbuf_1 wire8520 (.A(net8523),
    .X(net8520));
 sky130_fd_sc_hd__clkbuf_1 wire8521 (.A(net8522),
    .X(net8521));
 sky130_fd_sc_hd__buf_1 wire8522 (.A(net8523),
    .X(net8522));
 sky130_fd_sc_hd__buf_1 wire8523 (.A(net8524),
    .X(net8523));
 sky130_fd_sc_hd__clkbuf_1 wire8524 (.A(net8529),
    .X(net8524));
 sky130_fd_sc_hd__clkbuf_1 wire8525 (.A(net8526),
    .X(net8525));
 sky130_fd_sc_hd__clkbuf_1 wire8526 (.A(net8527),
    .X(net8526));
 sky130_fd_sc_hd__clkbuf_1 wire8527 (.A(net8528),
    .X(net8527));
 sky130_fd_sc_hd__clkbuf_1 wire8528 (.A(net8518),
    .X(net8528));
 sky130_fd_sc_hd__clkbuf_1 max_length8529 (.A(net8518),
    .X(net8529));
 sky130_fd_sc_hd__buf_1 fanout8530 (.A(net8546),
    .X(net8530));
 sky130_fd_sc_hd__clkbuf_2 wire8531 (.A(net8532),
    .X(net8531));
 sky130_fd_sc_hd__clkbuf_2 wire8532 (.A(net8533),
    .X(net8532));
 sky130_fd_sc_hd__clkbuf_1 wire8533 (.A(net8534),
    .X(net8533));
 sky130_fd_sc_hd__clkbuf_1 wire8534 (.A(net8535),
    .X(net8534));
 sky130_fd_sc_hd__clkbuf_1 wire8535 (.A(net8536),
    .X(net8535));
 sky130_fd_sc_hd__clkbuf_1 wire8536 (.A(net8530),
    .X(net8536));
 sky130_fd_sc_hd__buf_1 fanout8537 (.A(net8844),
    .X(net8537));
 sky130_fd_sc_hd__clkbuf_1 wire8538 (.A(net8539),
    .X(net8538));
 sky130_fd_sc_hd__buf_1 wire8539 (.A(net8540),
    .X(net8539));
 sky130_fd_sc_hd__buf_1 wire8540 (.A(net8541),
    .X(net8540));
 sky130_fd_sc_hd__clkbuf_1 wire8541 (.A(net8542),
    .X(net8541));
 sky130_fd_sc_hd__clkbuf_1 wire8542 (.A(net8543),
    .X(net8542));
 sky130_fd_sc_hd__clkbuf_1 wire8543 (.A(net8544),
    .X(net8543));
 sky130_fd_sc_hd__clkbuf_1 wire8544 (.A(net8545),
    .X(net8544));
 sky130_fd_sc_hd__clkbuf_1 wire8545 (.A(net8537),
    .X(net8545));
 sky130_fd_sc_hd__clkbuf_1 wire8546 (.A(net8547),
    .X(net8546));
 sky130_fd_sc_hd__clkbuf_1 wire8547 (.A(net8548),
    .X(net8547));
 sky130_fd_sc_hd__clkbuf_1 wire8548 (.A(net8549),
    .X(net8548));
 sky130_fd_sc_hd__clkbuf_1 wire8549 (.A(net8550),
    .X(net8549));
 sky130_fd_sc_hd__clkbuf_1 wire8550 (.A(net8537),
    .X(net8550));
 sky130_fd_sc_hd__buf_1 fanout8551 (.A(net8554),
    .X(net8551));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8552 (.A(net8553),
    .X(net8552));
 sky130_fd_sc_hd__clkbuf_2 wire8553 (.A(net8551),
    .X(net8553));
 sky130_fd_sc_hd__clkbuf_2 fanout8554 (.A(net8560),
    .X(net8554));
 sky130_fd_sc_hd__buf_1 fanout8555 (.A(net8590),
    .X(net8555));
 sky130_fd_sc_hd__clkbuf_1 wire8556 (.A(net8557),
    .X(net8556));
 sky130_fd_sc_hd__clkbuf_1 wire8557 (.A(net8558),
    .X(net8557));
 sky130_fd_sc_hd__clkbuf_1 wire8558 (.A(net8559),
    .X(net8558));
 sky130_fd_sc_hd__clkbuf_2 wire8559 (.A(net8560),
    .X(net8559));
 sky130_fd_sc_hd__clkbuf_2 wire8560 (.A(net8555),
    .X(net8560));
 sky130_fd_sc_hd__clkbuf_2 fanout8561 (.A(net8564),
    .X(net8561));
 sky130_fd_sc_hd__clkbuf_2 wire8562 (.A(net8561),
    .X(net8562));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_length8563 (.A(net8561),
    .X(net8563));
 sky130_fd_sc_hd__buf_1 fanout8564 (.A(net8594),
    .X(net8564));
 sky130_fd_sc_hd__buf_1 max_length8565 (.A(net8566),
    .X(net8565));
 sky130_fd_sc_hd__buf_1 max_length8566 (.A(net8568),
    .X(net8566));
 sky130_fd_sc_hd__clkbuf_2 max_length8567 (.A(net8568),
    .X(net8567));
 sky130_fd_sc_hd__buf_1 wire8568 (.A(net8564),
    .X(net8568));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout8569 (.A(net8575),
    .X(net8569));
 sky130_fd_sc_hd__buf_1 wire8570 (.A(net8572),
    .X(net8570));
 sky130_fd_sc_hd__clkbuf_1 max_length8571 (.A(net8572),
    .X(net8571));
 sky130_fd_sc_hd__clkbuf_2 wire8572 (.A(net8569),
    .X(net8572));
 sky130_fd_sc_hd__clkbuf_2 fanout8573 (.A(net8578),
    .X(net8573));
 sky130_fd_sc_hd__buf_1 wire8574 (.A(net8573),
    .X(net8574));
 sky130_fd_sc_hd__buf_1 fanout8575 (.A(net8592),
    .X(net8575));
 sky130_fd_sc_hd__clkbuf_1 wire8576 (.A(net8577),
    .X(net8576));
 sky130_fd_sc_hd__buf_1 max_length8577 (.A(net8578),
    .X(net8577));
 sky130_fd_sc_hd__buf_1 wire8578 (.A(net8580),
    .X(net8578));
 sky130_fd_sc_hd__buf_1 wire8579 (.A(net8580),
    .X(net8579));
 sky130_fd_sc_hd__clkbuf_2 max_length8580 (.A(net8575),
    .X(net8580));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout8581 (.A(net8585),
    .X(net8581));
 sky130_fd_sc_hd__buf_1 wire8582 (.A(net8583),
    .X(net8582));
 sky130_fd_sc_hd__buf_1 wire8583 (.A(net8584),
    .X(net8583));
 sky130_fd_sc_hd__clkbuf_2 max_length8584 (.A(net8581),
    .X(net8584));
 sky130_fd_sc_hd__clkbuf_1 fanout8585 (.A(net8593),
    .X(net8585));
 sky130_fd_sc_hd__buf_1 wire8586 (.A(net8587),
    .X(net8586));
 sky130_fd_sc_hd__buf_1 wire8587 (.A(net8588),
    .X(net8587));
 sky130_fd_sc_hd__buf_1 wire8588 (.A(net8589),
    .X(net8588));
 sky130_fd_sc_hd__buf_1 wire8589 (.A(net8585),
    .X(net8589));
 sky130_fd_sc_hd__buf_1 fanout8590 (.A(net8815),
    .X(net8590));
 sky130_fd_sc_hd__clkbuf_1 wire8591 (.A(net8592),
    .X(net8591));
 sky130_fd_sc_hd__buf_1 wire8592 (.A(net8593),
    .X(net8592));
 sky130_fd_sc_hd__buf_1 wire8593 (.A(net8594),
    .X(net8593));
 sky130_fd_sc_hd__buf_1 wire8594 (.A(net8595),
    .X(net8594));
 sky130_fd_sc_hd__clkbuf_1 wire8595 (.A(net8596),
    .X(net8595));
 sky130_fd_sc_hd__clkbuf_1 wire8596 (.A(net8597),
    .X(net8596));
 sky130_fd_sc_hd__clkbuf_1 wire8597 (.A(net8598),
    .X(net8597));
 sky130_fd_sc_hd__clkbuf_1 wire8598 (.A(net8599),
    .X(net8598));
 sky130_fd_sc_hd__clkbuf_1 wire8599 (.A(net8600),
    .X(net8599));
 sky130_fd_sc_hd__clkbuf_1 wire8600 (.A(net8601),
    .X(net8600));
 sky130_fd_sc_hd__buf_1 wire8601 (.A(net8590),
    .X(net8601));
 sky130_fd_sc_hd__buf_1 fanout8602 (.A(net8607),
    .X(net8602));
 sky130_fd_sc_hd__buf_1 wire8603 (.A(net8604),
    .X(net8603));
 sky130_fd_sc_hd__clkbuf_2 wire8604 (.A(net8602),
    .X(net8604));
 sky130_fd_sc_hd__clkbuf_2 fanout8605 (.A(net8821),
    .X(net8605));
 sky130_fd_sc_hd__clkbuf_1 wire8606 (.A(net8607),
    .X(net8606));
 sky130_fd_sc_hd__buf_1 max_length8607 (.A(net8605),
    .X(net8607));
 sky130_fd_sc_hd__clkbuf_2 fanout8608 (.A(net8639),
    .X(net8608));
 sky130_fd_sc_hd__buf_1 wire8609 (.A(net8608),
    .X(net8609));
 sky130_fd_sc_hd__clkbuf_1 wire8610 (.A(net8611),
    .X(net8610));
 sky130_fd_sc_hd__clkbuf_1 wire8611 (.A(net8612),
    .X(net8611));
 sky130_fd_sc_hd__clkbuf_1 wire8612 (.A(net8613),
    .X(net8612));
 sky130_fd_sc_hd__clkbuf_1 wire8613 (.A(net8614),
    .X(net8613));
 sky130_fd_sc_hd__buf_1 wire8614 (.A(net8608),
    .X(net8614));
 sky130_fd_sc_hd__buf_1 fanout8615 (.A(net8634),
    .X(net8615));
 sky130_fd_sc_hd__clkbuf_2 wire8616 (.A(net8615),
    .X(net8616));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout8617 (.A(net8622),
    .X(net8617));
 sky130_fd_sc_hd__buf_1 max_length8618 (.A(net8619),
    .X(net8618));
 sky130_fd_sc_hd__clkbuf_2 wire8619 (.A(net8617),
    .X(net8619));
 sky130_fd_sc_hd__clkbuf_2 fanout8620 (.A(net8644),
    .X(net8620));
 sky130_fd_sc_hd__buf_2 wire8621 (.A(net8620),
    .X(net8621));
 sky130_fd_sc_hd__clkbuf_2 fanout8622 (.A(net8643),
    .X(net8622));
 sky130_fd_sc_hd__clkbuf_1 fanout8623 (.A(net8629),
    .X(net8623));
 sky130_fd_sc_hd__buf_1 wire8624 (.A(net8625),
    .X(net8624));
 sky130_fd_sc_hd__clkbuf_2 wire8625 (.A(net8623),
    .X(net8625));
 sky130_fd_sc_hd__buf_1 wire8626 (.A(net8623),
    .X(net8626));
 sky130_fd_sc_hd__buf_1 fanout8627 (.A(net8629),
    .X(net8627));
 sky130_fd_sc_hd__buf_1 wire8628 (.A(net8627),
    .X(net8628));
 sky130_fd_sc_hd__buf_1 fanout8629 (.A(net8642),
    .X(net8629));
 sky130_fd_sc_hd__clkbuf_2 wire8630 (.A(net8632),
    .X(net8630));
 sky130_fd_sc_hd__buf_1 wire8631 (.A(net8632),
    .X(net8631));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8632 (.A(net8629),
    .X(net8632));
 sky130_fd_sc_hd__clkbuf_1 fanout8633 (.A(net8826),
    .X(net8633));
 sky130_fd_sc_hd__clkbuf_1 wire8634 (.A(net8635),
    .X(net8634));
 sky130_fd_sc_hd__clkbuf_1 wire8635 (.A(net8636),
    .X(net8635));
 sky130_fd_sc_hd__clkbuf_1 wire8636 (.A(net8637),
    .X(net8636));
 sky130_fd_sc_hd__clkbuf_1 wire8637 (.A(net8638),
    .X(net8637));
 sky130_fd_sc_hd__clkbuf_1 wire8638 (.A(net8639),
    .X(net8638));
 sky130_fd_sc_hd__buf_1 wire8639 (.A(net8640),
    .X(net8639));
 sky130_fd_sc_hd__clkbuf_1 wire8640 (.A(net8641),
    .X(net8640));
 sky130_fd_sc_hd__clkbuf_1 wire8641 (.A(net8644),
    .X(net8641));
 sky130_fd_sc_hd__clkbuf_1 wire8642 (.A(net8643),
    .X(net8642));
 sky130_fd_sc_hd__buf_1 wire8643 (.A(net8633),
    .X(net8643));
 sky130_fd_sc_hd__buf_1 max_length8644 (.A(net8633),
    .X(net8644));
 sky130_fd_sc_hd__buf_1 fanout8645 (.A(net8660),
    .X(net8645));
 sky130_fd_sc_hd__buf_1 wire8646 (.A(net8645),
    .X(net8646));
 sky130_fd_sc_hd__clkbuf_2 wire8647 (.A(net8648),
    .X(net8647));
 sky130_fd_sc_hd__buf_1 wire8648 (.A(net8645),
    .X(net8648));
 sky130_fd_sc_hd__buf_1 fanout8649 (.A(net8653),
    .X(net8649));
 sky130_fd_sc_hd__clkbuf_2 wire8650 (.A(net8649),
    .X(net8650));
 sky130_fd_sc_hd__buf_1 wire8651 (.A(net8652),
    .X(net8651));
 sky130_fd_sc_hd__buf_1 max_length8652 (.A(net8649),
    .X(net8652));
 sky130_fd_sc_hd__clkbuf_1 fanout8653 (.A(net8658),
    .X(net8653));
 sky130_fd_sc_hd__buf_1 max_length8654 (.A(net8655),
    .X(net8654));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8655 (.A(net8656),
    .X(net8655));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8656 (.A(net8657),
    .X(net8656));
 sky130_fd_sc_hd__buf_1 wire8657 (.A(net8653),
    .X(net8657));
 sky130_fd_sc_hd__clkbuf_1 fanout8658 (.A(net8706),
    .X(net8658));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8659 (.A(net8660),
    .X(net8659));
 sky130_fd_sc_hd__buf_1 wire8660 (.A(net8658),
    .X(net8660));
 sky130_fd_sc_hd__buf_1 fanout8661 (.A(net8664),
    .X(net8661));
 sky130_fd_sc_hd__clkbuf_2 wire8662 (.A(net8661),
    .X(net8662));
 sky130_fd_sc_hd__clkbuf_2 wire8663 (.A(net8661),
    .X(net8663));
 sky130_fd_sc_hd__buf_1 fanout8664 (.A(net8670),
    .X(net8664));
 sky130_fd_sc_hd__buf_1 max_length8665 (.A(net8667),
    .X(net8665));
 sky130_fd_sc_hd__buf_1 max_length8666 (.A(net8667),
    .X(net8666));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8667 (.A(net8668),
    .X(net8667));
 sky130_fd_sc_hd__buf_1 max_length8668 (.A(net8664),
    .X(net8668));
 sky130_fd_sc_hd__buf_1 fanout8669 (.A(net8703),
    .X(net8669));
 sky130_fd_sc_hd__buf_1 wire8670 (.A(net8669),
    .X(net8670));
 sky130_fd_sc_hd__buf_1 max_length8671 (.A(net8672),
    .X(net8671));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8672 (.A(net8669),
    .X(net8672));
 sky130_fd_sc_hd__clkbuf_2 fanout8673 (.A(net8697),
    .X(net8673));
 sky130_fd_sc_hd__buf_1 wire8674 (.A(net8675),
    .X(net8674));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8675 (.A(net8673),
    .X(net8675));
 sky130_fd_sc_hd__buf_1 max_length8676 (.A(net8673),
    .X(net8676));
 sky130_fd_sc_hd__buf_1 fanout8677 (.A(net8699),
    .X(net8677));
 sky130_fd_sc_hd__buf_1 max_length8678 (.A(net8679),
    .X(net8678));
 sky130_fd_sc_hd__buf_1 wire8679 (.A(net8677),
    .X(net8679));
 sky130_fd_sc_hd__buf_1 fanout8680 (.A(net8685),
    .X(net8680));
 sky130_fd_sc_hd__buf_1 max_length8681 (.A(net8682),
    .X(net8681));
 sky130_fd_sc_hd__buf_1 max_length8682 (.A(net8683),
    .X(net8682));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8683 (.A(net8680),
    .X(net8683));
 sky130_fd_sc_hd__clkbuf_2 fanout8684 (.A(net8701),
    .X(net8684));
 sky130_fd_sc_hd__buf_1 wire8685 (.A(net8684),
    .X(net8685));
 sky130_fd_sc_hd__buf_1 wire8686 (.A(net8684),
    .X(net8686));
 sky130_fd_sc_hd__buf_1 fanout8687 (.A(net8695),
    .X(net8687));
 sky130_fd_sc_hd__buf_1 wire8688 (.A(net8689),
    .X(net8688));
 sky130_fd_sc_hd__buf_1 wire8689 (.A(net8690),
    .X(net8689));
 sky130_fd_sc_hd__buf_1 max_length8690 (.A(net8691),
    .X(net8690));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8691 (.A(net8687),
    .X(net8691));
 sky130_fd_sc_hd__buf_1 fanout8692 (.A(net8698),
    .X(net8692));
 sky130_fd_sc_hd__buf_1 wire8693 (.A(net8694),
    .X(net8693));
 sky130_fd_sc_hd__clkbuf_2 wire8694 (.A(net8695),
    .X(net8694));
 sky130_fd_sc_hd__buf_1 wire8695 (.A(net8692),
    .X(net8695));
 sky130_fd_sc_hd__buf_1 fanout8696 (.A(net8702),
    .X(net8696));
 sky130_fd_sc_hd__clkbuf_1 wire8697 (.A(net8701),
    .X(net8697));
 sky130_fd_sc_hd__clkbuf_1 wire8698 (.A(net8700),
    .X(net8698));
 sky130_fd_sc_hd__clkbuf_1 max_length8699 (.A(net8700),
    .X(net8699));
 sky130_fd_sc_hd__buf_1 wire8700 (.A(net8696),
    .X(net8700));
 sky130_fd_sc_hd__buf_1 max_length8701 (.A(net8696),
    .X(net8701));
 sky130_fd_sc_hd__buf_1 fanout8702 (.A(net8731),
    .X(net8702));
 sky130_fd_sc_hd__buf_1 wire8703 (.A(net8704),
    .X(net8703));
 sky130_fd_sc_hd__clkbuf_1 wire8704 (.A(net8705),
    .X(net8704));
 sky130_fd_sc_hd__clkbuf_1 max_length8705 (.A(net8706),
    .X(net8705));
 sky130_fd_sc_hd__buf_1 wire8706 (.A(net8707),
    .X(net8706));
 sky130_fd_sc_hd__buf_1 wire8707 (.A(net8702),
    .X(net8707));
 sky130_fd_sc_hd__buf_1 fanout8708 (.A(net8713),
    .X(net8708));
 sky130_fd_sc_hd__buf_1 wire8709 (.A(net8710),
    .X(net8709));
 sky130_fd_sc_hd__clkbuf_2 max_length8710 (.A(net8711),
    .X(net8710));
 sky130_fd_sc_hd__clkbuf_2 max_length8711 (.A(net8708),
    .X(net8711));
 sky130_fd_sc_hd__buf_1 fanout8712 (.A(net8720),
    .X(net8712));
 sky130_fd_sc_hd__buf_1 wire8713 (.A(net8712),
    .X(net8713));
 sky130_fd_sc_hd__buf_1 wire8714 (.A(net8715),
    .X(net8714));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8715 (.A(net8716),
    .X(net8715));
 sky130_fd_sc_hd__buf_1 max_length8716 (.A(net8712),
    .X(net8716));
 sky130_fd_sc_hd__buf_1 fanout8717 (.A(net8722),
    .X(net8717));
 sky130_fd_sc_hd__buf_1 wire8718 (.A(net8719),
    .X(net8718));
 sky130_fd_sc_hd__clkbuf_1 wire8719 (.A(net8720),
    .X(net8719));
 sky130_fd_sc_hd__buf_1 max_length8720 (.A(net8721),
    .X(net8720));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8721 (.A(net8717),
    .X(net8721));
 sky130_fd_sc_hd__buf_1 fanout8722 (.A(net8732),
    .X(net8722));
 sky130_fd_sc_hd__clkbuf_2 wire8723 (.A(net8724),
    .X(net8723));
 sky130_fd_sc_hd__clkbuf_1 wire8724 (.A(net8725),
    .X(net8724));
 sky130_fd_sc_hd__clkbuf_1 wire8725 (.A(net8726),
    .X(net8725));
 sky130_fd_sc_hd__buf_1 wire8726 (.A(net8722),
    .X(net8726));
 sky130_fd_sc_hd__buf_1 fanout8727 (.A(net8733),
    .X(net8727));
 sky130_fd_sc_hd__clkbuf_2 wire8728 (.A(net8729),
    .X(net8728));
 sky130_fd_sc_hd__clkbuf_2 wire8729 (.A(net8727),
    .X(net8729));
 sky130_fd_sc_hd__buf_2 fanout8730 (.A(net8733),
    .X(net8730));
 sky130_fd_sc_hd__buf_1 fanout8731 (.A(net8827),
    .X(net8731));
 sky130_fd_sc_hd__buf_1 wire8732 (.A(net8738),
    .X(net8732));
 sky130_fd_sc_hd__buf_1 wire8733 (.A(net8734),
    .X(net8733));
 sky130_fd_sc_hd__clkbuf_1 wire8734 (.A(net8735),
    .X(net8734));
 sky130_fd_sc_hd__clkbuf_1 wire8735 (.A(net8736),
    .X(net8735));
 sky130_fd_sc_hd__clkbuf_1 wire8736 (.A(net8737),
    .X(net8736));
 sky130_fd_sc_hd__clkbuf_1 wire8737 (.A(net8738),
    .X(net8737));
 sky130_fd_sc_hd__buf_1 wire8738 (.A(net8739),
    .X(net8738));
 sky130_fd_sc_hd__clkbuf_1 wire8739 (.A(net8740),
    .X(net8739));
 sky130_fd_sc_hd__clkbuf_1 wire8740 (.A(net8741),
    .X(net8740));
 sky130_fd_sc_hd__clkbuf_1 wire8741 (.A(net8742),
    .X(net8741));
 sky130_fd_sc_hd__clkbuf_1 wire8742 (.A(net8731),
    .X(net8742));
 sky130_fd_sc_hd__buf_1 fanout8743 (.A(net8747),
    .X(net8743));
 sky130_fd_sc_hd__buf_1 wire8744 (.A(net8745),
    .X(net8744));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8745 (.A(net8743),
    .X(net8745));
 sky130_fd_sc_hd__buf_1 wire8746 (.A(net8743),
    .X(net8746));
 sky130_fd_sc_hd__clkbuf_2 fanout8747 (.A(net8751),
    .X(net8747));
 sky130_fd_sc_hd__buf_1 wire8748 (.A(net8750),
    .X(net8748));
 sky130_fd_sc_hd__clkbuf_1 max_length8749 (.A(net8750),
    .X(net8749));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8750 (.A(net8747),
    .X(net8750));
 sky130_fd_sc_hd__clkbuf_1 fanout8751 (.A(net8793),
    .X(net8751));
 sky130_fd_sc_hd__buf_1 max_length8752 (.A(net8753),
    .X(net8752));
 sky130_fd_sc_hd__buf_1 wire8753 (.A(net8755),
    .X(net8753));
 sky130_fd_sc_hd__buf_1 wire8754 (.A(net8755),
    .X(net8754));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8755 (.A(net8751),
    .X(net8755));
 sky130_fd_sc_hd__clkbuf_1 fanout8756 (.A(net8763),
    .X(net8756));
 sky130_fd_sc_hd__buf_1 wire8757 (.A(net8758),
    .X(net8757));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8758 (.A(net8759),
    .X(net8758));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8759 (.A(net8756),
    .X(net8759));
 sky130_fd_sc_hd__clkbuf_1 fanout8760 (.A(net8766),
    .X(net8760));
 sky130_fd_sc_hd__buf_1 max_length8761 (.A(net8762),
    .X(net8761));
 sky130_fd_sc_hd__clkbuf_2 wire8762 (.A(net8760),
    .X(net8762));
 sky130_fd_sc_hd__buf_1 fanout8763 (.A(net8798),
    .X(net8763));
 sky130_fd_sc_hd__buf_1 wire8764 (.A(net8765),
    .X(net8764));
 sky130_fd_sc_hd__buf_1 wire8765 (.A(net8763),
    .X(net8765));
 sky130_fd_sc_hd__clkbuf_1 max_length8766 (.A(net8763),
    .X(net8766));
 sky130_fd_sc_hd__buf_2 fanout8767 (.A(net8772),
    .X(net8767));
 sky130_fd_sc_hd__buf_1 wire8768 (.A(net8767),
    .X(net8768));
 sky130_fd_sc_hd__buf_1 fanout8769 (.A(net8796),
    .X(net8769));
 sky130_fd_sc_hd__buf_1 wire8770 (.A(net8771),
    .X(net8770));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8771 (.A(net8772),
    .X(net8771));
 sky130_fd_sc_hd__buf_1 wire8772 (.A(net8769),
    .X(net8772));
 sky130_fd_sc_hd__buf_1 fanout8773 (.A(net8800),
    .X(net8773));
 sky130_fd_sc_hd__clkbuf_1 wire8774 (.A(net8775),
    .X(net8774));
 sky130_fd_sc_hd__buf_1 max_length8775 (.A(net8776),
    .X(net8775));
 sky130_fd_sc_hd__buf_1 wire8776 (.A(net8777),
    .X(net8776));
 sky130_fd_sc_hd__clkbuf_2 wire8777 (.A(net8773),
    .X(net8777));
 sky130_fd_sc_hd__buf_1 fanout8778 (.A(net8799),
    .X(net8778));
 sky130_fd_sc_hd__buf_1 wire8779 (.A(net8780),
    .X(net8779));
 sky130_fd_sc_hd__buf_1 wire8780 (.A(net8778),
    .X(net8780));
 sky130_fd_sc_hd__buf_2 fanout8781 (.A(net8790),
    .X(net8781));
 sky130_fd_sc_hd__buf_1 wire8782 (.A(net8781),
    .X(net8782));
 sky130_fd_sc_hd__buf_1 wire8783 (.A(net8781),
    .X(net8783));
 sky130_fd_sc_hd__buf_1 fanout8784 (.A(net8790),
    .X(net8784));
 sky130_fd_sc_hd__clkbuf_2 wire8785 (.A(net8784),
    .X(net8785));
 sky130_fd_sc_hd__buf_1 fanout8786 (.A(net8791),
    .X(net8786));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8787 (.A(net8788),
    .X(net8787));
 sky130_fd_sc_hd__buf_1 wire8788 (.A(net8789),
    .X(net8788));
 sky130_fd_sc_hd__buf_1 wire8789 (.A(net8786),
    .X(net8789));
 sky130_fd_sc_hd__buf_1 fanout8790 (.A(net8801),
    .X(net8790));
 sky130_fd_sc_hd__buf_1 wire8791 (.A(net8790),
    .X(net8791));
 sky130_fd_sc_hd__buf_1 fanout8792 (.A(net8839),
    .X(net8792));
 sky130_fd_sc_hd__clkbuf_1 wire8793 (.A(net8794),
    .X(net8793));
 sky130_fd_sc_hd__clkbuf_1 wire8794 (.A(net8795),
    .X(net8794));
 sky130_fd_sc_hd__clkbuf_1 wire8795 (.A(net8796),
    .X(net8795));
 sky130_fd_sc_hd__buf_1 wire8796 (.A(net8792),
    .X(net8796));
 sky130_fd_sc_hd__buf_1 wire8797 (.A(net8798),
    .X(net8797));
 sky130_fd_sc_hd__buf_1 wire8798 (.A(net8800),
    .X(net8798));
 sky130_fd_sc_hd__clkbuf_1 max_length8799 (.A(net8800),
    .X(net8799));
 sky130_fd_sc_hd__buf_1 wire8800 (.A(net8801),
    .X(net8800));
 sky130_fd_sc_hd__buf_1 wire8801 (.A(net8802),
    .X(net8801));
 sky130_fd_sc_hd__clkbuf_1 wire8802 (.A(net8792),
    .X(net8802));
 sky130_fd_sc_hd__clkbuf_2 fanout8803 (.A(net8808),
    .X(net8803));
 sky130_fd_sc_hd__clkbuf_1 wire8804 (.A(net8805),
    .X(net8804));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8805 (.A(net8803),
    .X(net8805));
 sky130_fd_sc_hd__buf_1 max_length8806 (.A(net8803),
    .X(net8806));
 sky130_fd_sc_hd__clkbuf_2 fanout8807 (.A(net8812),
    .X(net8807));
 sky130_fd_sc_hd__buf_1 fanout8808 (.A(net8834),
    .X(net8808));
 sky130_fd_sc_hd__buf_1 wire8809 (.A(net8810),
    .X(net8809));
 sky130_fd_sc_hd__buf_1 max_length8810 (.A(net8811),
    .X(net8810));
 sky130_fd_sc_hd__buf_1 wire8811 (.A(net8808),
    .X(net8811));
 sky130_fd_sc_hd__clkbuf_1 wire8812 (.A(net8813),
    .X(net8812));
 sky130_fd_sc_hd__clkbuf_1 max_length8813 (.A(net8808),
    .X(net8813));
 sky130_fd_sc_hd__buf_1 fanout8814 (.A(net8856),
    .X(net8814));
 sky130_fd_sc_hd__clkbuf_1 wire8815 (.A(net8816),
    .X(net8815));
 sky130_fd_sc_hd__clkbuf_1 wire8816 (.A(net8817),
    .X(net8816));
 sky130_fd_sc_hd__clkbuf_1 wire8817 (.A(net8818),
    .X(net8817));
 sky130_fd_sc_hd__clkbuf_1 wire8818 (.A(net8819),
    .X(net8818));
 sky130_fd_sc_hd__clkbuf_1 wire8819 (.A(net8820),
    .X(net8819));
 sky130_fd_sc_hd__clkbuf_1 wire8820 (.A(net8821),
    .X(net8820));
 sky130_fd_sc_hd__buf_1 wire8821 (.A(net8822),
    .X(net8821));
 sky130_fd_sc_hd__buf_1 wire8822 (.A(net8823),
    .X(net8822));
 sky130_fd_sc_hd__clkbuf_1 wire8823 (.A(net8824),
    .X(net8823));
 sky130_fd_sc_hd__clkbuf_1 wire8824 (.A(net8825),
    .X(net8824));
 sky130_fd_sc_hd__clkbuf_1 wire8825 (.A(net8826),
    .X(net8825));
 sky130_fd_sc_hd__buf_1 wire8826 (.A(net8814),
    .X(net8826));
 sky130_fd_sc_hd__clkbuf_1 wire8827 (.A(net8828),
    .X(net8827));
 sky130_fd_sc_hd__clkbuf_1 wire8828 (.A(net8829),
    .X(net8828));
 sky130_fd_sc_hd__clkbuf_1 wire8829 (.A(net8830),
    .X(net8829));
 sky130_fd_sc_hd__clkbuf_1 wire8830 (.A(net8831),
    .X(net8830));
 sky130_fd_sc_hd__clkbuf_1 wire8831 (.A(net8839),
    .X(net8831));
 sky130_fd_sc_hd__clkbuf_1 wire8832 (.A(net8833),
    .X(net8832));
 sky130_fd_sc_hd__clkbuf_1 wire8833 (.A(net8834),
    .X(net8833));
 sky130_fd_sc_hd__buf_1 wire8834 (.A(net8835),
    .X(net8834));
 sky130_fd_sc_hd__clkbuf_1 wire8835 (.A(net8836),
    .X(net8835));
 sky130_fd_sc_hd__clkbuf_1 wire8836 (.A(net8837),
    .X(net8836));
 sky130_fd_sc_hd__clkbuf_1 wire8837 (.A(net8838),
    .X(net8837));
 sky130_fd_sc_hd__clkbuf_1 wire8838 (.A(net8839),
    .X(net8838));
 sky130_fd_sc_hd__buf_1 wire8839 (.A(net8840),
    .X(net8839));
 sky130_fd_sc_hd__clkbuf_1 wire8840 (.A(net8841),
    .X(net8840));
 sky130_fd_sc_hd__clkbuf_1 wire8841 (.A(net8842),
    .X(net8841));
 sky130_fd_sc_hd__clkbuf_1 wire8842 (.A(net8843),
    .X(net8842));
 sky130_fd_sc_hd__clkbuf_1 wire8843 (.A(net8814),
    .X(net8843));
 sky130_fd_sc_hd__clkbuf_1 wire8844 (.A(net8845),
    .X(net8844));
 sky130_fd_sc_hd__clkbuf_1 wire8845 (.A(net8846),
    .X(net8845));
 sky130_fd_sc_hd__clkbuf_1 wire8846 (.A(net8847),
    .X(net8846));
 sky130_fd_sc_hd__clkbuf_1 wire8847 (.A(net8848),
    .X(net8847));
 sky130_fd_sc_hd__clkbuf_1 wire8848 (.A(net8849),
    .X(net8848));
 sky130_fd_sc_hd__clkbuf_1 wire8849 (.A(net8850),
    .X(net8849));
 sky130_fd_sc_hd__clkbuf_1 wire8850 (.A(net8851),
    .X(net8850));
 sky130_fd_sc_hd__clkbuf_1 wire8851 (.A(net8852),
    .X(net8851));
 sky130_fd_sc_hd__clkbuf_1 wire8852 (.A(net8853),
    .X(net8852));
 sky130_fd_sc_hd__clkbuf_1 wire8853 (.A(net8854),
    .X(net8853));
 sky130_fd_sc_hd__clkbuf_1 wire8854 (.A(net8855),
    .X(net8854));
 sky130_fd_sc_hd__clkbuf_1 max_length8855 (.A(net8856),
    .X(net8855));
 sky130_fd_sc_hd__buf_1 wire8856 (.A(net8857),
    .X(net8856));
 sky130_fd_sc_hd__clkbuf_1 wire8857 (.A(net8858),
    .X(net8857));
 sky130_fd_sc_hd__clkbuf_1 wire8858 (.A(net8859),
    .X(net8858));
 sky130_fd_sc_hd__clkbuf_1 wire8859 (.A(net8860),
    .X(net8859));
 sky130_fd_sc_hd__clkbuf_1 wire8860 (.A(net8861),
    .X(net8860));
 sky130_fd_sc_hd__clkbuf_1 wire8861 (.A(net147),
    .X(net8861));
 sky130_fd_sc_hd__clkbuf_1 fanout8862 (.A(net8874),
    .X(net8862));
 sky130_fd_sc_hd__buf_1 wire8863 (.A(net8865),
    .X(net8863));
 sky130_fd_sc_hd__buf_1 wire8864 (.A(net8865),
    .X(net8864));
 sky130_fd_sc_hd__buf_1 wire8865 (.A(net8862),
    .X(net8865));
 sky130_fd_sc_hd__buf_1 fanout8866 (.A(net8870),
    .X(net8866));
 sky130_fd_sc_hd__buf_1 wire8867 (.A(net8868),
    .X(net8867));
 sky130_fd_sc_hd__buf_1 wire8868 (.A(net8866),
    .X(net8868));
 sky130_fd_sc_hd__buf_1 fanout8869 (.A(net8873),
    .X(net8869));
 sky130_fd_sc_hd__buf_1 wire8870 (.A(net8871),
    .X(net8870));
 sky130_fd_sc_hd__buf_1 max_length8871 (.A(net8872),
    .X(net8871));
 sky130_fd_sc_hd__clkbuf_1 wire8872 (.A(net8869),
    .X(net8872));
 sky130_fd_sc_hd__clkbuf_1 fanout8873 (.A(net146),
    .X(net8873));
 sky130_fd_sc_hd__buf_1 wire8874 (.A(net8876),
    .X(net8874));
 sky130_fd_sc_hd__clkbuf_1 max_length8875 (.A(net8876),
    .X(net8875));
 sky130_fd_sc_hd__buf_1 wire8876 (.A(net8877),
    .X(net8876));
 sky130_fd_sc_hd__clkbuf_1 wire8877 (.A(net8878),
    .X(net8877));
 sky130_fd_sc_hd__clkbuf_1 wire8878 (.A(net8879),
    .X(net8878));
 sky130_fd_sc_hd__clkbuf_1 wire8879 (.A(net8880),
    .X(net8879));
 sky130_fd_sc_hd__clkbuf_1 wire8880 (.A(net8873),
    .X(net8880));
 sky130_fd_sc_hd__clkbuf_1 wire8881 (.A(net134),
    .X(net8881));
 sky130_fd_sc_hd__clkbuf_1 wire8882 (.A(net8883),
    .X(net8882));
 sky130_fd_sc_hd__clkbuf_1 wire8883 (.A(net8884),
    .X(net8883));
 sky130_fd_sc_hd__clkbuf_1 wire8884 (.A(net131),
    .X(net8884));
 sky130_fd_sc_hd__clkbuf_1 wire8885 (.A(net128),
    .X(net8885));
 sky130_fd_sc_hd__clkbuf_1 wire8886 (.A(net127),
    .X(net8886));
 sky130_fd_sc_hd__buf_1 fanout8887 (.A(net8890),
    .X(net8887));
 sky130_fd_sc_hd__buf_1 max_length8888 (.A(net8889),
    .X(net8888));
 sky130_fd_sc_hd__buf_1 wire8889 (.A(net8887),
    .X(net8889));
 sky130_fd_sc_hd__buf_1 fanout8890 (.A(net8900),
    .X(net8890));
 sky130_fd_sc_hd__buf_1 wire8891 (.A(net8892),
    .X(net8891));
 sky130_fd_sc_hd__buf_1 wire8892 (.A(net8894),
    .X(net8892));
 sky130_fd_sc_hd__buf_1 wire8893 (.A(net8894),
    .X(net8893));
 sky130_fd_sc_hd__buf_1 wire8894 (.A(net8890),
    .X(net8894));
 sky130_fd_sc_hd__buf_1 fanout8895 (.A(net8899),
    .X(net8895));
 sky130_fd_sc_hd__clkbuf_1 max_length8896 (.A(net8897),
    .X(net8896));
 sky130_fd_sc_hd__clkbuf_2 wire8897 (.A(net8898),
    .X(net8897));
 sky130_fd_sc_hd__buf_1 wire8898 (.A(net8895),
    .X(net8898));
 sky130_fd_sc_hd__buf_1 fanout8899 (.A(net8907),
    .X(net8899));
 sky130_fd_sc_hd__clkbuf_1 max_length8900 (.A(net8901),
    .X(net8900));
 sky130_fd_sc_hd__buf_1 wire8901 (.A(net8902),
    .X(net8901));
 sky130_fd_sc_hd__buf_1 wire8902 (.A(net8903),
    .X(net8902));
 sky130_fd_sc_hd__buf_1 wire8903 (.A(net8899),
    .X(net8903));
 sky130_fd_sc_hd__buf_1 fanout8904 (.A(net8911),
    .X(net8904));
 sky130_fd_sc_hd__buf_1 wire8905 (.A(net8906),
    .X(net8905));
 sky130_fd_sc_hd__buf_1 wire8906 (.A(net8904),
    .X(net8906));
 sky130_fd_sc_hd__buf_1 wire8907 (.A(net8908),
    .X(net8907));
 sky130_fd_sc_hd__clkbuf_1 wire8908 (.A(net8904),
    .X(net8908));
 sky130_fd_sc_hd__clkbuf_1 wire8909 (.A(net8915),
    .X(net8909));
 sky130_fd_sc_hd__clkbuf_1 wire8910 (.A(net8911),
    .X(net8910));
 sky130_fd_sc_hd__buf_1 wire8911 (.A(net8912),
    .X(net8911));
 sky130_fd_sc_hd__clkbuf_1 wire8912 (.A(net8913),
    .X(net8912));
 sky130_fd_sc_hd__clkbuf_1 wire8913 (.A(net8914),
    .X(net8913));
 sky130_fd_sc_hd__clkbuf_1 wire8914 (.A(net8916),
    .X(net8914));
 sky130_fd_sc_hd__clkbuf_1 max_length8915 (.A(net8916),
    .X(net8915));
 sky130_fd_sc_hd__buf_1 wire8916 (.A(net8917),
    .X(net8916));
 sky130_fd_sc_hd__clkbuf_1 wire8917 (.A(net8918),
    .X(net8917));
 sky130_fd_sc_hd__clkbuf_1 wire8918 (.A(net8919),
    .X(net8918));
 sky130_fd_sc_hd__clkbuf_1 wire8919 (.A(net8920),
    .X(net8919));
 sky130_fd_sc_hd__clkbuf_1 wire8920 (.A(net8921),
    .X(net8920));
 sky130_fd_sc_hd__buf_1 wire8921 (.A(net8922),
    .X(net8921));
 sky130_fd_sc_hd__clkbuf_1 wire8922 (.A(net8923),
    .X(net8922));
 sky130_fd_sc_hd__clkbuf_1 wire8923 (.A(net113),
    .X(net8923));
 sky130_fd_sc_hd__clkbuf_1 wire8924 (.A(net8925),
    .X(net8924));
 sky130_fd_sc_hd__clkbuf_1 wire8925 (.A(net8926),
    .X(net8925));
 sky130_fd_sc_hd__clkbuf_1 wire8926 (.A(net8927),
    .X(net8926));
 sky130_fd_sc_hd__clkbuf_1 wire8927 (.A(net112),
    .X(net8927));
 sky130_fd_sc_hd__clkbuf_1 wire8928 (.A(net8929),
    .X(net8928));
 sky130_fd_sc_hd__clkbuf_1 wire8929 (.A(net8930),
    .X(net8929));
 sky130_fd_sc_hd__clkbuf_1 wire8930 (.A(net8931),
    .X(net8930));
 sky130_fd_sc_hd__clkbuf_1 wire8931 (.A(net111),
    .X(net8931));
 sky130_fd_sc_hd__clkbuf_1 wire8932 (.A(net8933),
    .X(net8932));
 sky130_fd_sc_hd__clkbuf_1 wire8933 (.A(net8934),
    .X(net8933));
 sky130_fd_sc_hd__clkbuf_1 wire8934 (.A(net8935),
    .X(net8934));
 sky130_fd_sc_hd__clkbuf_1 wire8935 (.A(net103),
    .X(net8935));
 sky130_fd_sc_hd__clkbuf_1 wire8936 (.A(net8937),
    .X(net8936));
 sky130_fd_sc_hd__clkbuf_1 wire8937 (.A(net8938),
    .X(net8937));
 sky130_fd_sc_hd__clkbuf_1 wire8938 (.A(net8939),
    .X(net8938));
 sky130_fd_sc_hd__clkbuf_1 wire8939 (.A(net102),
    .X(net8939));
 sky130_fd_sc_hd__clkbuf_1 wire8940 (.A(net8941),
    .X(net8940));
 sky130_fd_sc_hd__clkbuf_1 wire8941 (.A(net8942),
    .X(net8941));
 sky130_fd_sc_hd__clkbuf_1 wire8942 (.A(net8943),
    .X(net8942));
 sky130_fd_sc_hd__clkbuf_1 wire8943 (.A(net8944),
    .X(net8943));
 sky130_fd_sc_hd__clkbuf_1 wire8944 (.A(net8945),
    .X(net8944));
 sky130_fd_sc_hd__clkbuf_1 wire8945 (.A(net101),
    .X(net8945));
 sky130_fd_sc_hd__clkbuf_1 wire8946 (.A(net8947),
    .X(net8946));
 sky130_fd_sc_hd__clkbuf_1 wire8947 (.A(net8948),
    .X(net8947));
 sky130_fd_sc_hd__clkbuf_1 wire8948 (.A(net8949),
    .X(net8948));
 sky130_fd_sc_hd__clkbuf_1 wire8949 (.A(net8950),
    .X(net8949));
 sky130_fd_sc_hd__clkbuf_1 wire8950 (.A(net8951),
    .X(net8950));
 sky130_fd_sc_hd__clkbuf_1 wire8951 (.A(net8952),
    .X(net8951));
 sky130_fd_sc_hd__clkbuf_1 wire8952 (.A(net100),
    .X(net8952));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire8953 (.A(net1),
    .X(net8953));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_8__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_10__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_11__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_12__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_15__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\matmul0.matmul_stage_inst.c[9] ),
    .X(net8954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\matmul0.matmul_stage_inst.c[6] ),
    .X(net8955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\matmul0.matmul_stage_inst.a[10] ),
    .X(net8956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\pid_d.curr_error[5] ),
    .X(net8957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\matmul0.matmul_stage_inst.a[7] ),
    .X(net8958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\matmul0.matmul_stage_inst.a[2] ),
    .X(net8959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\matmul0.matmul_stage_inst.a[0] ),
    .X(net8960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\matmul0.matmul_stage_inst.a[5] ),
    .X(net8961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net150),
    .X(net8962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_00408_),
    .X(net8963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\svm0.vC[9] ),
    .X(net8964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\matmul0.matmul_stage_inst.a[9] ),
    .X(net8965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\cordic0.sin[3] ),
    .X(net8966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\svm0.vC[11] ),
    .X(net8967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\cordic0.cos[3] ),
    .X(net8968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\matmul0.matmul_stage_inst.a[4] ),
    .X(net8969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\matmul0.matmul_stage_inst.a[8] ),
    .X(net8970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\svm0.tA[9] ),
    .X(net8971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\cordic0.cos[9] ),
    .X(net8972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\matmul0.matmul_stage_inst.b[15] ),
    .X(net8973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\matmul0.matmul_stage_inst.c[5] ),
    .X(net8974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\cordic0.cos[6] ),
    .X(net8975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\matmul0.matmul_stage_inst.start ),
    .X(net8976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_00014_),
    .X(net8977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\matmul0.matmul_stage_inst.d[10] ),
    .X(net8978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\matmul0.matmul_stage_inst.a[1] ),
    .X(net8979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\matmul0.matmul_stage_inst.b[0] ),
    .X(net8980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\matmul0.matmul_stage_inst.a[3] ),
    .X(net8981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\matmul0.matmul_stage_inst.a[12] ),
    .X(net8982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\pid_q.curr_error[13] ),
    .X(net8983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\matmul0.matmul_stage_inst.a[14] ),
    .X(net8984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\pid_q.target[3] ),
    .X(net8985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\pid_q.target[1] ),
    .X(net8986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\pid_d.curr_error[0] ),
    .X(net8987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\pid_d.prev_error[14] ),
    .X(net8988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\matmul0.matmul_stage_inst.a[6] ),
    .X(net8989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\pid_q.target[14] ),
    .X(net8990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\matmul0.matmul_stage_inst.b[13] ),
    .X(net8991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\pid_d.iterate_enable ),
    .X(net8992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\pid_d.curr_error[13] ),
    .X(net8993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\matmul0.matmul_stage_inst.b[5] ),
    .X(net8994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\svm0.vC[13] ),
    .X(net8995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\pid_q.curr_int[2] ),
    .X(net8996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\cordic0.cos[5] ),
    .X(net8997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\cordic0.out_valid ),
    .X(net8998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\pid_q.target[9] ),
    .X(net8999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net151),
    .X(net9000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_00407_),
    .X(net9001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\matmul0.matmul_stage_inst.d[6] ),
    .X(net9002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\matmul0.matmul_stage_inst.c[10] ),
    .X(net9003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\pid_q.target[4] ),
    .X(net9004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\svm0.vC[6] ),
    .X(net9005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\cordic0.cos[10] ),
    .X(net9006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\matmul0.matmul_stage_inst.d[0] ),
    .X(net9007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\matmul0.matmul_stage_inst.d[7] ),
    .X(net9008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\pid_d.curr_int[1] ),
    .X(net9009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\pid_q.target[0] ),
    .X(net9010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\pid_q.target[11] ),
    .X(net9011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\pid_d.prev_error[12] ),
    .X(net9012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\pid_d.curr_error[9] ),
    .X(net9013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\pid_q.target[5] ),
    .X(net9014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\pid_q.curr_int[15] ),
    .X(net9015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\cordic0.sin[5] ),
    .X(net9016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\matmul0.matmul_stage_inst.c[4] ),
    .X(net9017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\pid_d.curr_int[9] ),
    .X(net9018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\matmul0.matmul_stage_inst.d[4] ),
    .X(net9019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\matmul0.matmul_stage_inst.d[5] ),
    .X(net9020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\matmul0.matmul_stage_inst.a[11] ),
    .X(net9021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\pid_d.curr_int[7] ),
    .X(net9022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\pid_q.target[2] ),
    .X(net9023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\matmul0.matmul_stage_inst.a[13] ),
    .X(net9024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\cordic0.cos[8] ),
    .X(net9025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\matmul0.matmul_stage_inst.d[12] ),
    .X(net9026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\cordic0.sin[1] ),
    .X(net9027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\pid_d.curr_error[3] ),
    .X(net9028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\cordic0.cos[1] ),
    .X(net9029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\svm0.vC[8] ),
    .X(net9030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\matmul0.matmul_stage_inst.b[4] ),
    .X(net9031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\pid_q.prev_error[12] ),
    .X(net9032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\matmul0.matmul_stage_inst.b[3] ),
    .X(net9033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\matmul0.matmul_stage_inst.c[8] ),
    .X(net9034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\pid_d.curr_int[8] ),
    .X(net9035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\matmul0.matmul_stage_inst.b[6] ),
    .X(net9036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\pid_d.curr_error[1] ),
    .X(net9037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\cordic0.cos[7] ),
    .X(net9038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\matmul0.matmul_stage_inst.b[9] ),
    .X(net9039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\matmul0.matmul_stage_inst.c[11] ),
    .X(net9040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\svm0.counter[15] ),
    .X(net9041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\pid_q.target[13] ),
    .X(net9042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\pid_d.curr_error[11] ),
    .X(net9043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\matmul0.matmul_stage_inst.d[11] ),
    .X(net9044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\matmul0.matmul_stage_inst.d[8] ),
    .X(net9045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\cordic0.cos[12] ),
    .X(net9046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\svm0.vC[4] ),
    .X(net9047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net149),
    .X(net9048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\cordic0.cos[0] ),
    .X(net9049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\pid_d.curr_error[2] ),
    .X(net9050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\svm0.vC[3] ),
    .X(net9051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\matmul0.matmul_stage_inst.d[1] ),
    .X(net9052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\pid_q.target[6] ),
    .X(net9053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\svm0.tB[1] ),
    .X(net9054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\pid_q.curr_error[1] ),
    .X(net9055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\svm0.vC[10] ),
    .X(net9056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\matmul0.matmul_stage_inst.c[15] ),
    .X(net9057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\svm0.vC[5] ),
    .X(net9058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\cordic0.sin[0] ),
    .X(net9059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\pid_q.target[7] ),
    .X(net9060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\pid_d.curr_error[15] ),
    .X(net9061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\cordic0.sin[10] ),
    .X(net9062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\matmul0.matmul_stage_inst.c[3] ),
    .X(net9063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\cordic0.sin[6] ),
    .X(net9064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\matmul0.matmul_stage_inst.d[9] ),
    .X(net9065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\pid_q.curr_int[13] ),
    .X(net9066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\pid_q.prev_error[14] ),
    .X(net9067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\svm0.vC[7] ),
    .X(net9068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\matmul0.matmul_stage_inst.d[2] ),
    .X(net9069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\svm0.vC[1] ),
    .X(net9070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\matmul0.matmul_stage_inst.c[1] ),
    .X(net9071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\svm0.vC[0] ),
    .X(net9072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\cordic0.sin[13] ),
    .X(net9073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\cordic0.sin[11] ),
    .X(net9074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\cordic0.sin[4] ),
    .X(net9075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\cordic0.sin[9] ),
    .X(net9076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\pid_q.curr_int[11] ),
    .X(net9077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\pid_q.target[10] ),
    .X(net9078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\pid_d.curr_int[2] ),
    .X(net9079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\svm0.tB[9] ),
    .X(net9080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\matmul0.matmul_stage_inst.b[1] ),
    .X(net9081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\matmul0.matmul_stage_inst.b[10] ),
    .X(net9082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\pid_d.prev_error[15] ),
    .X(net9083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\svm0.vC[14] ),
    .X(net9084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\cordic0.sin[8] ),
    .X(net9085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\matmul0.op_in[1] ),
    .X(net9086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\matmul0.matmul_stage_inst.d[13] ),
    .X(net9087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\cordic0.sin[2] ),
    .X(net9088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\svm0.tA[0] ),
    .X(net9089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\svm0.tB[6] ),
    .X(net9090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\svm0.tC[14] ),
    .X(net9091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\matmul0.matmul_stage_inst.b[12] ),
    .X(net9092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\svm0.tA[6] ),
    .X(net9093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\matmul0.matmul_stage_inst.b[7] ),
    .X(net9094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\svm0.vC[2] ),
    .X(net9095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\svm0.tB[14] ),
    .X(net9096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\svm0.vC[15] ),
    .X(net9097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\cordic0.sin[7] ),
    .X(net9098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\svm0.tB[8] ),
    .X(net9099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\svm0.tA[8] ),
    .X(net9100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\cordic0.sin[12] ),
    .X(net9101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\cordic0.in_valid ),
    .X(net9102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\pid_q.target[8] ),
    .X(net9103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\matmul0.matmul_stage_inst.c[2] ),
    .X(net9104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\pid_d.prev_error[9] ),
    .X(net9105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\pid_d.prev_error[3] ),
    .X(net9106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\pid_q.prev_error[15] ),
    .X(net9107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\svm0.tA[1] ),
    .X(net9108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\pid_d.prev_int[13] ),
    .X(net9109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\svm0.in_valid ),
    .X(net9110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\svm0.tA[14] ),
    .X(net9111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\svm0.tC[9] ),
    .X(net9112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\matmul0.matmul_stage_inst.b[8] ),
    .X(net9113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\pid_d.prev_error[7] ),
    .X(net9114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\svm0.vC[12] ),
    .X(net9115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\matmul0.matmul_stage_inst.c[12] ),
    .X(net9116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\pid_d.prev_error[6] ),
    .X(net9117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\svm0.tC[6] ),
    .X(net9118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\pid_d.prev_error[8] ),
    .X(net9119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\matmul0.matmul_stage_inst.b[14] ),
    .X(net9120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\pid_d.prev_error[10] ),
    .X(net9121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\pid_q.prev_int[15] ),
    .X(net9122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\pid_q.prev_error[7] ),
    .X(net9123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\pid_d.prev_error[5] ),
    .X(net9124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\pid_q.prev_int[13] ),
    .X(net9125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\svm0.tC[12] ),
    .X(net9126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\pid_q.prev_error[10] ),
    .X(net9127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\matmul0.matmul_stage_inst.c[7] ),
    .X(net9128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\svm0.tB[13] ),
    .X(net9129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\matmul0.matmul_stage_inst.b[11] ),
    .X(net9130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\svm0.tA[13] ),
    .X(net9131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\svm0.tB[5] ),
    .X(net9132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\pid_q.prev_error[9] ),
    .X(net9133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\pid_d.prev_int[15] ),
    .X(net9134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\pid_d.prev_error[2] ),
    .X(net9135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\svm0.tA[5] ),
    .X(net9136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\svm0.tC[4] ),
    .X(net9137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\pid_d.prev_error[4] ),
    .X(net9138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\pid_q.prev_error[4] ),
    .X(net9139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\svm0.tB[4] ),
    .X(net9140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\svm0.tB[12] ),
    .X(net9141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\pid_q.prev_error[8] ),
    .X(net9142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\svm0.tA[12] ),
    .X(net9143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\pid_q.prev_error[5] ),
    .X(net9144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\pid_q.prev_error[6] ),
    .X(net9145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\matmul0.matmul_stage_inst.c[14] ),
    .X(net9146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\svm0.tC[3] ),
    .X(net9147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\matmul0.matmul_stage_inst.state[0] ),
    .X(net9148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\svm0.tC[2] ),
    .X(net9149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\matmul0.state[0] ),
    .X(net9150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\pid_q.curr_error[14] ),
    .X(net9151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\svm0.tC[0] ),
    .X(net9152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\cordic0.slte0.opA[16] ),
    .X(net9153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\pid_d.mult0.b[8] ),
    .X(net9154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\svm0.tB[0] ),
    .X(net9155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\pid_d.mult0.b[11] ),
    .X(net9156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\svm0.tC[13] ),
    .X(net9157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\matmul0.a_in[3] ),
    .X(net9158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\pid_d.prev_error[13] ),
    .X(net9159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\cordic0.slte0.opA[1] ),
    .X(net9160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\svm0.tC[8] ),
    .X(net9161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\svm0.delta[13] ),
    .X(net9162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\pid_q.out[0] ),
    .X(net9163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\pid_q.curr_error[15] ),
    .X(net9164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\svm0.tB[10] ),
    .X(net9165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\pid_q.out[5] ),
    .X(net9166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\svm0.tB[3] ),
    .X(net9167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\cordic0.slte0.opA[5] ),
    .X(net9168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\pid_d.curr_int[10] ),
    .X(net9169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_00803_),
    .X(net9170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\pid_d.mult0.b[9] ),
    .X(net9171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\svm0.tA[10] ),
    .X(net9172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\pid_q.out[8] ),
    .X(net9173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\pid_q.out[6] ),
    .X(net9174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\pid_q.prev_error[3] ),
    .X(net9175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\svm0.tB[11] ),
    .X(net9176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\pid_q.prev_error[0] ),
    .X(net9177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\pid_q.prev_error[2] ),
    .X(net9178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\pid_q.prev_error[13] ),
    .X(net9179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\svm0.tC[5] ),
    .X(net9180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\pid_d.prev_error[11] ),
    .X(net9181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\pid_d.prev_error[1] ),
    .X(net9182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\matmul0.a[13] ),
    .X(net9183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\pid_q.prev_error[11] ),
    .X(net9184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\pid_q.prev_int[12] ),
    .X(net9185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\svm0.tA[4] ),
    .X(net9186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\cordic0.slte0.opA[2] ),
    .X(net9187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\cordic0.slte0.opA[8] ),
    .X(net9188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\pid_q.prev_int[14] ),
    .X(net9189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\svm0.tA[15] ),
    .X(net9190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\cordic0.slte0.opA[14] ),
    .X(net9191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\matmul0.op_in[0] ),
    .X(net9192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\pid_q.curr_error[10] ),
    .X(net9193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\svm0.tC[15] ),
    .X(net9194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\pid_d.curr_int[15] ),
    .X(net9195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\pid_d.curr_int[6] ),
    .X(net9196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_00799_),
    .X(net9197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\svm0.tC[10] ),
    .X(net9198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\svm0.calc_ready ),
    .X(net9199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\pid_q.prev_int[8] ),
    .X(net9200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\pid_q.prev_int[11] ),
    .X(net9201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\pid_q.curr_int[10] ),
    .X(net9202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_00424_),
    .X(net9203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\svm0.tB[2] ),
    .X(net9204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\pid_d.prev_int[9] ),
    .X(net9205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\pid_d.curr_int[0] ),
    .X(net9206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\pid_q.prev_int[3] ),
    .X(net9207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\cordic0.slte0.opA[0] ),
    .X(net9208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\pid_d.prev_int[4] ),
    .X(net9209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\cordic0.cos[11] ),
    .X(net9210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\pid_q.prev_int[6] ),
    .X(net9211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\pid_q.prev_int[5] ),
    .X(net9212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\svm0.delta[15] ),
    .X(net9213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\svm0.tB[15] ),
    .X(net9214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\pid_d.prev_int[7] ),
    .X(net9215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\cordic0.slte0.opA[17] ),
    .X(net9216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\pid_d.prev_int[8] ),
    .X(net9217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\cordic0.slte0.opA[4] ),
    .X(net9218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\svm0.tB[7] ),
    .X(net9219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\svm0.tA[7] ),
    .X(net9220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\pid_q.prev_int[7] ),
    .X(net9221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\svm0.tC[11] ),
    .X(net9222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\pid_q.prev_int[9] ),
    .X(net9223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\pid_d.prev_int[11] ),
    .X(net9224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\matmul0.b[11] ),
    .X(net9225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\matmul0.b_in[4] ),
    .X(net9226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\matmul0.a[9] ),
    .X(net9227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\pid_q.prev_error[1] ),
    .X(net9228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\pid_q.out[7] ),
    .X(net9229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\matmul0.b[12] ),
    .X(net9230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\matmul0.a[4] ),
    .X(net9231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\svm0.tA[11] ),
    .X(net9232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\cordic0.cos[13] ),
    .X(net9233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\pid_d.ki[7] ),
    .X(net9234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\matmul0.beta_pass[13] ),
    .X(net9235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\pid_d.prev_int[5] ),
    .X(net9236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\matmul0.b[13] ),
    .X(net9237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\matmul0.beta_pass[5] ),
    .X(net9238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\pid_q.prev_int[4] ),
    .X(net9239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\cordic0.cos[1] ),
    .X(net9240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\cordic0.cos[5] ),
    .X(net9241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\matmul0.b[11] ),
    .X(net9242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\pid_d.curr_int[6] ),
    .X(net9243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\svm0.calc_ready ),
    .X(net9244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\cordic0.sin[6] ),
    .X(net9245));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net3152));
 sky130_fd_sc_hd__clkbuf_1 max_cap1 (.A(net9247),
    .X(net9246));
 sky130_fd_sc_hd__clkbuf_1 wire2 (.A(_08877_),
    .X(net9247));
 sky130_fd_sc_hd__buf_1 max_cap3 (.A(_02716_),
    .X(net9248));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_954 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1095 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1010 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1066 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1092 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1008 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1094 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_870 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_983 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1087 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1098 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_898 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1095 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1157 ();
endmodule
