module fpga_wrapper (clk_mosi,
    clk_sys,
    cs,
    pwmA,
    pwmB,
    pwmC,
    ready,
    rstb,
    spi_mosi);
 input clk_mosi;
 input clk_sys;
 input cs;
 output pwmA;
 output pwmB;
 output pwmC;
 output ready;
 input rstb;
 input spi_mosi;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire \spi0.cs_sync[0] ;
 wire \spi0.cs_sync[1] ;
 wire \spi0.cs_sync[2] ;
 wire \spi0.data_packed[0] ;
 wire \spi0.data_packed[10] ;
 wire \spi0.data_packed[11] ;
 wire \spi0.data_packed[12] ;
 wire \spi0.data_packed[13] ;
 wire \spi0.data_packed[14] ;
 wire \spi0.data_packed[15] ;
 wire \spi0.data_packed[16] ;
 wire \spi0.data_packed[17] ;
 wire \spi0.data_packed[18] ;
 wire \spi0.data_packed[19] ;
 wire \spi0.data_packed[1] ;
 wire \spi0.data_packed[20] ;
 wire \spi0.data_packed[21] ;
 wire \spi0.data_packed[22] ;
 wire \spi0.data_packed[23] ;
 wire \spi0.data_packed[24] ;
 wire \spi0.data_packed[25] ;
 wire \spi0.data_packed[26] ;
 wire \spi0.data_packed[27] ;
 wire \spi0.data_packed[28] ;
 wire \spi0.data_packed[29] ;
 wire \spi0.data_packed[2] ;
 wire \spi0.data_packed[30] ;
 wire \spi0.data_packed[31] ;
 wire \spi0.data_packed[32] ;
 wire \spi0.data_packed[33] ;
 wire \spi0.data_packed[34] ;
 wire \spi0.data_packed[35] ;
 wire \spi0.data_packed[36] ;
 wire \spi0.data_packed[37] ;
 wire \spi0.data_packed[38] ;
 wire \spi0.data_packed[39] ;
 wire \spi0.data_packed[3] ;
 wire \spi0.data_packed[40] ;
 wire \spi0.data_packed[41] ;
 wire \spi0.data_packed[42] ;
 wire \spi0.data_packed[43] ;
 wire \spi0.data_packed[44] ;
 wire \spi0.data_packed[45] ;
 wire \spi0.data_packed[46] ;
 wire \spi0.data_packed[47] ;
 wire \spi0.data_packed[48] ;
 wire \spi0.data_packed[49] ;
 wire \spi0.data_packed[4] ;
 wire \spi0.data_packed[50] ;
 wire \spi0.data_packed[51] ;
 wire \spi0.data_packed[52] ;
 wire \spi0.data_packed[53] ;
 wire \spi0.data_packed[54] ;
 wire \spi0.data_packed[55] ;
 wire \spi0.data_packed[56] ;
 wire \spi0.data_packed[57] ;
 wire \spi0.data_packed[58] ;
 wire \spi0.data_packed[59] ;
 wire \spi0.data_packed[5] ;
 wire \spi0.data_packed[60] ;
 wire \spi0.data_packed[61] ;
 wire \spi0.data_packed[62] ;
 wire \spi0.data_packed[63] ;
 wire \spi0.data_packed[64] ;
 wire \spi0.data_packed[65] ;
 wire \spi0.data_packed[66] ;
 wire \spi0.data_packed[67] ;
 wire \spi0.data_packed[68] ;
 wire \spi0.data_packed[69] ;
 wire \spi0.data_packed[6] ;
 wire \spi0.data_packed[70] ;
 wire \spi0.data_packed[71] ;
 wire \spi0.data_packed[72] ;
 wire \spi0.data_packed[73] ;
 wire \spi0.data_packed[74] ;
 wire \spi0.data_packed[75] ;
 wire \spi0.data_packed[76] ;
 wire \spi0.data_packed[77] ;
 wire \spi0.data_packed[78] ;
 wire \spi0.data_packed[79] ;
 wire \spi0.data_packed[7] ;
 wire \spi0.data_packed[8] ;
 wire \spi0.data_packed[9] ;
 wire \spi0.opcode[0] ;
 wire \spi0.opcode[1] ;
 wire \spi0.opcode[2] ;
 wire \spi0.opcode[3] ;
 wire \spi0.opcode[4] ;
 wire \spi0.opcode[5] ;
 wire \spi0.opcode[6] ;
 wire \spi0.opcode[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \top0.a_in_matmul[0] ;
 wire \top0.a_in_matmul[10] ;
 wire \top0.a_in_matmul[11] ;
 wire \top0.a_in_matmul[12] ;
 wire \top0.a_in_matmul[13] ;
 wire \top0.a_in_matmul[14] ;
 wire \top0.a_in_matmul[15] ;
 wire \top0.a_in_matmul[1] ;
 wire \top0.a_in_matmul[2] ;
 wire \top0.a_in_matmul[3] ;
 wire \top0.a_in_matmul[4] ;
 wire \top0.a_in_matmul[5] ;
 wire \top0.a_in_matmul[6] ;
 wire \top0.a_in_matmul[7] ;
 wire \top0.a_in_matmul[8] ;
 wire \top0.a_in_matmul[9] ;
 wire \top0.b_in_matmul[0] ;
 wire \top0.b_in_matmul[10] ;
 wire \top0.b_in_matmul[11] ;
 wire \top0.b_in_matmul[12] ;
 wire \top0.b_in_matmul[13] ;
 wire \top0.b_in_matmul[14] ;
 wire \top0.b_in_matmul[15] ;
 wire \top0.b_in_matmul[1] ;
 wire \top0.b_in_matmul[2] ;
 wire \top0.b_in_matmul[3] ;
 wire \top0.b_in_matmul[4] ;
 wire \top0.b_in_matmul[5] ;
 wire \top0.b_in_matmul[6] ;
 wire \top0.b_in_matmul[7] ;
 wire \top0.b_in_matmul[8] ;
 wire \top0.b_in_matmul[9] ;
 wire \top0.c_out_calc[0] ;
 wire \top0.c_out_calc[10] ;
 wire \top0.c_out_calc[11] ;
 wire \top0.c_out_calc[12] ;
 wire \top0.c_out_calc[13] ;
 wire \top0.c_out_calc[14] ;
 wire \top0.c_out_calc[15] ;
 wire \top0.c_out_calc[1] ;
 wire \top0.c_out_calc[2] ;
 wire \top0.c_out_calc[3] ;
 wire \top0.c_out_calc[4] ;
 wire \top0.c_out_calc[5] ;
 wire \top0.c_out_calc[6] ;
 wire \top0.c_out_calc[7] ;
 wire \top0.c_out_calc[8] ;
 wire \top0.c_out_calc[9] ;
 wire \top0.clarke_done ;
 wire \top0.cordic0.cos[0] ;
 wire \top0.cordic0.cos[10] ;
 wire \top0.cordic0.cos[11] ;
 wire \top0.cordic0.cos[12] ;
 wire \top0.cordic0.cos[13] ;
 wire \top0.cordic0.cos[1] ;
 wire \top0.cordic0.cos[2] ;
 wire \top0.cordic0.cos[3] ;
 wire \top0.cordic0.cos[4] ;
 wire \top0.cordic0.cos[5] ;
 wire \top0.cordic0.cos[6] ;
 wire \top0.cordic0.cos[7] ;
 wire \top0.cordic0.cos[8] ;
 wire \top0.cordic0.cos[9] ;
 wire \top0.cordic0.domain[0] ;
 wire \top0.cordic0.domain[1] ;
 wire \top0.cordic0.gm0.iter[0] ;
 wire \top0.cordic0.gm0.iter[1] ;
 wire \top0.cordic0.gm0.iter[2] ;
 wire \top0.cordic0.gm0.iter[3] ;
 wire \top0.cordic0.gm0.iter[4] ;
 wire \top0.cordic0.in_valid ;
 wire \top0.cordic0.out_valid ;
 wire \top0.cordic0.sin[0] ;
 wire \top0.cordic0.sin[10] ;
 wire \top0.cordic0.sin[11] ;
 wire \top0.cordic0.sin[12] ;
 wire \top0.cordic0.sin[13] ;
 wire \top0.cordic0.sin[1] ;
 wire \top0.cordic0.sin[2] ;
 wire \top0.cordic0.sin[3] ;
 wire \top0.cordic0.sin[4] ;
 wire \top0.cordic0.sin[5] ;
 wire \top0.cordic0.sin[6] ;
 wire \top0.cordic0.sin[7] ;
 wire \top0.cordic0.sin[8] ;
 wire \top0.cordic0.sin[9] ;
 wire \top0.cordic0.slte0.opA[0] ;
 wire \top0.cordic0.slte0.opA[10] ;
 wire \top0.cordic0.slte0.opA[11] ;
 wire \top0.cordic0.slte0.opA[12] ;
 wire \top0.cordic0.slte0.opA[13] ;
 wire \top0.cordic0.slte0.opA[14] ;
 wire \top0.cordic0.slte0.opA[15] ;
 wire \top0.cordic0.slte0.opA[16] ;
 wire \top0.cordic0.slte0.opA[17] ;
 wire \top0.cordic0.slte0.opA[1] ;
 wire \top0.cordic0.slte0.opA[2] ;
 wire \top0.cordic0.slte0.opA[3] ;
 wire \top0.cordic0.slte0.opA[4] ;
 wire \top0.cordic0.slte0.opA[5] ;
 wire \top0.cordic0.slte0.opA[6] ;
 wire \top0.cordic0.slte0.opA[7] ;
 wire \top0.cordic0.slte0.opA[8] ;
 wire \top0.cordic0.slte0.opA[9] ;
 wire \top0.cordic0.slte0.opB[10] ;
 wire \top0.cordic0.slte0.opB[11] ;
 wire \top0.cordic0.slte0.opB[12] ;
 wire \top0.cordic0.slte0.opB[13] ;
 wire \top0.cordic0.slte0.opB[14] ;
 wire \top0.cordic0.slte0.opB[15] ;
 wire \top0.cordic0.slte0.opB[2] ;
 wire \top0.cordic0.slte0.opB[3] ;
 wire \top0.cordic0.slte0.opB[4] ;
 wire \top0.cordic0.slte0.opB[5] ;
 wire \top0.cordic0.slte0.opB[6] ;
 wire \top0.cordic0.slte0.opB[7] ;
 wire \top0.cordic0.slte0.opB[8] ;
 wire \top0.cordic0.slte0.opB[9] ;
 wire \top0.cordic0.state[0] ;
 wire \top0.cordic0.vec[0][0] ;
 wire \top0.cordic0.vec[0][10] ;
 wire \top0.cordic0.vec[0][11] ;
 wire \top0.cordic0.vec[0][12] ;
 wire \top0.cordic0.vec[0][13] ;
 wire \top0.cordic0.vec[0][14] ;
 wire \top0.cordic0.vec[0][15] ;
 wire \top0.cordic0.vec[0][16] ;
 wire \top0.cordic0.vec[0][17] ;
 wire \top0.cordic0.vec[0][1] ;
 wire \top0.cordic0.vec[0][2] ;
 wire \top0.cordic0.vec[0][3] ;
 wire \top0.cordic0.vec[0][4] ;
 wire \top0.cordic0.vec[0][5] ;
 wire \top0.cordic0.vec[0][6] ;
 wire \top0.cordic0.vec[0][7] ;
 wire \top0.cordic0.vec[0][8] ;
 wire \top0.cordic0.vec[0][9] ;
 wire \top0.cordic0.vec[1][0] ;
 wire \top0.cordic0.vec[1][10] ;
 wire \top0.cordic0.vec[1][11] ;
 wire \top0.cordic0.vec[1][12] ;
 wire \top0.cordic0.vec[1][13] ;
 wire \top0.cordic0.vec[1][14] ;
 wire \top0.cordic0.vec[1][15] ;
 wire \top0.cordic0.vec[1][16] ;
 wire \top0.cordic0.vec[1][17] ;
 wire \top0.cordic0.vec[1][1] ;
 wire \top0.cordic0.vec[1][2] ;
 wire \top0.cordic0.vec[1][3] ;
 wire \top0.cordic0.vec[1][4] ;
 wire \top0.cordic0.vec[1][5] ;
 wire \top0.cordic0.vec[1][6] ;
 wire \top0.cordic0.vec[1][7] ;
 wire \top0.cordic0.vec[1][8] ;
 wire \top0.cordic0.vec[1][9] ;
 wire \top0.cordic_done ;
 wire \top0.currT_r[0] ;
 wire \top0.currT_r[10] ;
 wire \top0.currT_r[11] ;
 wire \top0.currT_r[12] ;
 wire \top0.currT_r[13] ;
 wire \top0.currT_r[14] ;
 wire \top0.currT_r[15] ;
 wire \top0.currT_r[1] ;
 wire \top0.currT_r[2] ;
 wire \top0.currT_r[3] ;
 wire \top0.currT_r[4] ;
 wire \top0.currT_r[5] ;
 wire \top0.currT_r[6] ;
 wire \top0.currT_r[7] ;
 wire \top0.currT_r[8] ;
 wire \top0.currT_r[9] ;
 wire \top0.kid[0] ;
 wire \top0.kid[10] ;
 wire \top0.kid[11] ;
 wire \top0.kid[12] ;
 wire \top0.kid[13] ;
 wire \top0.kid[14] ;
 wire \top0.kid[15] ;
 wire \top0.kid[1] ;
 wire \top0.kid[2] ;
 wire \top0.kid[3] ;
 wire \top0.kid[4] ;
 wire \top0.kid[5] ;
 wire \top0.kid[6] ;
 wire \top0.kid[7] ;
 wire \top0.kid[8] ;
 wire \top0.kid[9] ;
 wire \top0.kiq[0] ;
 wire \top0.kiq[10] ;
 wire \top0.kiq[11] ;
 wire \top0.kiq[12] ;
 wire \top0.kiq[13] ;
 wire \top0.kiq[14] ;
 wire \top0.kiq[15] ;
 wire \top0.kiq[1] ;
 wire \top0.kiq[2] ;
 wire \top0.kiq[3] ;
 wire \top0.kiq[4] ;
 wire \top0.kiq[5] ;
 wire \top0.kiq[6] ;
 wire \top0.kiq[7] ;
 wire \top0.kiq[8] ;
 wire \top0.kiq[9] ;
 wire \top0.kpd[0] ;
 wire \top0.kpd[10] ;
 wire \top0.kpd[11] ;
 wire \top0.kpd[12] ;
 wire \top0.kpd[13] ;
 wire \top0.kpd[14] ;
 wire \top0.kpd[15] ;
 wire \top0.kpd[1] ;
 wire \top0.kpd[2] ;
 wire \top0.kpd[3] ;
 wire \top0.kpd[4] ;
 wire \top0.kpd[5] ;
 wire \top0.kpd[6] ;
 wire \top0.kpd[7] ;
 wire \top0.kpd[8] ;
 wire \top0.kpd[9] ;
 wire \top0.kpq[0] ;
 wire \top0.kpq[10] ;
 wire \top0.kpq[11] ;
 wire \top0.kpq[12] ;
 wire \top0.kpq[13] ;
 wire \top0.kpq[14] ;
 wire \top0.kpq[15] ;
 wire \top0.kpq[1] ;
 wire \top0.kpq[2] ;
 wire \top0.kpq[3] ;
 wire \top0.kpq[4] ;
 wire \top0.kpq[5] ;
 wire \top0.kpq[6] ;
 wire \top0.kpq[7] ;
 wire \top0.kpq[8] ;
 wire \top0.kpq[9] ;
 wire \top0.matmul0.a[0] ;
 wire \top0.matmul0.a[10] ;
 wire \top0.matmul0.a[11] ;
 wire \top0.matmul0.a[12] ;
 wire \top0.matmul0.a[13] ;
 wire \top0.matmul0.a[14] ;
 wire \top0.matmul0.a[15] ;
 wire \top0.matmul0.a[1] ;
 wire \top0.matmul0.a[2] ;
 wire \top0.matmul0.a[3] ;
 wire \top0.matmul0.a[4] ;
 wire \top0.matmul0.a[5] ;
 wire \top0.matmul0.a[6] ;
 wire \top0.matmul0.a[7] ;
 wire \top0.matmul0.a[8] ;
 wire \top0.matmul0.a[9] ;
 wire \top0.matmul0.alpha_pass[0] ;
 wire \top0.matmul0.alpha_pass[10] ;
 wire \top0.matmul0.alpha_pass[11] ;
 wire \top0.matmul0.alpha_pass[12] ;
 wire \top0.matmul0.alpha_pass[13] ;
 wire \top0.matmul0.alpha_pass[14] ;
 wire \top0.matmul0.alpha_pass[15] ;
 wire \top0.matmul0.alpha_pass[1] ;
 wire \top0.matmul0.alpha_pass[2] ;
 wire \top0.matmul0.alpha_pass[3] ;
 wire \top0.matmul0.alpha_pass[4] ;
 wire \top0.matmul0.alpha_pass[5] ;
 wire \top0.matmul0.alpha_pass[6] ;
 wire \top0.matmul0.alpha_pass[7] ;
 wire \top0.matmul0.alpha_pass[8] ;
 wire \top0.matmul0.alpha_pass[9] ;
 wire \top0.matmul0.b[0] ;
 wire \top0.matmul0.b[10] ;
 wire \top0.matmul0.b[11] ;
 wire \top0.matmul0.b[12] ;
 wire \top0.matmul0.b[13] ;
 wire \top0.matmul0.b[14] ;
 wire \top0.matmul0.b[15] ;
 wire \top0.matmul0.b[1] ;
 wire \top0.matmul0.b[2] ;
 wire \top0.matmul0.b[3] ;
 wire \top0.matmul0.b[4] ;
 wire \top0.matmul0.b[5] ;
 wire \top0.matmul0.b[6] ;
 wire \top0.matmul0.b[7] ;
 wire \top0.matmul0.b[8] ;
 wire \top0.matmul0.b[9] ;
 wire \top0.matmul0.beta_pass[0] ;
 wire \top0.matmul0.beta_pass[10] ;
 wire \top0.matmul0.beta_pass[11] ;
 wire \top0.matmul0.beta_pass[12] ;
 wire \top0.matmul0.beta_pass[13] ;
 wire \top0.matmul0.beta_pass[14] ;
 wire \top0.matmul0.beta_pass[15] ;
 wire \top0.matmul0.beta_pass[1] ;
 wire \top0.matmul0.beta_pass[2] ;
 wire \top0.matmul0.beta_pass[3] ;
 wire \top0.matmul0.beta_pass[4] ;
 wire \top0.matmul0.beta_pass[5] ;
 wire \top0.matmul0.beta_pass[6] ;
 wire \top0.matmul0.beta_pass[7] ;
 wire \top0.matmul0.beta_pass[8] ;
 wire \top0.matmul0.beta_pass[9] ;
 wire \top0.matmul0.cos[0] ;
 wire \top0.matmul0.cos[10] ;
 wire \top0.matmul0.cos[11] ;
 wire \top0.matmul0.cos[12] ;
 wire \top0.matmul0.cos[13] ;
 wire \top0.matmul0.cos[1] ;
 wire \top0.matmul0.cos[2] ;
 wire \top0.matmul0.cos[3] ;
 wire \top0.matmul0.cos[4] ;
 wire \top0.matmul0.cos[5] ;
 wire \top0.matmul0.cos[6] ;
 wire \top0.matmul0.cos[7] ;
 wire \top0.matmul0.cos[8] ;
 wire \top0.matmul0.cos[9] ;
 wire \top0.matmul0.done_pass ;
 wire \top0.matmul0.matmul_stage_inst.a[0] ;
 wire \top0.matmul0.matmul_stage_inst.a[10] ;
 wire \top0.matmul0.matmul_stage_inst.a[11] ;
 wire \top0.matmul0.matmul_stage_inst.a[12] ;
 wire \top0.matmul0.matmul_stage_inst.a[13] ;
 wire \top0.matmul0.matmul_stage_inst.a[14] ;
 wire \top0.matmul0.matmul_stage_inst.a[1] ;
 wire \top0.matmul0.matmul_stage_inst.a[2] ;
 wire \top0.matmul0.matmul_stage_inst.a[3] ;
 wire \top0.matmul0.matmul_stage_inst.a[4] ;
 wire \top0.matmul0.matmul_stage_inst.a[5] ;
 wire \top0.matmul0.matmul_stage_inst.a[6] ;
 wire \top0.matmul0.matmul_stage_inst.a[7] ;
 wire \top0.matmul0.matmul_stage_inst.a[8] ;
 wire \top0.matmul0.matmul_stage_inst.a[9] ;
 wire \top0.matmul0.matmul_stage_inst.b[0] ;
 wire \top0.matmul0.matmul_stage_inst.b[10] ;
 wire \top0.matmul0.matmul_stage_inst.b[11] ;
 wire \top0.matmul0.matmul_stage_inst.b[12] ;
 wire \top0.matmul0.matmul_stage_inst.b[13] ;
 wire \top0.matmul0.matmul_stage_inst.b[14] ;
 wire \top0.matmul0.matmul_stage_inst.b[15] ;
 wire \top0.matmul0.matmul_stage_inst.b[1] ;
 wire \top0.matmul0.matmul_stage_inst.b[2] ;
 wire \top0.matmul0.matmul_stage_inst.b[3] ;
 wire \top0.matmul0.matmul_stage_inst.b[4] ;
 wire \top0.matmul0.matmul_stage_inst.b[5] ;
 wire \top0.matmul0.matmul_stage_inst.b[6] ;
 wire \top0.matmul0.matmul_stage_inst.b[7] ;
 wire \top0.matmul0.matmul_stage_inst.b[8] ;
 wire \top0.matmul0.matmul_stage_inst.b[9] ;
 wire \top0.matmul0.matmul_stage_inst.c[10] ;
 wire \top0.matmul0.matmul_stage_inst.c[11] ;
 wire \top0.matmul0.matmul_stage_inst.c[12] ;
 wire \top0.matmul0.matmul_stage_inst.c[13] ;
 wire \top0.matmul0.matmul_stage_inst.c[14] ;
 wire \top0.matmul0.matmul_stage_inst.c[15] ;
 wire \top0.matmul0.matmul_stage_inst.c[1] ;
 wire \top0.matmul0.matmul_stage_inst.c[2] ;
 wire \top0.matmul0.matmul_stage_inst.c[3] ;
 wire \top0.matmul0.matmul_stage_inst.c[4] ;
 wire \top0.matmul0.matmul_stage_inst.c[5] ;
 wire \top0.matmul0.matmul_stage_inst.c[6] ;
 wire \top0.matmul0.matmul_stage_inst.c[7] ;
 wire \top0.matmul0.matmul_stage_inst.c[8] ;
 wire \top0.matmul0.matmul_stage_inst.c[9] ;
 wire \top0.matmul0.matmul_stage_inst.d[0] ;
 wire \top0.matmul0.matmul_stage_inst.d[10] ;
 wire \top0.matmul0.matmul_stage_inst.d[11] ;
 wire \top0.matmul0.matmul_stage_inst.d[12] ;
 wire \top0.matmul0.matmul_stage_inst.d[13] ;
 wire \top0.matmul0.matmul_stage_inst.d[1] ;
 wire \top0.matmul0.matmul_stage_inst.d[2] ;
 wire \top0.matmul0.matmul_stage_inst.d[4] ;
 wire \top0.matmul0.matmul_stage_inst.d[5] ;
 wire \top0.matmul0.matmul_stage_inst.d[6] ;
 wire \top0.matmul0.matmul_stage_inst.d[7] ;
 wire \top0.matmul0.matmul_stage_inst.d[8] ;
 wire \top0.matmul0.matmul_stage_inst.d[9] ;
 wire \top0.matmul0.matmul_stage_inst.e[0] ;
 wire \top0.matmul0.matmul_stage_inst.e[10] ;
 wire \top0.matmul0.matmul_stage_inst.e[11] ;
 wire \top0.matmul0.matmul_stage_inst.e[12] ;
 wire \top0.matmul0.matmul_stage_inst.e[13] ;
 wire \top0.matmul0.matmul_stage_inst.e[14] ;
 wire \top0.matmul0.matmul_stage_inst.e[15] ;
 wire \top0.matmul0.matmul_stage_inst.e[1] ;
 wire \top0.matmul0.matmul_stage_inst.e[2] ;
 wire \top0.matmul0.matmul_stage_inst.e[3] ;
 wire \top0.matmul0.matmul_stage_inst.e[4] ;
 wire \top0.matmul0.matmul_stage_inst.e[5] ;
 wire \top0.matmul0.matmul_stage_inst.e[6] ;
 wire \top0.matmul0.matmul_stage_inst.e[7] ;
 wire \top0.matmul0.matmul_stage_inst.e[8] ;
 wire \top0.matmul0.matmul_stage_inst.e[9] ;
 wire \top0.matmul0.matmul_stage_inst.f[0] ;
 wire \top0.matmul0.matmul_stage_inst.f[10] ;
 wire \top0.matmul0.matmul_stage_inst.f[11] ;
 wire \top0.matmul0.matmul_stage_inst.f[12] ;
 wire \top0.matmul0.matmul_stage_inst.f[13] ;
 wire \top0.matmul0.matmul_stage_inst.f[14] ;
 wire \top0.matmul0.matmul_stage_inst.f[15] ;
 wire \top0.matmul0.matmul_stage_inst.f[1] ;
 wire \top0.matmul0.matmul_stage_inst.f[2] ;
 wire \top0.matmul0.matmul_stage_inst.f[3] ;
 wire \top0.matmul0.matmul_stage_inst.f[4] ;
 wire \top0.matmul0.matmul_stage_inst.f[5] ;
 wire \top0.matmul0.matmul_stage_inst.f[6] ;
 wire \top0.matmul0.matmul_stage_inst.f[7] ;
 wire \top0.matmul0.matmul_stage_inst.f[8] ;
 wire \top0.matmul0.matmul_stage_inst.f[9] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[0] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[10] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[11] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[12] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[13] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[14] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[15] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[1] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[2] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[3] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[4] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[5] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[6] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[7] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[8] ;
 wire \top0.matmul0.matmul_stage_inst.mult1[9] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[0] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[10] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[11] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[12] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[13] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[14] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[15] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[1] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[2] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[3] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[4] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[5] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[6] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[7] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[8] ;
 wire \top0.matmul0.matmul_stage_inst.mult2[9] ;
 wire \top0.matmul0.matmul_stage_inst.start ;
 wire \top0.matmul0.matmul_stage_inst.state[0] ;
 wire \top0.matmul0.matmul_stage_inst.state[1] ;
 wire \top0.matmul0.matmul_stage_inst.state[2] ;
 wire \top0.matmul0.matmul_stage_inst.state[4] ;
 wire \top0.matmul0.matmul_stage_inst.state[5] ;
 wire \top0.matmul0.matmul_stage_inst.state[6] ;
 wire \top0.matmul0.op[0] ;
 wire \top0.matmul0.op[1] ;
 wire \top0.matmul0.op_in[0] ;
 wire \top0.matmul0.op_in[1] ;
 wire \top0.matmul0.sin[0] ;
 wire \top0.matmul0.sin[10] ;
 wire \top0.matmul0.sin[11] ;
 wire \top0.matmul0.sin[12] ;
 wire \top0.matmul0.sin[13] ;
 wire \top0.matmul0.sin[1] ;
 wire \top0.matmul0.sin[2] ;
 wire \top0.matmul0.sin[3] ;
 wire \top0.matmul0.sin[4] ;
 wire \top0.matmul0.sin[5] ;
 wire \top0.matmul0.sin[6] ;
 wire \top0.matmul0.sin[7] ;
 wire \top0.matmul0.sin[8] ;
 wire \top0.matmul0.sin[9] ;
 wire \top0.matmul0.start ;
 wire \top0.matmul0.state[0] ;
 wire \top0.matmul0.state[1] ;
 wire \top0.periodTop[0] ;
 wire \top0.periodTop[10] ;
 wire \top0.periodTop[11] ;
 wire \top0.periodTop[12] ;
 wire \top0.periodTop[13] ;
 wire \top0.periodTop[14] ;
 wire \top0.periodTop[15] ;
 wire \top0.periodTop[1] ;
 wire \top0.periodTop[2] ;
 wire \top0.periodTop[3] ;
 wire \top0.periodTop[4] ;
 wire \top0.periodTop[5] ;
 wire \top0.periodTop[6] ;
 wire \top0.periodTop[7] ;
 wire \top0.periodTop[8] ;
 wire \top0.periodTop[9] ;
 wire \top0.periodTop_r[0] ;
 wire \top0.periodTop_r[10] ;
 wire \top0.periodTop_r[11] ;
 wire \top0.periodTop_r[12] ;
 wire \top0.periodTop_r[13] ;
 wire \top0.periodTop_r[14] ;
 wire \top0.periodTop_r[15] ;
 wire \top0.periodTop_r[1] ;
 wire \top0.periodTop_r[2] ;
 wire \top0.periodTop_r[3] ;
 wire \top0.periodTop_r[4] ;
 wire \top0.periodTop_r[5] ;
 wire \top0.periodTop_r[6] ;
 wire \top0.periodTop_r[7] ;
 wire \top0.periodTop_r[8] ;
 wire \top0.periodTop_r[9] ;
 wire \top0.pid_d.curr_error[0] ;
 wire \top0.pid_d.curr_error[10] ;
 wire \top0.pid_d.curr_error[11] ;
 wire \top0.pid_d.curr_error[12] ;
 wire \top0.pid_d.curr_error[13] ;
 wire \top0.pid_d.curr_error[14] ;
 wire \top0.pid_d.curr_error[15] ;
 wire \top0.pid_d.curr_error[1] ;
 wire \top0.pid_d.curr_error[2] ;
 wire \top0.pid_d.curr_error[3] ;
 wire \top0.pid_d.curr_error[4] ;
 wire \top0.pid_d.curr_error[5] ;
 wire \top0.pid_d.curr_error[6] ;
 wire \top0.pid_d.curr_error[7] ;
 wire \top0.pid_d.curr_error[8] ;
 wire \top0.pid_d.curr_error[9] ;
 wire \top0.pid_d.curr_int[0] ;
 wire \top0.pid_d.curr_int[10] ;
 wire \top0.pid_d.curr_int[11] ;
 wire \top0.pid_d.curr_int[12] ;
 wire \top0.pid_d.curr_int[13] ;
 wire \top0.pid_d.curr_int[14] ;
 wire \top0.pid_d.curr_int[15] ;
 wire \top0.pid_d.curr_int[1] ;
 wire \top0.pid_d.curr_int[2] ;
 wire \top0.pid_d.curr_int[3] ;
 wire \top0.pid_d.curr_int[4] ;
 wire \top0.pid_d.curr_int[5] ;
 wire \top0.pid_d.curr_int[6] ;
 wire \top0.pid_d.curr_int[7] ;
 wire \top0.pid_d.curr_int[8] ;
 wire \top0.pid_d.curr_int[9] ;
 wire \top0.pid_d.iterate_enable ;
 wire \top0.pid_d.mult0.a[0] ;
 wire \top0.pid_d.mult0.a[10] ;
 wire \top0.pid_d.mult0.a[11] ;
 wire \top0.pid_d.mult0.a[12] ;
 wire \top0.pid_d.mult0.a[13] ;
 wire \top0.pid_d.mult0.a[14] ;
 wire \top0.pid_d.mult0.a[15] ;
 wire \top0.pid_d.mult0.a[1] ;
 wire \top0.pid_d.mult0.a[2] ;
 wire \top0.pid_d.mult0.a[3] ;
 wire \top0.pid_d.mult0.a[4] ;
 wire \top0.pid_d.mult0.a[5] ;
 wire \top0.pid_d.mult0.a[6] ;
 wire \top0.pid_d.mult0.a[7] ;
 wire \top0.pid_d.mult0.a[8] ;
 wire \top0.pid_d.mult0.a[9] ;
 wire \top0.pid_d.mult0.b[0] ;
 wire \top0.pid_d.mult0.b[10] ;
 wire \top0.pid_d.mult0.b[11] ;
 wire \top0.pid_d.mult0.b[12] ;
 wire \top0.pid_d.mult0.b[13] ;
 wire \top0.pid_d.mult0.b[14] ;
 wire \top0.pid_d.mult0.b[15] ;
 wire \top0.pid_d.mult0.b[1] ;
 wire \top0.pid_d.mult0.b[2] ;
 wire \top0.pid_d.mult0.b[3] ;
 wire \top0.pid_d.mult0.b[4] ;
 wire \top0.pid_d.mult0.b[5] ;
 wire \top0.pid_d.mult0.b[6] ;
 wire \top0.pid_d.mult0.b[7] ;
 wire \top0.pid_d.mult0.b[8] ;
 wire \top0.pid_d.mult0.b[9] ;
 wire \top0.pid_d.out[0] ;
 wire \top0.pid_d.out[10] ;
 wire \top0.pid_d.out[11] ;
 wire \top0.pid_d.out[12] ;
 wire \top0.pid_d.out[13] ;
 wire \top0.pid_d.out[14] ;
 wire \top0.pid_d.out[15] ;
 wire \top0.pid_d.out[1] ;
 wire \top0.pid_d.out[2] ;
 wire \top0.pid_d.out[3] ;
 wire \top0.pid_d.out[4] ;
 wire \top0.pid_d.out[5] ;
 wire \top0.pid_d.out[6] ;
 wire \top0.pid_d.out[7] ;
 wire \top0.pid_d.out[8] ;
 wire \top0.pid_d.out[9] ;
 wire \top0.pid_d.out_valid ;
 wire \top0.pid_d.prev_error[0] ;
 wire \top0.pid_d.prev_error[10] ;
 wire \top0.pid_d.prev_error[11] ;
 wire \top0.pid_d.prev_error[12] ;
 wire \top0.pid_d.prev_error[13] ;
 wire \top0.pid_d.prev_error[14] ;
 wire \top0.pid_d.prev_error[15] ;
 wire \top0.pid_d.prev_error[1] ;
 wire \top0.pid_d.prev_error[2] ;
 wire \top0.pid_d.prev_error[3] ;
 wire \top0.pid_d.prev_error[4] ;
 wire \top0.pid_d.prev_error[5] ;
 wire \top0.pid_d.prev_error[6] ;
 wire \top0.pid_d.prev_error[7] ;
 wire \top0.pid_d.prev_error[8] ;
 wire \top0.pid_d.prev_error[9] ;
 wire \top0.pid_d.prev_int[0] ;
 wire \top0.pid_d.prev_int[10] ;
 wire \top0.pid_d.prev_int[11] ;
 wire \top0.pid_d.prev_int[12] ;
 wire \top0.pid_d.prev_int[13] ;
 wire \top0.pid_d.prev_int[14] ;
 wire \top0.pid_d.prev_int[15] ;
 wire \top0.pid_d.prev_int[1] ;
 wire \top0.pid_d.prev_int[2] ;
 wire \top0.pid_d.prev_int[3] ;
 wire \top0.pid_d.prev_int[4] ;
 wire \top0.pid_d.prev_int[5] ;
 wire \top0.pid_d.prev_int[6] ;
 wire \top0.pid_d.prev_int[7] ;
 wire \top0.pid_d.prev_int[8] ;
 wire \top0.pid_d.prev_int[9] ;
 wire \top0.pid_d.state[0] ;
 wire \top0.pid_d.state[1] ;
 wire \top0.pid_d.state[2] ;
 wire \top0.pid_d.state[3] ;
 wire \top0.pid_d.state[4] ;
 wire \top0.pid_d.state[5] ;
 wire \top0.pid_q.curr_error[0] ;
 wire \top0.pid_q.curr_error[10] ;
 wire \top0.pid_q.curr_error[11] ;
 wire \top0.pid_q.curr_error[12] ;
 wire \top0.pid_q.curr_error[13] ;
 wire \top0.pid_q.curr_error[14] ;
 wire \top0.pid_q.curr_error[15] ;
 wire \top0.pid_q.curr_error[1] ;
 wire \top0.pid_q.curr_error[2] ;
 wire \top0.pid_q.curr_error[3] ;
 wire \top0.pid_q.curr_error[4] ;
 wire \top0.pid_q.curr_error[5] ;
 wire \top0.pid_q.curr_error[6] ;
 wire \top0.pid_q.curr_error[7] ;
 wire \top0.pid_q.curr_error[8] ;
 wire \top0.pid_q.curr_error[9] ;
 wire \top0.pid_q.curr_int[0] ;
 wire \top0.pid_q.curr_int[10] ;
 wire \top0.pid_q.curr_int[11] ;
 wire \top0.pid_q.curr_int[12] ;
 wire \top0.pid_q.curr_int[13] ;
 wire \top0.pid_q.curr_int[14] ;
 wire \top0.pid_q.curr_int[15] ;
 wire \top0.pid_q.curr_int[1] ;
 wire \top0.pid_q.curr_int[2] ;
 wire \top0.pid_q.curr_int[3] ;
 wire \top0.pid_q.curr_int[4] ;
 wire \top0.pid_q.curr_int[5] ;
 wire \top0.pid_q.curr_int[6] ;
 wire \top0.pid_q.curr_int[7] ;
 wire \top0.pid_q.curr_int[8] ;
 wire \top0.pid_q.curr_int[9] ;
 wire \top0.pid_q.mult0.a[0] ;
 wire \top0.pid_q.mult0.a[10] ;
 wire \top0.pid_q.mult0.a[11] ;
 wire \top0.pid_q.mult0.a[12] ;
 wire \top0.pid_q.mult0.a[13] ;
 wire \top0.pid_q.mult0.a[14] ;
 wire \top0.pid_q.mult0.a[15] ;
 wire \top0.pid_q.mult0.a[1] ;
 wire \top0.pid_q.mult0.a[2] ;
 wire \top0.pid_q.mult0.a[3] ;
 wire \top0.pid_q.mult0.a[4] ;
 wire \top0.pid_q.mult0.a[5] ;
 wire \top0.pid_q.mult0.a[6] ;
 wire \top0.pid_q.mult0.a[7] ;
 wire \top0.pid_q.mult0.a[8] ;
 wire \top0.pid_q.mult0.a[9] ;
 wire \top0.pid_q.mult0.b[0] ;
 wire \top0.pid_q.mult0.b[10] ;
 wire \top0.pid_q.mult0.b[11] ;
 wire \top0.pid_q.mult0.b[12] ;
 wire \top0.pid_q.mult0.b[13] ;
 wire \top0.pid_q.mult0.b[14] ;
 wire \top0.pid_q.mult0.b[15] ;
 wire \top0.pid_q.mult0.b[1] ;
 wire \top0.pid_q.mult0.b[2] ;
 wire \top0.pid_q.mult0.b[3] ;
 wire \top0.pid_q.mult0.b[4] ;
 wire \top0.pid_q.mult0.b[5] ;
 wire \top0.pid_q.mult0.b[6] ;
 wire \top0.pid_q.mult0.b[7] ;
 wire \top0.pid_q.mult0.b[8] ;
 wire \top0.pid_q.mult0.b[9] ;
 wire \top0.pid_q.out[0] ;
 wire \top0.pid_q.out[10] ;
 wire \top0.pid_q.out[11] ;
 wire \top0.pid_q.out[12] ;
 wire \top0.pid_q.out[13] ;
 wire \top0.pid_q.out[14] ;
 wire \top0.pid_q.out[15] ;
 wire \top0.pid_q.out[1] ;
 wire \top0.pid_q.out[2] ;
 wire \top0.pid_q.out[3] ;
 wire \top0.pid_q.out[4] ;
 wire \top0.pid_q.out[5] ;
 wire \top0.pid_q.out[6] ;
 wire \top0.pid_q.out[7] ;
 wire \top0.pid_q.out[8] ;
 wire \top0.pid_q.out[9] ;
 wire \top0.pid_q.prev_error[0] ;
 wire \top0.pid_q.prev_error[10] ;
 wire \top0.pid_q.prev_error[11] ;
 wire \top0.pid_q.prev_error[12] ;
 wire \top0.pid_q.prev_error[13] ;
 wire \top0.pid_q.prev_error[14] ;
 wire \top0.pid_q.prev_error[15] ;
 wire \top0.pid_q.prev_error[1] ;
 wire \top0.pid_q.prev_error[2] ;
 wire \top0.pid_q.prev_error[3] ;
 wire \top0.pid_q.prev_error[4] ;
 wire \top0.pid_q.prev_error[5] ;
 wire \top0.pid_q.prev_error[6] ;
 wire \top0.pid_q.prev_error[7] ;
 wire \top0.pid_q.prev_error[8] ;
 wire \top0.pid_q.prev_error[9] ;
 wire \top0.pid_q.prev_int[0] ;
 wire \top0.pid_q.prev_int[10] ;
 wire \top0.pid_q.prev_int[11] ;
 wire \top0.pid_q.prev_int[12] ;
 wire \top0.pid_q.prev_int[13] ;
 wire \top0.pid_q.prev_int[14] ;
 wire \top0.pid_q.prev_int[15] ;
 wire \top0.pid_q.prev_int[1] ;
 wire \top0.pid_q.prev_int[2] ;
 wire \top0.pid_q.prev_int[3] ;
 wire \top0.pid_q.prev_int[4] ;
 wire \top0.pid_q.prev_int[5] ;
 wire \top0.pid_q.prev_int[6] ;
 wire \top0.pid_q.prev_int[7] ;
 wire \top0.pid_q.prev_int[8] ;
 wire \top0.pid_q.prev_int[9] ;
 wire \top0.pid_q.state[0] ;
 wire \top0.pid_q.state[1] ;
 wire \top0.pid_q.state[2] ;
 wire \top0.pid_q.state[3] ;
 wire \top0.pid_q.state[4] ;
 wire \top0.pid_q.state[5] ;
 wire \top0.ready ;
 wire \top0.start_svm ;
 wire \top0.state[0] ;
 wire \top0.state[1] ;
 wire \top0.state[2] ;
 wire \top0.svm0.calc_ready ;
 wire \top0.svm0.counter[0] ;
 wire \top0.svm0.counter[10] ;
 wire \top0.svm0.counter[11] ;
 wire \top0.svm0.counter[12] ;
 wire \top0.svm0.counter[13] ;
 wire \top0.svm0.counter[14] ;
 wire \top0.svm0.counter[15] ;
 wire \top0.svm0.counter[1] ;
 wire \top0.svm0.counter[2] ;
 wire \top0.svm0.counter[3] ;
 wire \top0.svm0.counter[4] ;
 wire \top0.svm0.counter[5] ;
 wire \top0.svm0.counter[6] ;
 wire \top0.svm0.counter[7] ;
 wire \top0.svm0.counter[8] ;
 wire \top0.svm0.counter[9] ;
 wire \top0.svm0.delta[0] ;
 wire \top0.svm0.delta[10] ;
 wire \top0.svm0.delta[11] ;
 wire \top0.svm0.delta[12] ;
 wire \top0.svm0.delta[13] ;
 wire \top0.svm0.delta[14] ;
 wire \top0.svm0.delta[15] ;
 wire \top0.svm0.delta[1] ;
 wire \top0.svm0.delta[2] ;
 wire \top0.svm0.delta[3] ;
 wire \top0.svm0.delta[4] ;
 wire \top0.svm0.delta[5] ;
 wire \top0.svm0.delta[6] ;
 wire \top0.svm0.delta[7] ;
 wire \top0.svm0.delta[8] ;
 wire \top0.svm0.delta[9] ;
 wire \top0.svm0.out_valid ;
 wire \top0.svm0.rising ;
 wire \top0.svm0.state[0] ;
 wire \top0.svm0.state[1] ;
 wire \top0.svm0.state[2] ;
 wire \top0.svm0.tA[0] ;
 wire \top0.svm0.tA[10] ;
 wire \top0.svm0.tA[11] ;
 wire \top0.svm0.tA[12] ;
 wire \top0.svm0.tA[13] ;
 wire \top0.svm0.tA[14] ;
 wire \top0.svm0.tA[15] ;
 wire \top0.svm0.tA[1] ;
 wire \top0.svm0.tA[2] ;
 wire \top0.svm0.tA[3] ;
 wire \top0.svm0.tA[4] ;
 wire \top0.svm0.tA[5] ;
 wire \top0.svm0.tA[6] ;
 wire \top0.svm0.tA[7] ;
 wire \top0.svm0.tA[8] ;
 wire \top0.svm0.tA[9] ;
 wire \top0.svm0.tB[0] ;
 wire \top0.svm0.tB[10] ;
 wire \top0.svm0.tB[11] ;
 wire \top0.svm0.tB[12] ;
 wire \top0.svm0.tB[13] ;
 wire \top0.svm0.tB[14] ;
 wire \top0.svm0.tB[15] ;
 wire \top0.svm0.tB[1] ;
 wire \top0.svm0.tB[2] ;
 wire \top0.svm0.tB[3] ;
 wire \top0.svm0.tB[4] ;
 wire \top0.svm0.tB[5] ;
 wire \top0.svm0.tB[6] ;
 wire \top0.svm0.tB[7] ;
 wire \top0.svm0.tB[8] ;
 wire \top0.svm0.tB[9] ;
 wire \top0.svm0.tC[0] ;
 wire \top0.svm0.tC[10] ;
 wire \top0.svm0.tC[11] ;
 wire \top0.svm0.tC[12] ;
 wire \top0.svm0.tC[13] ;
 wire \top0.svm0.tC[14] ;
 wire \top0.svm0.tC[15] ;
 wire \top0.svm0.tC[1] ;
 wire \top0.svm0.tC[2] ;
 wire \top0.svm0.tC[3] ;
 wire \top0.svm0.tC[4] ;
 wire \top0.svm0.tC[5] ;
 wire \top0.svm0.tC[6] ;
 wire \top0.svm0.tC[7] ;
 wire \top0.svm0.tC[8] ;
 wire \top0.svm0.tC[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire clknet_leaf_0_clk_sys;
 wire clknet_leaf_1_clk_sys;
 wire clknet_leaf_2_clk_sys;
 wire clknet_leaf_3_clk_sys;
 wire clknet_leaf_4_clk_sys;
 wire clknet_leaf_5_clk_sys;
 wire clknet_leaf_6_clk_sys;
 wire clknet_leaf_7_clk_sys;
 wire clknet_leaf_8_clk_sys;
 wire clknet_leaf_9_clk_sys;
 wire clknet_leaf_10_clk_sys;
 wire clknet_leaf_11_clk_sys;
 wire clknet_leaf_12_clk_sys;
 wire clknet_leaf_13_clk_sys;
 wire clknet_leaf_14_clk_sys;
 wire clknet_leaf_15_clk_sys;
 wire clknet_leaf_16_clk_sys;
 wire clknet_leaf_17_clk_sys;
 wire clknet_leaf_18_clk_sys;
 wire clknet_leaf_20_clk_sys;
 wire clknet_leaf_21_clk_sys;
 wire clknet_leaf_22_clk_sys;
 wire clknet_leaf_23_clk_sys;
 wire clknet_leaf_24_clk_sys;
 wire clknet_leaf_25_clk_sys;
 wire clknet_leaf_26_clk_sys;
 wire clknet_leaf_27_clk_sys;
 wire clknet_leaf_28_clk_sys;
 wire clknet_leaf_29_clk_sys;
 wire clknet_leaf_30_clk_sys;
 wire clknet_leaf_31_clk_sys;
 wire clknet_leaf_32_clk_sys;
 wire clknet_leaf_33_clk_sys;
 wire clknet_leaf_36_clk_sys;
 wire clknet_leaf_37_clk_sys;
 wire clknet_leaf_38_clk_sys;
 wire clknet_leaf_39_clk_sys;
 wire clknet_leaf_40_clk_sys;
 wire clknet_leaf_41_clk_sys;
 wire clknet_leaf_42_clk_sys;
 wire clknet_leaf_43_clk_sys;
 wire clknet_leaf_44_clk_sys;
 wire clknet_leaf_45_clk_sys;
 wire clknet_leaf_46_clk_sys;
 wire clknet_leaf_47_clk_sys;
 wire clknet_leaf_48_clk_sys;
 wire clknet_leaf_49_clk_sys;
 wire clknet_leaf_50_clk_sys;
 wire clknet_leaf_51_clk_sys;
 wire clknet_leaf_52_clk_sys;
 wire clknet_leaf_53_clk_sys;
 wire clknet_leaf_54_clk_sys;
 wire clknet_leaf_55_clk_sys;
 wire clknet_leaf_56_clk_sys;
 wire clknet_leaf_57_clk_sys;
 wire clknet_leaf_58_clk_sys;
 wire clknet_leaf_59_clk_sys;
 wire clknet_leaf_60_clk_sys;
 wire clknet_leaf_61_clk_sys;
 wire clknet_leaf_62_clk_sys;
 wire clknet_leaf_63_clk_sys;
 wire clknet_leaf_64_clk_sys;
 wire clknet_leaf_65_clk_sys;
 wire clknet_leaf_66_clk_sys;
 wire clknet_leaf_67_clk_sys;
 wire clknet_leaf_68_clk_sys;
 wire clknet_leaf_69_clk_sys;
 wire clknet_leaf_70_clk_sys;
 wire clknet_leaf_71_clk_sys;
 wire clknet_leaf_72_clk_sys;
 wire clknet_leaf_73_clk_sys;
 wire clknet_leaf_74_clk_sys;
 wire clknet_leaf_75_clk_sys;
 wire clknet_leaf_76_clk_sys;
 wire clknet_leaf_77_clk_sys;
 wire clknet_leaf_78_clk_sys;
 wire clknet_leaf_79_clk_sys;
 wire clknet_leaf_80_clk_sys;
 wire clknet_leaf_81_clk_sys;
 wire clknet_leaf_82_clk_sys;
 wire clknet_leaf_83_clk_sys;
 wire clknet_leaf_84_clk_sys;
 wire clknet_leaf_85_clk_sys;
 wire clknet_leaf_86_clk_sys;
 wire clknet_leaf_87_clk_sys;
 wire clknet_leaf_88_clk_sys;
 wire clknet_leaf_89_clk_sys;
 wire clknet_leaf_90_clk_sys;
 wire clknet_leaf_91_clk_sys;
 wire clknet_leaf_92_clk_sys;
 wire clknet_leaf_93_clk_sys;
 wire clknet_leaf_94_clk_sys;
 wire clknet_leaf_96_clk_sys;
 wire clknet_leaf_97_clk_sys;
 wire clknet_leaf_98_clk_sys;
 wire clknet_leaf_99_clk_sys;
 wire clknet_leaf_100_clk_sys;
 wire clknet_leaf_101_clk_sys;
 wire clknet_leaf_102_clk_sys;
 wire clknet_leaf_103_clk_sys;
 wire clknet_leaf_104_clk_sys;
 wire clknet_leaf_105_clk_sys;
 wire clknet_leaf_106_clk_sys;
 wire clknet_leaf_107_clk_sys;
 wire clknet_leaf_108_clk_sys;
 wire clknet_leaf_109_clk_sys;
 wire clknet_leaf_110_clk_sys;
 wire clknet_0_clk_sys;
 wire clknet_3_0__leaf_clk_sys;
 wire clknet_3_1__leaf_clk_sys;
 wire clknet_3_2__leaf_clk_sys;
 wire clknet_3_3__leaf_clk_sys;
 wire clknet_3_4__leaf_clk_sys;
 wire clknet_3_5__leaf_clk_sys;
 wire clknet_3_6__leaf_clk_sys;
 wire clknet_3_7__leaf_clk_sys;
 wire clknet_0_clk_mosi;
 wire clknet_3_0__leaf_clk_mosi;
 wire clknet_3_1__leaf_clk_mosi;
 wire clknet_3_2__leaf_clk_mosi;
 wire clknet_3_3__leaf_clk_mosi;
 wire clknet_3_4__leaf_clk_mosi;
 wire clknet_3_5__leaf_clk_mosi;
 wire clknet_3_6__leaf_clk_mosi;
 wire clknet_3_7__leaf_clk_mosi;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;

 sky130_fd_sc_hd__inv_2 _13189_ (.A(\top0.matmul0.matmul_stage_inst.start ),
    .Y(_05421_));
 sky130_fd_sc_hd__a21o_1 _13190_ (.A1(\top0.matmul0.matmul_stage_inst.state[0] ),
    .A2(_05421_),
    .B1(\top0.matmul0.done_pass ),
    .X(_00014_));
 sky130_fd_sc_hd__inv_2 _13191_ (.A(\top0.ready ),
    .Y(_05422_));
 sky130_fd_sc_hd__and4b_1 _13192_ (.A_N(\spi0.cs_sync[2] ),
    .B(\spi0.opcode[6] ),
    .C(\spi0.opcode[7] ),
    .D(\spi0.cs_sync[1] ),
    .X(_05423_));
 sky130_fd_sc_hd__and4_1 _13193_ (.A(\spi0.opcode[0] ),
    .B(\spi0.opcode[2] ),
    .C(\spi0.opcode[3] ),
    .D(\spi0.opcode[4] ),
    .X(_05424_));
 sky130_fd_sc_hd__nand4_4 _13194_ (.A(\spi0.opcode[1] ),
    .B(\spi0.opcode[5] ),
    .C(_05423_),
    .D(_05424_),
    .Y(_05425_));
 sky130_fd_sc_hd__inv_2 _13195_ (.A(_05425_),
    .Y(_05426_));
 sky130_fd_sc_hd__a22o_1 _13196_ (.A1(net744),
    .A2(_05422_),
    .B1(\state[0] ),
    .B2(_05426_),
    .X(_00013_));
 sky130_fd_sc_hd__inv_2 _13197_ (.A(\top0.pid_d.iterate_enable ),
    .Y(_05427_));
 sky130_fd_sc_hd__or4_2 _13198_ (.A(\spi0.opcode[1] ),
    .B(\spi0.opcode[5] ),
    .C(\spi0.opcode[6] ),
    .D(\spi0.opcode[7] ),
    .X(_05428_));
 sky130_fd_sc_hd__or4_2 _13199_ (.A(\spi0.opcode[0] ),
    .B(\spi0.opcode[2] ),
    .C(\spi0.opcode[3] ),
    .D(\spi0.opcode[4] ),
    .X(_05429_));
 sky130_fd_sc_hd__nor4b_4 _13200_ (.A(\spi0.cs_sync[2] ),
    .B(_05428_),
    .C(_05429_),
    .D_N(\spi0.cs_sync[1] ),
    .Y(_05430_));
 sky130_fd_sc_hd__a211o_1 _13201_ (.A1(\top0.pid_q.state[0] ),
    .A2(_05427_),
    .B1(net16),
    .C1(net544),
    .X(_00018_));
 sky130_fd_sc_hd__a211o_1 _13202_ (.A1(\top0.pid_d.state[0] ),
    .A2(_05427_),
    .B1(net16),
    .C1(net433),
    .X(_00017_));
 sky130_fd_sc_hd__a22o_1 _13203_ (.A1(net744),
    .A2(\top0.ready ),
    .B1(\state[0] ),
    .B2(_05425_),
    .X(_00012_));
 sky130_fd_sc_hd__inv_2 _13204_ (.A(\top0.matmul0.done_pass ),
    .Y(_05431_));
 sky130_fd_sc_hd__a21o_1 _13205_ (.A1(_05431_),
    .A2(\top0.matmul0.state[1] ),
    .B1(net748),
    .X(_00016_));
 sky130_fd_sc_hd__inv_2 _13206_ (.A(\top0.matmul0.start ),
    .Y(_05432_));
 sky130_fd_sc_hd__and2_1 _13207_ (.A(\top0.matmul0.done_pass ),
    .B(\top0.matmul0.state[1] ),
    .X(_05433_));
 sky130_fd_sc_hd__buf_6 _13208_ (.A(_05433_),
    .X(_05434_));
 sky130_fd_sc_hd__clkbuf_8 _13209_ (.A(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__buf_4 _13210_ (.A(_05435_),
    .X(_05436_));
 sky130_fd_sc_hd__clkbuf_4 _13211_ (.A(_05436_),
    .X(_05437_));
 sky130_fd_sc_hd__clkbuf_4 _13212_ (.A(_05437_),
    .X(_05438_));
 sky130_fd_sc_hd__buf_4 _13213_ (.A(_05438_),
    .X(_05439_));
 sky130_fd_sc_hd__a21o_1 _13214_ (.A1(net997),
    .A2(_05432_),
    .B1(_05439_),
    .X(_00015_));
 sky130_fd_sc_hd__or4b_1 _13215_ (.A(\spi0.cs_sync[2] ),
    .B(_05428_),
    .C(_05429_),
    .D_N(\spi0.cs_sync[1] ),
    .X(_05440_));
 sky130_fd_sc_hd__clkbuf_4 _13216_ (.A(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__clkbuf_4 _13217_ (.A(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__buf_4 _13218_ (.A(_05442_),
    .X(_05443_));
 sky130_fd_sc_hd__clkbuf_2 _13219_ (.A(_05443_),
    .X(_05444_));
 sky130_fd_sc_hd__and3_1 _13220_ (.A(\top0.pid_d.state[0] ),
    .B(\top0.pid_d.iterate_enable ),
    .C(net1019),
    .X(_05445_));
 sky130_fd_sc_hd__clkbuf_1 _13221_ (.A(_05445_),
    .X(_00004_));
 sky130_fd_sc_hd__and2_1 _13222_ (.A(\top0.pid_d.state[3] ),
    .B(_05441_),
    .X(_05446_));
 sky130_fd_sc_hd__clkbuf_1 _13223_ (.A(_05446_),
    .X(_00003_));
 sky130_fd_sc_hd__and2_1 _13224_ (.A(net551),
    .B(_05441_),
    .X(_05447_));
 sky130_fd_sc_hd__buf_2 _13225_ (.A(_05447_),
    .X(_05448_));
 sky130_fd_sc_hd__clkbuf_4 _13226_ (.A(_05448_),
    .X(_00011_));
 sky130_fd_sc_hd__clkbuf_4 _13227_ (.A(_05443_),
    .X(_05449_));
 sky130_fd_sc_hd__and2_1 _13228_ (.A(net553),
    .B(_05449_),
    .X(_05450_));
 sky130_fd_sc_hd__clkbuf_1 _13229_ (.A(_05450_),
    .X(_00010_));
 sky130_fd_sc_hd__and3_1 _13230_ (.A(\top0.pid_q.state[0] ),
    .B(\top0.pid_d.iterate_enable ),
    .C(net1019),
    .X(_05451_));
 sky130_fd_sc_hd__clkbuf_1 _13231_ (.A(_05451_),
    .X(_00009_));
 sky130_fd_sc_hd__and2_1 _13232_ (.A(net547),
    .B(_05441_),
    .X(_05452_));
 sky130_fd_sc_hd__buf_1 _13233_ (.A(_05452_),
    .X(_00008_));
 sky130_fd_sc_hd__and2_1 _13234_ (.A(net543),
    .B(_05442_),
    .X(_05453_));
 sky130_fd_sc_hd__clkbuf_1 _13235_ (.A(_05453_),
    .X(_00007_));
 sky130_fd_sc_hd__and2_1 _13236_ (.A(net437),
    .B(_05441_),
    .X(_05454_));
 sky130_fd_sc_hd__buf_1 _13237_ (.A(_05454_),
    .X(_00006_));
 sky130_fd_sc_hd__and2_1 _13238_ (.A(net441),
    .B(_05449_),
    .X(_05455_));
 sky130_fd_sc_hd__clkbuf_1 _13239_ (.A(_05455_),
    .X(_00005_));
 sky130_fd_sc_hd__nand2_4 _13240_ (.A(\top0.matmul0.matmul_stage_inst.state[0] ),
    .B(\top0.matmul0.matmul_stage_inst.start ),
    .Y(_05456_));
 sky130_fd_sc_hd__inv_2 _13241_ (.A(_05456_),
    .Y(_05457_));
 sky130_fd_sc_hd__clkbuf_4 _13242_ (.A(_05457_),
    .X(_05458_));
 sky130_fd_sc_hd__clkbuf_4 _13243_ (.A(_05458_),
    .X(_00000_));
 sky130_fd_sc_hd__and2_1 _13244_ (.A(\top0.pid_d.state[5] ),
    .B(net1019),
    .X(_05459_));
 sky130_fd_sc_hd__clkbuf_1 _13245_ (.A(_05459_),
    .X(_00002_));
 sky130_fd_sc_hd__nand2_4 _13246_ (.A(\top0.matmul0.state[0] ),
    .B(\top0.matmul0.start ),
    .Y(_05460_));
 sky130_fd_sc_hd__buf_4 _13247_ (.A(_05460_),
    .X(_05461_));
 sky130_fd_sc_hd__inv_2 _13248_ (.A(_05461_),
    .Y(_00001_));
 sky130_fd_sc_hd__and3b_1 _13249_ (.A_N(net173),
    .B(\top0.svm0.state[1] ),
    .C(\top0.svm0.state[0] ),
    .X(_05462_));
 sky130_fd_sc_hd__buf_6 _13250_ (.A(_05462_),
    .X(_05463_));
 sky130_fd_sc_hd__clkbuf_8 _13251_ (.A(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__buf_4 _13252_ (.A(_05464_),
    .X(_05465_));
 sky130_fd_sc_hd__clkbuf_4 _13253_ (.A(_05433_),
    .X(_05466_));
 sky130_fd_sc_hd__nor3b_4 _13254_ (.A(net173),
    .B(\top0.svm0.state[1] ),
    .C_N(\top0.svm0.state[0] ),
    .Y(_05467_));
 sky130_fd_sc_hd__and3_1 _13255_ (.A(net76),
    .B(_05466_),
    .C(_05467_),
    .X(_05468_));
 sky130_fd_sc_hd__nor3b_4 _13256_ (.A(net173),
    .B(\top0.svm0.state[0] ),
    .C_N(\top0.svm0.state[1] ),
    .Y(_05469_));
 sky130_fd_sc_hd__buf_6 _13257_ (.A(_05469_),
    .X(_05470_));
 sky130_fd_sc_hd__a32o_1 _13258_ (.A1(\top0.matmul0.beta_pass[5] ),
    .A2(_05466_),
    .A3(_05470_),
    .B1(_05464_),
    .B2(\top0.c_out_calc[5] ),
    .X(_05471_));
 sky130_fd_sc_hd__nor2_4 _13259_ (.A(_05468_),
    .B(_05471_),
    .Y(_05472_));
 sky130_fd_sc_hd__nand2_2 _13260_ (.A(net47),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__buf_6 _13261_ (.A(_05467_),
    .X(_05474_));
 sky130_fd_sc_hd__nand3_2 _13262_ (.A(\top0.matmul0.alpha_pass[4] ),
    .B(_05466_),
    .C(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__a32oi_4 _13263_ (.A1(\top0.matmul0.beta_pass[4] ),
    .A2(_05434_),
    .A3(_05470_),
    .B1(_05463_),
    .B2(\top0.c_out_calc[4] ),
    .Y(_05476_));
 sky130_fd_sc_hd__and3_1 _13264_ (.A(net43),
    .B(_05475_),
    .C(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__nand3_2 _13265_ (.A(\top0.matmul0.alpha_pass[3] ),
    .B(_05466_),
    .C(_05474_),
    .Y(_05478_));
 sky130_fd_sc_hd__a32oi_4 _13266_ (.A1(\top0.matmul0.beta_pass[3] ),
    .A2(_05434_),
    .A3(_05469_),
    .B1(_05463_),
    .B2(\top0.c_out_calc[3] ),
    .Y(_05479_));
 sky130_fd_sc_hd__and3_1 _13267_ (.A(net42),
    .B(_05478_),
    .C(_05479_),
    .X(_05480_));
 sky130_fd_sc_hd__xor2_1 _13268_ (.A(_05477_),
    .B(_05480_),
    .X(_05481_));
 sky130_fd_sc_hd__xnor2_2 _13269_ (.A(_05473_),
    .B(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__nand3_1 _13270_ (.A(\top0.matmul0.alpha_pass[0] ),
    .B(_05435_),
    .C(_05474_),
    .Y(_05483_));
 sky130_fd_sc_hd__clkbuf_4 _13271_ (.A(_05483_),
    .X(_05484_));
 sky130_fd_sc_hd__a32oi_2 _13272_ (.A1(\top0.matmul0.beta_pass[0] ),
    .A2(_05435_),
    .A3(_05470_),
    .B1(_05464_),
    .B2(\top0.c_out_calc[0] ),
    .Y(_05485_));
 sky130_fd_sc_hd__buf_2 _13273_ (.A(_05485_),
    .X(_05486_));
 sky130_fd_sc_hd__and3_1 _13274_ (.A(net38),
    .B(_05484_),
    .C(_05486_),
    .X(_05487_));
 sky130_fd_sc_hd__nand3_2 _13275_ (.A(\top0.matmul0.alpha_pass[1] ),
    .B(_05435_),
    .C(_05474_),
    .Y(_05488_));
 sky130_fd_sc_hd__buf_2 _13276_ (.A(_05488_),
    .X(_05489_));
 sky130_fd_sc_hd__a32oi_4 _13277_ (.A1(\top0.matmul0.beta_pass[1] ),
    .A2(_05466_),
    .A3(_05470_),
    .B1(_05464_),
    .B2(\top0.c_out_calc[1] ),
    .Y(_05490_));
 sky130_fd_sc_hd__buf_2 _13278_ (.A(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__and3_1 _13279_ (.A(net40),
    .B(_05489_),
    .C(_05491_),
    .X(_05492_));
 sky130_fd_sc_hd__and3_1 _13280_ (.A(\top0.matmul0.alpha_pass[2] ),
    .B(_05466_),
    .C(_05474_),
    .X(_05493_));
 sky130_fd_sc_hd__a32o_1 _13281_ (.A1(\top0.matmul0.beta_pass[2] ),
    .A2(_05466_),
    .A3(_05470_),
    .B1(_05463_),
    .B2(\top0.c_out_calc[2] ),
    .X(_05494_));
 sky130_fd_sc_hd__nor2_1 _13282_ (.A(_05493_),
    .B(_05494_),
    .Y(_05495_));
 sky130_fd_sc_hd__clkbuf_4 _13283_ (.A(_05495_),
    .X(_05496_));
 sky130_fd_sc_hd__clkbuf_4 _13284_ (.A(_05496_),
    .X(_05497_));
 sky130_fd_sc_hd__o211a_1 _13285_ (.A1(_05487_),
    .A2(_05492_),
    .B1(_05497_),
    .C1(net42),
    .X(_05498_));
 sky130_fd_sc_hd__a21o_1 _13286_ (.A1(_05487_),
    .A2(_05492_),
    .B1(_05498_),
    .X(_05499_));
 sky130_fd_sc_hd__clkinv_4 _13287_ (.A(net33),
    .Y(_05500_));
 sky130_fd_sc_hd__nand2_1 _13288_ (.A(_05484_),
    .B(_05486_),
    .Y(_05501_));
 sky130_fd_sc_hd__nor2_1 _13289_ (.A(_05500_),
    .B(_05501_),
    .Y(_05502_));
 sky130_fd_sc_hd__and3_1 _13290_ (.A(net38),
    .B(_05489_),
    .C(_05491_),
    .X(_05503_));
 sky130_fd_sc_hd__inv_1 _13291_ (.A(net40),
    .Y(_05504_));
 sky130_fd_sc_hd__nor3_1 _13292_ (.A(_05504_),
    .B(_05493_),
    .C(_05494_),
    .Y(_05505_));
 sky130_fd_sc_hd__xnor2_1 _13293_ (.A(_05503_),
    .B(_05505_),
    .Y(_05506_));
 sky130_fd_sc_hd__xnor2_2 _13294_ (.A(_05502_),
    .B(_05506_),
    .Y(_05507_));
 sky130_fd_sc_hd__xnor2_1 _13295_ (.A(_05499_),
    .B(_05507_),
    .Y(_05508_));
 sky130_fd_sc_hd__xnor2_2 _13296_ (.A(_05482_),
    .B(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hd__nand2_1 _13297_ (.A(net42),
    .B(_05497_),
    .Y(_05510_));
 sky130_fd_sc_hd__xor2_1 _13298_ (.A(_05487_),
    .B(_05492_),
    .X(_05511_));
 sky130_fd_sc_hd__xnor2_2 _13299_ (.A(_05510_),
    .B(_05511_),
    .Y(_05512_));
 sky130_fd_sc_hd__and3_1 _13300_ (.A(net42),
    .B(_05489_),
    .C(_05491_),
    .X(_05513_));
 sky130_fd_sc_hd__and3_1 _13301_ (.A(net40),
    .B(_05484_),
    .C(_05486_),
    .X(_05514_));
 sky130_fd_sc_hd__a22o_1 _13302_ (.A1(net43),
    .A2(_05497_),
    .B1(_05513_),
    .B2(_05514_),
    .X(_05515_));
 sky130_fd_sc_hd__o21a_1 _13303_ (.A1(_05513_),
    .A2(_05514_),
    .B1(_05515_),
    .X(_05516_));
 sky130_fd_sc_hd__clkbuf_4 _13304_ (.A(_05472_),
    .X(_05517_));
 sky130_fd_sc_hd__buf_1 _13305_ (.A(_05517_),
    .X(_05518_));
 sky130_fd_sc_hd__nand2_2 _13306_ (.A(net49),
    .B(net1015),
    .Y(_05519_));
 sky130_fd_sc_hd__buf_2 _13307_ (.A(_05475_),
    .X(_05520_));
 sky130_fd_sc_hd__buf_2 _13308_ (.A(_05476_),
    .X(_05521_));
 sky130_fd_sc_hd__and3_1 _13309_ (.A(net47),
    .B(_05520_),
    .C(_05521_),
    .X(_05522_));
 sky130_fd_sc_hd__buf_2 _13310_ (.A(_05478_),
    .X(_05523_));
 sky130_fd_sc_hd__buf_2 _13311_ (.A(_05479_),
    .X(_05524_));
 sky130_fd_sc_hd__and3_1 _13312_ (.A(net43),
    .B(_05523_),
    .C(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__xor2_2 _13313_ (.A(_05522_),
    .B(_05525_),
    .X(_05526_));
 sky130_fd_sc_hd__xnor2_4 _13314_ (.A(_05519_),
    .B(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__a21o_1 _13315_ (.A1(_05512_),
    .A2(_05516_),
    .B1(_05527_),
    .X(_05528_));
 sky130_fd_sc_hd__o21a_1 _13316_ (.A1(_05512_),
    .A2(_05516_),
    .B1(_05528_),
    .X(_05529_));
 sky130_fd_sc_hd__inv_2 _13317_ (.A(net48),
    .Y(_05530_));
 sky130_fd_sc_hd__and3_2 _13318_ (.A(\top0.matmul0.alpha_pass[6] ),
    .B(_05434_),
    .C(_05467_),
    .X(_05531_));
 sky130_fd_sc_hd__a32o_2 _13319_ (.A1(\top0.matmul0.beta_pass[6] ),
    .A2(_05434_),
    .A3(_05469_),
    .B1(_05463_),
    .B2(\top0.c_out_calc[6] ),
    .X(_05532_));
 sky130_fd_sc_hd__or2_1 _13320_ (.A(_05531_),
    .B(_05532_),
    .X(_05533_));
 sky130_fd_sc_hd__buf_6 _13321_ (.A(_05533_),
    .X(_05534_));
 sky130_fd_sc_hd__nor2_1 _13322_ (.A(_05530_),
    .B(_05534_),
    .Y(_05535_));
 sky130_fd_sc_hd__inv_2 _13323_ (.A(net54),
    .Y(_05536_));
 sky130_fd_sc_hd__and3_1 _13324_ (.A(\top0.matmul0.beta_pass[8] ),
    .B(_05434_),
    .C(_05469_),
    .X(_05537_));
 sky130_fd_sc_hd__buf_6 _13325_ (.A(_05537_),
    .X(_05538_));
 sky130_fd_sc_hd__a32o_2 _13326_ (.A1(net1024),
    .A2(_05466_),
    .A3(_05467_),
    .B1(_05464_),
    .B2(\top0.c_out_calc[8] ),
    .X(_05539_));
 sky130_fd_sc_hd__nor3_1 _13327_ (.A(_05536_),
    .B(_05538_),
    .C(_05539_),
    .Y(_05540_));
 sky130_fd_sc_hd__inv_2 _13328_ (.A(net51),
    .Y(_05541_));
 sky130_fd_sc_hd__and3_1 _13329_ (.A(\top0.matmul0.alpha_pass[7] ),
    .B(_05434_),
    .C(_05467_),
    .X(_05542_));
 sky130_fd_sc_hd__buf_6 _13330_ (.A(_05542_),
    .X(_05543_));
 sky130_fd_sc_hd__a32o_1 _13331_ (.A1(\top0.matmul0.beta_pass[7] ),
    .A2(_05434_),
    .A3(_05469_),
    .B1(_05463_),
    .B2(\top0.c_out_calc[7] ),
    .X(_05544_));
 sky130_fd_sc_hd__buf_6 _13332_ (.A(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__or3_1 _13333_ (.A(_05541_),
    .B(_05543_),
    .C(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__xor2_1 _13334_ (.A(_05540_),
    .B(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__xnor2_2 _13335_ (.A(_05535_),
    .B(_05547_),
    .Y(_05548_));
 sky130_fd_sc_hd__or3_1 _13336_ (.A(_05541_),
    .B(_05531_),
    .C(_05532_),
    .X(_05549_));
 sky130_fd_sc_hd__or3_1 _13337_ (.A(_05536_),
    .B(_05543_),
    .C(_05545_),
    .X(_05550_));
 sky130_fd_sc_hd__nor2_2 _13338_ (.A(_05538_),
    .B(_05539_),
    .Y(_05551_));
 sky130_fd_sc_hd__o2bb2a_1 _13339_ (.A1_N(net57),
    .A2_N(_05551_),
    .B1(_05549_),
    .B2(_05550_),
    .X(_05552_));
 sky130_fd_sc_hd__a21o_1 _13340_ (.A1(_05549_),
    .A2(_05550_),
    .B1(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__o211a_1 _13341_ (.A1(_05522_),
    .A2(_05525_),
    .B1(net50),
    .C1(net1015),
    .X(_05554_));
 sky130_fd_sc_hd__a21o_1 _13342_ (.A1(_05522_),
    .A2(_05525_),
    .B1(_05554_),
    .X(_05555_));
 sky130_fd_sc_hd__xnor2_1 _13343_ (.A(_05553_),
    .B(_05555_),
    .Y(_05556_));
 sky130_fd_sc_hd__xnor2_1 _13344_ (.A(_05548_),
    .B(_05556_),
    .Y(_05557_));
 sky130_fd_sc_hd__xor2_1 _13345_ (.A(_05529_),
    .B(_05557_),
    .X(_05558_));
 sky130_fd_sc_hd__xnor2_2 _13346_ (.A(_05509_),
    .B(_05558_),
    .Y(_05559_));
 sky130_fd_sc_hd__nand2_1 _13347_ (.A(net52),
    .B(_05517_),
    .Y(_05560_));
 sky130_fd_sc_hd__and3_1 _13348_ (.A(net50),
    .B(_05520_),
    .C(_05521_),
    .X(_05561_));
 sky130_fd_sc_hd__and3_1 _13349_ (.A(net47),
    .B(_05523_),
    .C(_05524_),
    .X(_05562_));
 sky130_fd_sc_hd__xor2_1 _13350_ (.A(_05561_),
    .B(_05562_),
    .X(_05563_));
 sky130_fd_sc_hd__xnor2_2 _13351_ (.A(_05560_),
    .B(_05563_),
    .Y(_05564_));
 sky130_fd_sc_hd__inv_2 _13352_ (.A(net43),
    .Y(_05565_));
 sky130_fd_sc_hd__or2_1 _13353_ (.A(_05493_),
    .B(_05494_),
    .X(_05566_));
 sky130_fd_sc_hd__buf_2 _13354_ (.A(_05566_),
    .X(_05567_));
 sky130_fd_sc_hd__nor2_1 _13355_ (.A(_05565_),
    .B(_05567_),
    .Y(_05568_));
 sky130_fd_sc_hd__xnor2_1 _13356_ (.A(_05513_),
    .B(_05514_),
    .Y(_05569_));
 sky130_fd_sc_hd__xnor2_2 _13357_ (.A(_05568_),
    .B(_05569_),
    .Y(_05570_));
 sky130_fd_sc_hd__and3_1 _13358_ (.A(net43),
    .B(_05489_),
    .C(_05491_),
    .X(_05571_));
 sky130_fd_sc_hd__and3_1 _13359_ (.A(net42),
    .B(_05484_),
    .C(_05486_),
    .X(_05572_));
 sky130_fd_sc_hd__inv_2 _13360_ (.A(net46),
    .Y(_05573_));
 sky130_fd_sc_hd__nor2_1 _13361_ (.A(_05573_),
    .B(_05567_),
    .Y(_05574_));
 sky130_fd_sc_hd__a21o_1 _13362_ (.A1(_05571_),
    .A2(_05572_),
    .B1(_05574_),
    .X(_05575_));
 sky130_fd_sc_hd__o21ai_1 _13363_ (.A1(_05571_),
    .A2(_05572_),
    .B1(_05575_),
    .Y(_05576_));
 sky130_fd_sc_hd__a21bo_1 _13364_ (.A1(_05564_),
    .A2(_05570_),
    .B1_N(_05576_),
    .X(_05577_));
 sky130_fd_sc_hd__o21a_1 _13365_ (.A1(_05564_),
    .A2(_05570_),
    .B1(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__clkbuf_4 _13366_ (.A(_05551_),
    .X(_05579_));
 sky130_fd_sc_hd__nand2_1 _13367_ (.A(net57),
    .B(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__xnor2_1 _13368_ (.A(_05549_),
    .B(_05550_),
    .Y(_05581_));
 sky130_fd_sc_hd__xnor2_2 _13369_ (.A(_05580_),
    .B(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__o211a_1 _13370_ (.A1(_05561_),
    .A2(_05562_),
    .B1(net52),
    .C1(_05518_),
    .X(_05583_));
 sky130_fd_sc_hd__a21o_1 _13371_ (.A1(_05561_),
    .A2(_05562_),
    .B1(_05583_),
    .X(_05584_));
 sky130_fd_sc_hd__nor2_2 _13372_ (.A(_05531_),
    .B(_05532_),
    .Y(_05585_));
 sky130_fd_sc_hd__buf_4 _13373_ (.A(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__nor2_2 _13374_ (.A(_05543_),
    .B(_05545_),
    .Y(_05587_));
 sky130_fd_sc_hd__clkbuf_4 _13375_ (.A(_05587_),
    .X(_05588_));
 sky130_fd_sc_hd__a22o_1 _13376_ (.A1(net54),
    .A2(_05586_),
    .B1(_05588_),
    .B2(net57),
    .X(_05589_));
 sky130_fd_sc_hd__and2_1 _13377_ (.A(net61),
    .B(_05551_),
    .X(_05590_));
 sky130_fd_sc_hd__a41o_1 _13378_ (.A1(net57),
    .A2(net54),
    .A3(_05586_),
    .A4(_05588_),
    .B1(_05590_),
    .X(_05591_));
 sky130_fd_sc_hd__nand2_1 _13379_ (.A(_05589_),
    .B(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__xnor2_1 _13380_ (.A(_05584_),
    .B(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__xnor2_2 _13381_ (.A(_05582_),
    .B(_05593_),
    .Y(_05594_));
 sky130_fd_sc_hd__xnor2_2 _13382_ (.A(_05512_),
    .B(_05516_),
    .Y(_05595_));
 sky130_fd_sc_hd__xnor2_4 _13383_ (.A(_05527_),
    .B(_05595_),
    .Y(_05596_));
 sky130_fd_sc_hd__a21o_1 _13384_ (.A1(_05578_),
    .A2(_05594_),
    .B1(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__o21a_1 _13385_ (.A1(_05578_),
    .A2(_05594_),
    .B1(_05597_),
    .X(_05598_));
 sky130_fd_sc_hd__nand3b_1 _13386_ (.A_N(\top0.svm0.state[1] ),
    .B(\top0.svm0.state[0] ),
    .C(\top0.matmul0.alpha_pass[10] ),
    .Y(_05599_));
 sky130_fd_sc_hd__nand3b_1 _13387_ (.A_N(\top0.svm0.state[0] ),
    .B(net430),
    .C(\top0.svm0.state[1] ),
    .Y(_05600_));
 sky130_fd_sc_hd__nand2_4 _13388_ (.A(\top0.matmul0.done_pass ),
    .B(\top0.matmul0.state[1] ),
    .Y(_05601_));
 sky130_fd_sc_hd__a211o_2 _13389_ (.A1(_05599_),
    .A2(_05600_),
    .B1(net173),
    .C1(_05601_),
    .X(_05602_));
 sky130_fd_sc_hd__nand2_4 _13390_ (.A(\top0.c_out_calc[10] ),
    .B(_05464_),
    .Y(_05603_));
 sky130_fd_sc_hd__and2_1 _13391_ (.A(_05602_),
    .B(_05603_),
    .X(_05604_));
 sky130_fd_sc_hd__buf_4 _13392_ (.A(_05604_),
    .X(_05605_));
 sky130_fd_sc_hd__nand2_2 _13393_ (.A(net61),
    .B(_05605_),
    .Y(_05606_));
 sky130_fd_sc_hd__inv_2 _13394_ (.A(net63),
    .Y(_05607_));
 sky130_fd_sc_hd__and3_2 _13395_ (.A(\top0.matmul0.alpha_pass[11] ),
    .B(_05434_),
    .C(_05467_),
    .X(_05608_));
 sky130_fd_sc_hd__a32o_2 _13396_ (.A1(\top0.matmul0.beta_pass[11] ),
    .A2(_05434_),
    .A3(_05469_),
    .B1(_05463_),
    .B2(\top0.c_out_calc[11] ),
    .X(_05609_));
 sky130_fd_sc_hd__or3_2 _13397_ (.A(_05607_),
    .B(_05608_),
    .C(_05609_),
    .X(_05610_));
 sky130_fd_sc_hd__nand3_4 _13398_ (.A(\top0.matmul0.alpha_pass[9] ),
    .B(_05435_),
    .C(_05474_),
    .Y(_05611_));
 sky130_fd_sc_hd__a32oi_4 _13399_ (.A1(\top0.matmul0.beta_pass[9] ),
    .A2(_05435_),
    .A3(_05470_),
    .B1(_05464_),
    .B2(\top0.c_out_calc[9] ),
    .Y(_05612_));
 sky130_fd_sc_hd__and3_2 _13400_ (.A(net56),
    .B(_05611_),
    .C(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__xnor2_4 _13401_ (.A(_05610_),
    .B(_05613_),
    .Y(_05614_));
 sky130_fd_sc_hd__xnor2_4 _13402_ (.A(_05606_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__nand3_1 _13403_ (.A(\top0.matmul0.alpha_pass[12] ),
    .B(_05435_),
    .C(_05474_),
    .Y(_05616_));
 sky130_fd_sc_hd__a32oi_4 _13404_ (.A1(\top0.matmul0.beta_pass[12] ),
    .A2(_05435_),
    .A3(_05470_),
    .B1(_05464_),
    .B2(\top0.c_out_calc[12] ),
    .Y(_05617_));
 sky130_fd_sc_hd__and2_1 _13405_ (.A(_05616_),
    .B(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__buf_4 _13406_ (.A(_05618_),
    .X(_05619_));
 sky130_fd_sc_hd__and3_1 _13407_ (.A(net64),
    .B(_05602_),
    .C(_05603_),
    .X(_05620_));
 sky130_fd_sc_hd__buf_2 _13408_ (.A(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__and3_2 _13409_ (.A(net60),
    .B(_05611_),
    .C(_05612_),
    .X(_05622_));
 sky130_fd_sc_hd__nor2_1 _13410_ (.A(_05621_),
    .B(_05622_),
    .Y(_05623_));
 sky130_fd_sc_hd__nor2_2 _13411_ (.A(_05608_),
    .B(_05609_),
    .Y(_05624_));
 sky130_fd_sc_hd__buf_4 _13412_ (.A(_05624_),
    .X(_05625_));
 sky130_fd_sc_hd__clkbuf_4 _13413_ (.A(_05625_),
    .X(_05626_));
 sky130_fd_sc_hd__a21oi_1 _13414_ (.A1(_05621_),
    .A2(_05622_),
    .B1(_05626_),
    .Y(_05627_));
 sky130_fd_sc_hd__nor2_1 _13415_ (.A(_05623_),
    .B(_05627_),
    .Y(_05628_));
 sky130_fd_sc_hd__or2_2 _13416_ (.A(_05608_),
    .B(_05609_),
    .X(_05629_));
 sky130_fd_sc_hd__nor2_1 _13417_ (.A(_05629_),
    .B(_05623_),
    .Y(_05630_));
 sky130_fd_sc_hd__a21o_1 _13418_ (.A1(_05621_),
    .A2(_05622_),
    .B1(_05619_),
    .X(_05631_));
 sky130_fd_sc_hd__a21o_1 _13419_ (.A1(_05621_),
    .A2(_05622_),
    .B1(net65),
    .X(_05632_));
 sky130_fd_sc_hd__o21a_1 _13420_ (.A1(_05630_),
    .A2(_05631_),
    .B1(_05632_),
    .X(_05633_));
 sky130_fd_sc_hd__inv_2 _13421_ (.A(_05633_),
    .Y(_05634_));
 sky130_fd_sc_hd__a31o_1 _13422_ (.A1(net65),
    .A2(_05619_),
    .A3(_05628_),
    .B1(_05634_),
    .X(_05635_));
 sky130_fd_sc_hd__xnor2_2 _13423_ (.A(_05615_),
    .B(_05635_),
    .Y(_05636_));
 sky130_fd_sc_hd__and3_2 _13424_ (.A(\top0.matmul0.alpha_pass[9] ),
    .B(_05466_),
    .C(_05467_),
    .X(_05637_));
 sky130_fd_sc_hd__a32o_1 _13425_ (.A1(\top0.matmul0.beta_pass[9] ),
    .A2(_05466_),
    .A3(_05470_),
    .B1(_05463_),
    .B2(\top0.c_out_calc[9] ),
    .X(_05638_));
 sky130_fd_sc_hd__nor2_4 _13426_ (.A(_05637_),
    .B(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__clkbuf_4 _13427_ (.A(_05639_),
    .X(_05640_));
 sky130_fd_sc_hd__xnor2_1 _13428_ (.A(net61),
    .B(_05625_),
    .Y(_05641_));
 sky130_fd_sc_hd__and3_1 _13429_ (.A(_05605_),
    .B(_05640_),
    .C(_05641_),
    .X(_05642_));
 sky130_fd_sc_hd__and3_1 _13430_ (.A(net65),
    .B(net63),
    .C(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__a21bo_1 _13431_ (.A1(_05582_),
    .A2(_05592_),
    .B1_N(_05584_),
    .X(_05644_));
 sky130_fd_sc_hd__o21a_1 _13432_ (.A1(_05582_),
    .A2(_05592_),
    .B1(_05644_),
    .X(_05645_));
 sky130_fd_sc_hd__xnor2_1 _13433_ (.A(_05643_),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__xnor2_1 _13434_ (.A(_05636_),
    .B(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__a21bo_1 _13435_ (.A1(_05559_),
    .A2(_05598_),
    .B1_N(_05647_),
    .X(_05648_));
 sky130_fd_sc_hd__o21ai_2 _13436_ (.A1(_05559_),
    .A2(_05598_),
    .B1(_05648_),
    .Y(_05649_));
 sky130_fd_sc_hd__a21bo_1 _13437_ (.A1(_05643_),
    .A2(_05636_),
    .B1_N(_05645_),
    .X(_05650_));
 sky130_fd_sc_hd__o21ai_2 _13438_ (.A1(_05643_),
    .A2(_05636_),
    .B1(_05650_),
    .Y(_05651_));
 sky130_fd_sc_hd__a21o_1 _13439_ (.A1(_05619_),
    .A2(_05628_),
    .B1(_05615_),
    .X(_05652_));
 sky130_fd_sc_hd__o211ai_4 _13440_ (.A1(net65),
    .A2(_05615_),
    .B1(_05652_),
    .C1(_05633_),
    .Y(_05653_));
 sky130_fd_sc_hd__a21bo_1 _13441_ (.A1(_05548_),
    .A2(_05555_),
    .B1_N(_05553_),
    .X(_05654_));
 sky130_fd_sc_hd__o21ai_2 _13442_ (.A1(_05548_),
    .A2(_05555_),
    .B1(_05654_),
    .Y(_05655_));
 sky130_fd_sc_hd__and3_1 _13443_ (.A(net56),
    .B(_05602_),
    .C(_05603_),
    .X(_05656_));
 sky130_fd_sc_hd__inv_2 _13444_ (.A(net60),
    .Y(_05657_));
 sky130_fd_sc_hd__or3_1 _13445_ (.A(_05657_),
    .B(_05608_),
    .C(_05609_),
    .X(_05658_));
 sky130_fd_sc_hd__or3_1 _13446_ (.A(_05536_),
    .B(_05637_),
    .C(_05638_),
    .X(_05659_));
 sky130_fd_sc_hd__xor2_1 _13447_ (.A(_05658_),
    .B(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__xnor2_2 _13448_ (.A(_05656_),
    .B(_05660_),
    .Y(_05661_));
 sky130_fd_sc_hd__inv_2 _13449_ (.A(\top0.matmul0.beta_pass[13] ),
    .Y(_05662_));
 sky130_fd_sc_hd__or3b_1 _13450_ (.A(_05662_),
    .B(_05601_),
    .C_N(_05470_),
    .X(_05663_));
 sky130_fd_sc_hd__a32oi_4 _13451_ (.A1(\top0.matmul0.alpha_pass[13] ),
    .A2(_05435_),
    .A3(_05474_),
    .B1(_05464_),
    .B2(\top0.c_out_calc[13] ),
    .Y(_05664_));
 sky130_fd_sc_hd__and2_1 _13452_ (.A(_05663_),
    .B(_05664_),
    .X(_05665_));
 sky130_fd_sc_hd__buf_4 _13453_ (.A(_05665_),
    .X(_05666_));
 sky130_fd_sc_hd__nand2_1 _13454_ (.A(net65),
    .B(_05666_),
    .Y(_05667_));
 sky130_fd_sc_hd__nand2_1 _13455_ (.A(net63),
    .B(_05619_),
    .Y(_05668_));
 sky130_fd_sc_hd__xnor2_1 _13456_ (.A(_05667_),
    .B(_05668_),
    .Y(_05669_));
 sky130_fd_sc_hd__a32o_1 _13457_ (.A1(net60),
    .A2(_05604_),
    .A3(_05613_),
    .B1(_05624_),
    .B2(net64),
    .X(_05670_));
 sky130_fd_sc_hd__a21o_1 _13458_ (.A1(net60),
    .A2(_05604_),
    .B1(_05613_),
    .X(_05671_));
 sky130_fd_sc_hd__nand2_2 _13459_ (.A(_05670_),
    .B(_05671_),
    .Y(_05672_));
 sky130_fd_sc_hd__xnor2_1 _13460_ (.A(_05669_),
    .B(_05672_),
    .Y(_05673_));
 sky130_fd_sc_hd__xor2_1 _13461_ (.A(_05661_),
    .B(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__xnor2_1 _13462_ (.A(_05655_),
    .B(_05674_),
    .Y(_05675_));
 sky130_fd_sc_hd__xnor2_1 _13463_ (.A(_05653_),
    .B(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__nand2_1 _13464_ (.A(net43),
    .B(_05517_),
    .Y(_05677_));
 sky130_fd_sc_hd__and3_1 _13465_ (.A(net42),
    .B(_05520_),
    .C(_05521_),
    .X(_05678_));
 sky130_fd_sc_hd__and3_1 _13466_ (.A(net39),
    .B(_05523_),
    .C(_05524_),
    .X(_05679_));
 sky130_fd_sc_hd__xor2_1 _13467_ (.A(_05678_),
    .B(_05679_),
    .X(_05680_));
 sky130_fd_sc_hd__xnor2_2 _13468_ (.A(_05677_),
    .B(_05680_),
    .Y(_05681_));
 sky130_fd_sc_hd__and2_1 _13469_ (.A(_05483_),
    .B(_05485_),
    .X(_05682_));
 sky130_fd_sc_hd__clkbuf_4 _13470_ (.A(_05682_),
    .X(_05683_));
 sky130_fd_sc_hd__a31o_1 _13471_ (.A1(net35),
    .A2(_05683_),
    .A3(_05503_),
    .B1(_05505_),
    .X(_05684_));
 sky130_fd_sc_hd__o21a_1 _13472_ (.A1(_05502_),
    .A2(_05503_),
    .B1(_05684_),
    .X(_05685_));
 sky130_fd_sc_hd__nand2_1 _13473_ (.A(net32),
    .B(_05683_),
    .Y(_05686_));
 sky130_fd_sc_hd__and3_1 _13474_ (.A(net35),
    .B(_05488_),
    .C(_05490_),
    .X(_05687_));
 sky130_fd_sc_hd__inv_1 _13475_ (.A(net38),
    .Y(_05688_));
 sky130_fd_sc_hd__nor3_1 _13476_ (.A(_05688_),
    .B(_05493_),
    .C(_05494_),
    .Y(_05689_));
 sky130_fd_sc_hd__xor2_1 _13477_ (.A(_05687_),
    .B(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__xnor2_2 _13478_ (.A(_05686_),
    .B(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hd__xnor2_1 _13479_ (.A(_05685_),
    .B(_05691_),
    .Y(_05692_));
 sky130_fd_sc_hd__xnor2_2 _13480_ (.A(_05681_),
    .B(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__a21o_1 _13481_ (.A1(_05499_),
    .A2(_05507_),
    .B1(_05482_),
    .X(_05694_));
 sky130_fd_sc_hd__o21a_1 _13482_ (.A1(_05499_),
    .A2(_05507_),
    .B1(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__nand2_1 _13483_ (.A(net45),
    .B(_05585_),
    .Y(_05696_));
 sky130_fd_sc_hd__nor3_1 _13484_ (.A(_05541_),
    .B(_05538_),
    .C(_05539_),
    .Y(_05697_));
 sky130_fd_sc_hd__or3_1 _13485_ (.A(_05530_),
    .B(_05543_),
    .C(_05545_),
    .X(_05698_));
 sky130_fd_sc_hd__xor2_1 _13486_ (.A(_05697_),
    .B(_05698_),
    .X(_05699_));
 sky130_fd_sc_hd__xor2_2 _13487_ (.A(_05696_),
    .B(_05699_),
    .X(_05700_));
 sky130_fd_sc_hd__nor2_1 _13488_ (.A(_05477_),
    .B(_05480_),
    .Y(_05701_));
 sky130_fd_sc_hd__nand2_1 _13489_ (.A(_05477_),
    .B(_05480_),
    .Y(_05702_));
 sky130_fd_sc_hd__o21ai_2 _13490_ (.A1(_05701_),
    .A2(_05473_),
    .B1(_05702_),
    .Y(_05703_));
 sky130_fd_sc_hd__and2_1 _13491_ (.A(net52),
    .B(_05587_),
    .X(_05704_));
 sky130_fd_sc_hd__a41o_1 _13492_ (.A1(net52),
    .A2(net49),
    .A3(_05585_),
    .A4(_05587_),
    .B1(_05540_),
    .X(_05705_));
 sky130_fd_sc_hd__o21a_1 _13493_ (.A1(_05535_),
    .A2(_05704_),
    .B1(_05705_),
    .X(_05706_));
 sky130_fd_sc_hd__xnor2_1 _13494_ (.A(_05703_),
    .B(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__xnor2_1 _13495_ (.A(_05700_),
    .B(_05707_),
    .Y(_05708_));
 sky130_fd_sc_hd__xnor2_1 _13496_ (.A(_05695_),
    .B(_05708_),
    .Y(_05709_));
 sky130_fd_sc_hd__xnor2_2 _13497_ (.A(_05693_),
    .B(_05709_),
    .Y(_05710_));
 sky130_fd_sc_hd__o21ba_1 _13498_ (.A1(_05509_),
    .A2(_05529_),
    .B1_N(_05557_),
    .X(_05711_));
 sky130_fd_sc_hd__a21o_1 _13499_ (.A1(_05509_),
    .A2(_05529_),
    .B1(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__xnor2_1 _13500_ (.A(_05710_),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__xnor2_1 _13501_ (.A(_05676_),
    .B(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__a21bo_1 _13502_ (.A1(_05649_),
    .A2(_05651_),
    .B1_N(_05714_),
    .X(_05715_));
 sky130_fd_sc_hd__o21a_1 _13503_ (.A1(_05649_),
    .A2(_05651_),
    .B1(_05715_),
    .X(_05716_));
 sky130_fd_sc_hd__buf_6 _13504_ (.A(_05474_),
    .X(_05717_));
 sky130_fd_sc_hd__and3_1 _13505_ (.A(\top0.matmul0.alpha_pass[14] ),
    .B(_05436_),
    .C(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__buf_6 _13506_ (.A(_05470_),
    .X(_05719_));
 sky130_fd_sc_hd__a32o_1 _13507_ (.A1(\top0.matmul0.beta_pass[14] ),
    .A2(_05436_),
    .A3(_05719_),
    .B1(_05464_),
    .B2(\top0.c_out_calc[14] ),
    .X(_05720_));
 sky130_fd_sc_hd__nor2_4 _13508_ (.A(_05718_),
    .B(_05720_),
    .Y(_05721_));
 sky130_fd_sc_hd__nand2_1 _13509_ (.A(\top0.periodTop_r[0] ),
    .B(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__clkbuf_4 _13510_ (.A(_05616_),
    .X(_05723_));
 sky130_fd_sc_hd__clkbuf_4 _13511_ (.A(_05617_),
    .X(_05724_));
 sky130_fd_sc_hd__and3_1 _13512_ (.A(net60),
    .B(_05723_),
    .C(_05724_),
    .X(_05725_));
 sky130_fd_sc_hd__clkbuf_4 _13513_ (.A(_05663_),
    .X(_05726_));
 sky130_fd_sc_hd__clkbuf_4 _13514_ (.A(_05664_),
    .X(_05727_));
 sky130_fd_sc_hd__and3_1 _13515_ (.A(net64),
    .B(_05726_),
    .C(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__xnor2_1 _13516_ (.A(_05725_),
    .B(_05728_),
    .Y(_05729_));
 sky130_fd_sc_hd__xnor2_2 _13517_ (.A(_05722_),
    .B(_05729_),
    .Y(_05730_));
 sky130_fd_sc_hd__nand2_4 _13518_ (.A(_05611_),
    .B(_05612_),
    .Y(_05731_));
 sky130_fd_sc_hd__nor2_1 _13519_ (.A(_05536_),
    .B(_05731_),
    .Y(_05732_));
 sky130_fd_sc_hd__a32o_1 _13520_ (.A1(net1025),
    .A2(_05656_),
    .A3(_05639_),
    .B1(_05624_),
    .B2(net60),
    .X(_05733_));
 sky130_fd_sc_hd__o21a_1 _13521_ (.A1(_05656_),
    .A2(_05732_),
    .B1(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__inv_2 _13522_ (.A(net57),
    .Y(_05735_));
 sky130_fd_sc_hd__nor2_1 _13523_ (.A(_05735_),
    .B(_05629_),
    .Y(_05736_));
 sky130_fd_sc_hd__and3_1 _13524_ (.A(net1025),
    .B(_05602_),
    .C(_05603_),
    .X(_05737_));
 sky130_fd_sc_hd__or3_1 _13525_ (.A(_05541_),
    .B(_05637_),
    .C(_05638_),
    .X(_05738_));
 sky130_fd_sc_hd__xor2_1 _13526_ (.A(_05737_),
    .B(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__xnor2_2 _13527_ (.A(_05736_),
    .B(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__xnor2_1 _13528_ (.A(_05734_),
    .B(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__xnor2_2 _13529_ (.A(_05730_),
    .B(_05741_),
    .Y(_05742_));
 sky130_fd_sc_hd__nor2_1 _13530_ (.A(_05700_),
    .B(_05703_),
    .Y(_05743_));
 sky130_fd_sc_hd__a21oi_1 _13531_ (.A1(_05700_),
    .A2(_05703_),
    .B1(_05706_),
    .Y(_05744_));
 sky130_fd_sc_hd__o21ai_2 _13532_ (.A1(_05672_),
    .A2(_05661_),
    .B1(_05669_),
    .Y(_05745_));
 sky130_fd_sc_hd__nand2_1 _13533_ (.A(_05672_),
    .B(_05661_),
    .Y(_05746_));
 sky130_fd_sc_hd__a2bb2o_1 _13534_ (.A1_N(_05743_),
    .A2_N(_05744_),
    .B1(_05745_),
    .B2(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__nand4bb_2 _13535_ (.A_N(_05743_),
    .B_N(_05744_),
    .C(_05745_),
    .D(_05746_),
    .Y(_05748_));
 sky130_fd_sc_hd__and3_1 _13536_ (.A(_05742_),
    .B(_05747_),
    .C(_05748_),
    .X(_05749_));
 sky130_fd_sc_hd__a21oi_1 _13537_ (.A1(_05747_),
    .A2(_05748_),
    .B1(_05742_),
    .Y(_05750_));
 sky130_fd_sc_hd__or2_1 _13538_ (.A(_05749_),
    .B(_05750_),
    .X(_05751_));
 sky130_fd_sc_hd__a21o_1 _13539_ (.A1(_05708_),
    .A2(_05693_),
    .B1(_05695_),
    .X(_05752_));
 sky130_fd_sc_hd__or2_1 _13540_ (.A(_05708_),
    .B(_05693_),
    .X(_05753_));
 sky130_fd_sc_hd__nand3b_1 _13541_ (.A_N(_05751_),
    .B(_05752_),
    .C(_05753_),
    .Y(_05754_));
 sky130_fd_sc_hd__a21bo_1 _13542_ (.A1(_05752_),
    .A2(_05753_),
    .B1_N(_05751_),
    .X(_05755_));
 sky130_fd_sc_hd__and3_2 _13543_ (.A(net1030),
    .B(_05484_),
    .C(_05486_),
    .X(_05756_));
 sky130_fd_sc_hd__and3_2 _13544_ (.A(net32),
    .B(_05488_),
    .C(_05490_),
    .X(_05757_));
 sky130_fd_sc_hd__or3_1 _13545_ (.A(_05500_),
    .B(_05493_),
    .C(_05494_),
    .X(_05758_));
 sky130_fd_sc_hd__xor2_2 _13546_ (.A(_05757_),
    .B(_05758_),
    .X(_05759_));
 sky130_fd_sc_hd__xnor2_4 _13547_ (.A(_05756_),
    .B(_05759_),
    .Y(_05760_));
 sky130_fd_sc_hd__a21o_1 _13548_ (.A1(net32),
    .A2(_05682_),
    .B1(_05687_),
    .X(_05761_));
 sky130_fd_sc_hd__and3_1 _13549_ (.A(net32),
    .B(_05682_),
    .C(_05687_),
    .X(_05762_));
 sky130_fd_sc_hd__a21o_1 _13550_ (.A1(_05689_),
    .A2(_05761_),
    .B1(_05762_),
    .X(_05763_));
 sky130_fd_sc_hd__nand2_1 _13551_ (.A(net42),
    .B(_05472_),
    .Y(_05764_));
 sky130_fd_sc_hd__and3_1 _13552_ (.A(net37),
    .B(_05478_),
    .C(_05479_),
    .X(_05765_));
 sky130_fd_sc_hd__and3_1 _13553_ (.A(net39),
    .B(_05475_),
    .C(_05476_),
    .X(_05766_));
 sky130_fd_sc_hd__xor2_1 _13554_ (.A(_05765_),
    .B(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__xnor2_2 _13555_ (.A(_05764_),
    .B(_05767_),
    .Y(_05768_));
 sky130_fd_sc_hd__xnor2_2 _13556_ (.A(_05763_),
    .B(_05768_),
    .Y(_05769_));
 sky130_fd_sc_hd__xnor2_4 _13557_ (.A(_05760_),
    .B(_05769_),
    .Y(_05770_));
 sky130_fd_sc_hd__a21o_1 _13558_ (.A1(_05685_),
    .A2(_05691_),
    .B1(_05681_),
    .X(_05771_));
 sky130_fd_sc_hd__o21a_2 _13559_ (.A1(_05685_),
    .A2(_05691_),
    .B1(_05771_),
    .X(_05772_));
 sky130_fd_sc_hd__nand2_1 _13560_ (.A(net44),
    .B(_05586_),
    .Y(_05773_));
 sky130_fd_sc_hd__nor3_1 _13561_ (.A(_05530_),
    .B(_05538_),
    .C(_05539_),
    .Y(_05774_));
 sky130_fd_sc_hd__or3_1 _13562_ (.A(_05573_),
    .B(_05542_),
    .C(_05544_),
    .X(_05775_));
 sky130_fd_sc_hd__xnor2_1 _13563_ (.A(_05774_),
    .B(_05775_),
    .Y(_05776_));
 sky130_fd_sc_hd__xnor2_2 _13564_ (.A(_05773_),
    .B(_05776_),
    .Y(_05777_));
 sky130_fd_sc_hd__a41o_1 _13565_ (.A1(net49),
    .A2(net46),
    .A3(_05585_),
    .A4(_05587_),
    .B1(_05697_),
    .X(_05778_));
 sky130_fd_sc_hd__a21bo_1 _13566_ (.A1(_05696_),
    .A2(_05698_),
    .B1_N(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__a22o_1 _13567_ (.A1(net43),
    .A2(_05472_),
    .B1(_05678_),
    .B2(_05679_),
    .X(_05780_));
 sky130_fd_sc_hd__o21ai_2 _13568_ (.A1(_05678_),
    .A2(_05679_),
    .B1(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__xnor2_1 _13569_ (.A(_05779_),
    .B(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__xnor2_2 _13570_ (.A(_05777_),
    .B(_05782_),
    .Y(_05783_));
 sky130_fd_sc_hd__xnor2_1 _13571_ (.A(_05772_),
    .B(_05783_),
    .Y(_05784_));
 sky130_fd_sc_hd__xnor2_2 _13572_ (.A(_05770_),
    .B(_05784_),
    .Y(_05785_));
 sky130_fd_sc_hd__a21oi_1 _13573_ (.A1(_05754_),
    .A2(_05755_),
    .B1(_05785_),
    .Y(_05786_));
 sky130_fd_sc_hd__and3_1 _13574_ (.A(_05785_),
    .B(_05754_),
    .C(_05755_),
    .X(_05787_));
 sky130_fd_sc_hd__nor2_1 _13575_ (.A(_05786_),
    .B(_05787_),
    .Y(_05788_));
 sky130_fd_sc_hd__o21a_1 _13576_ (.A1(_05710_),
    .A2(_05712_),
    .B1(_05676_),
    .X(_05789_));
 sky130_fd_sc_hd__nand4_2 _13577_ (.A(net66),
    .B(net63),
    .C(_05619_),
    .D(_05666_),
    .Y(_05790_));
 sky130_fd_sc_hd__o21ba_1 _13578_ (.A1(_05653_),
    .A2(_05655_),
    .B1_N(_05674_),
    .X(_05791_));
 sky130_fd_sc_hd__a21o_1 _13579_ (.A1(_05653_),
    .A2(_05655_),
    .B1(_05791_),
    .X(_05792_));
 sky130_fd_sc_hd__xor2_1 _13580_ (.A(_05790_),
    .B(_05792_),
    .X(_05793_));
 sky130_fd_sc_hd__a21o_1 _13581_ (.A1(_05710_),
    .A2(_05712_),
    .B1(_05793_),
    .X(_05794_));
 sky130_fd_sc_hd__and2_1 _13582_ (.A(_05710_),
    .B(_05712_),
    .X(_05795_));
 sky130_fd_sc_hd__o21a_1 _13583_ (.A1(_05795_),
    .A2(_05789_),
    .B1(_05793_),
    .X(_05796_));
 sky130_fd_sc_hd__o21bai_1 _13584_ (.A1(_05789_),
    .A2(_05794_),
    .B1_N(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__xnor2_1 _13585_ (.A(_05788_),
    .B(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__or2_1 _13586_ (.A(_05716_),
    .B(_05798_),
    .X(_05799_));
 sky130_fd_sc_hd__xnor2_1 _13587_ (.A(_05651_),
    .B(_05714_),
    .Y(_05800_));
 sky130_fd_sc_hd__xnor2_1 _13588_ (.A(_05649_),
    .B(_05800_),
    .Y(_05801_));
 sky130_fd_sc_hd__xor2_1 _13589_ (.A(_05559_),
    .B(_05598_),
    .X(_05802_));
 sky130_fd_sc_hd__xnor2_1 _13590_ (.A(_05647_),
    .B(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__o22a_1 _13591_ (.A1(_05626_),
    .A2(_05639_),
    .B1(_05622_),
    .B2(net66),
    .X(_05804_));
 sky130_fd_sc_hd__inv_2 _13592_ (.A(net65),
    .Y(_05805_));
 sky130_fd_sc_hd__and3_1 _13593_ (.A(_05805_),
    .B(net61),
    .C(_05621_),
    .X(_05806_));
 sky130_fd_sc_hd__a211o_1 _13594_ (.A1(net66),
    .A2(_05641_),
    .B1(_05806_),
    .C1(_05731_),
    .X(_05807_));
 sky130_fd_sc_hd__a31o_1 _13595_ (.A1(net66),
    .A2(_05626_),
    .A3(_05621_),
    .B1(_05640_),
    .X(_05808_));
 sky130_fd_sc_hd__a2bb2oi_4 _13596_ (.A1_N(_05621_),
    .A2_N(_05804_),
    .B1(_05807_),
    .B2(_05808_),
    .Y(_05809_));
 sky130_fd_sc_hd__nand2_1 _13597_ (.A(net63),
    .B(_05551_),
    .Y(_05810_));
 sky130_fd_sc_hd__or3_2 _13598_ (.A(_05657_),
    .B(_05543_),
    .C(_05545_),
    .X(_05811_));
 sky130_fd_sc_hd__or3_2 _13599_ (.A(_05735_),
    .B(_05531_),
    .C(_05532_),
    .X(_05812_));
 sky130_fd_sc_hd__or2_1 _13600_ (.A(_05811_),
    .B(_05812_),
    .X(_05813_));
 sky130_fd_sc_hd__nand2_1 _13601_ (.A(_05811_),
    .B(_05812_),
    .Y(_05814_));
 sky130_fd_sc_hd__a21bo_1 _13602_ (.A1(_05810_),
    .A2(_05813_),
    .B1_N(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__and3_1 _13603_ (.A(net1027),
    .B(_05520_),
    .C(_05521_),
    .X(_05816_));
 sky130_fd_sc_hd__and3_1 _13604_ (.A(net50),
    .B(_05523_),
    .C(_05524_),
    .X(_05817_));
 sky130_fd_sc_hd__nor2_1 _13605_ (.A(_05816_),
    .B(_05817_),
    .Y(_05818_));
 sky130_fd_sc_hd__nand2_1 _13606_ (.A(\top0.periodTop_r[4] ),
    .B(_05517_),
    .Y(_05819_));
 sky130_fd_sc_hd__nand2_1 _13607_ (.A(_05816_),
    .B(_05817_),
    .Y(_05820_));
 sky130_fd_sc_hd__o21a_1 _13608_ (.A1(_05818_),
    .A2(_05819_),
    .B1(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__buf_6 _13609_ (.A(_05534_),
    .X(_05822_));
 sky130_fd_sc_hd__o211ai_1 _13610_ (.A1(_05536_),
    .A2(_05822_),
    .B1(_05588_),
    .C1(net56),
    .Y(_05823_));
 sky130_fd_sc_hd__a211o_1 _13611_ (.A1(net57),
    .A2(_05588_),
    .B1(_05822_),
    .C1(_05536_),
    .X(_05824_));
 sky130_fd_sc_hd__nand2_1 _13612_ (.A(_05823_),
    .B(_05824_),
    .Y(_05825_));
 sky130_fd_sc_hd__xnor2_2 _13613_ (.A(_05590_),
    .B(_05825_),
    .Y(_05826_));
 sky130_fd_sc_hd__a21o_1 _13614_ (.A1(_05815_),
    .A2(_05821_),
    .B1(_05826_),
    .X(_05827_));
 sky130_fd_sc_hd__o21ai_2 _13615_ (.A1(_05815_),
    .A2(_05821_),
    .B1(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__xor2_2 _13616_ (.A(_05578_),
    .B(_05594_),
    .X(_05829_));
 sky130_fd_sc_hd__xnor2_4 _13617_ (.A(_05596_),
    .B(_05829_),
    .Y(_05830_));
 sky130_fd_sc_hd__xor2_1 _13618_ (.A(_05815_),
    .B(_05821_),
    .X(_05831_));
 sky130_fd_sc_hd__xnor2_2 _13619_ (.A(_05826_),
    .B(_05831_),
    .Y(_05832_));
 sky130_fd_sc_hd__xnor2_1 _13620_ (.A(_05571_),
    .B(_05572_),
    .Y(_05833_));
 sky130_fd_sc_hd__nand2_1 _13621_ (.A(_05574_),
    .B(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__or2_1 _13622_ (.A(_05574_),
    .B(_05833_),
    .X(_05835_));
 sky130_fd_sc_hd__xnor2_1 _13623_ (.A(_05816_),
    .B(_05817_),
    .Y(_05836_));
 sky130_fd_sc_hd__xnor2_1 _13624_ (.A(_05819_),
    .B(_05836_),
    .Y(_05837_));
 sky130_fd_sc_hd__and3_1 _13625_ (.A(_05834_),
    .B(_05835_),
    .C(_05837_),
    .X(_05838_));
 sky130_fd_sc_hd__and3_1 _13626_ (.A(net47),
    .B(_05489_),
    .C(_05491_),
    .X(_05839_));
 sky130_fd_sc_hd__and3_1 _13627_ (.A(net43),
    .B(_05484_),
    .C(_05486_),
    .X(_05840_));
 sky130_fd_sc_hd__o211a_1 _13628_ (.A1(_05839_),
    .A2(_05840_),
    .B1(net50),
    .C1(_05496_),
    .X(_05841_));
 sky130_fd_sc_hd__a21oi_1 _13629_ (.A1(_05839_),
    .A2(_05840_),
    .B1(_05841_),
    .Y(_05842_));
 sky130_fd_sc_hd__a21o_1 _13630_ (.A1(_05834_),
    .A2(_05835_),
    .B1(_05837_),
    .X(_05843_));
 sky130_fd_sc_hd__o21ai_2 _13631_ (.A1(_05838_),
    .A2(_05842_),
    .B1(_05843_),
    .Y(_05844_));
 sky130_fd_sc_hd__xor2_1 _13632_ (.A(_05564_),
    .B(_05570_),
    .X(_05845_));
 sky130_fd_sc_hd__xnor2_1 _13633_ (.A(_05576_),
    .B(_05845_),
    .Y(_05846_));
 sky130_fd_sc_hd__o21a_1 _13634_ (.A1(_05832_),
    .A2(_05844_),
    .B1(_05846_),
    .X(_05847_));
 sky130_fd_sc_hd__a21oi_2 _13635_ (.A1(_05832_),
    .A2(_05844_),
    .B1(_05847_),
    .Y(_05848_));
 sky130_fd_sc_hd__nand2_1 _13636_ (.A(_05830_),
    .B(_05848_),
    .Y(_05849_));
 sky130_fd_sc_hd__or2_1 _13637_ (.A(_05828_),
    .B(_05849_),
    .X(_05850_));
 sky130_fd_sc_hd__nor2_1 _13638_ (.A(_05830_),
    .B(_05848_),
    .Y(_05851_));
 sky130_fd_sc_hd__o21a_1 _13639_ (.A1(_05828_),
    .A2(_05851_),
    .B1(_05849_),
    .X(_05852_));
 sky130_fd_sc_hd__a21o_1 _13640_ (.A1(_05809_),
    .A2(_05850_),
    .B1(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__nand3_1 _13641_ (.A(_05828_),
    .B(_05809_),
    .C(_05851_),
    .Y(_05854_));
 sky130_fd_sc_hd__a21bo_1 _13642_ (.A1(_05803_),
    .A2(_05853_),
    .B1_N(_05854_),
    .X(_05855_));
 sky130_fd_sc_hd__nand2_1 _13643_ (.A(_05801_),
    .B(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__and2_1 _13644_ (.A(_05716_),
    .B(_05798_),
    .X(_05857_));
 sky130_fd_sc_hd__a21o_1 _13645_ (.A1(_05799_),
    .A2(_05856_),
    .B1(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__o211a_1 _13646_ (.A1(_05809_),
    .A2(_05852_),
    .B1(_05850_),
    .C1(_05854_),
    .X(_05859_));
 sky130_fd_sc_hd__xnor2_1 _13647_ (.A(_05803_),
    .B(_05859_),
    .Y(_05860_));
 sky130_fd_sc_hd__nand2_1 _13648_ (.A(\top0.periodTop_r[1] ),
    .B(_05640_),
    .Y(_05861_));
 sky130_fd_sc_hd__nand2_1 _13649_ (.A(net66),
    .B(_05605_),
    .Y(_05862_));
 sky130_fd_sc_hd__xnor2_2 _13650_ (.A(_05861_),
    .B(_05862_),
    .Y(_05863_));
 sky130_fd_sc_hd__xor2_1 _13651_ (.A(_05811_),
    .B(_05812_),
    .X(_05864_));
 sky130_fd_sc_hd__xnor2_2 _13652_ (.A(_05810_),
    .B(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__a22o_1 _13653_ (.A1(net61),
    .A2(_05585_),
    .B1(_05588_),
    .B2(net63),
    .X(_05866_));
 sky130_fd_sc_hd__and4_1 _13654_ (.A(net63),
    .B(net61),
    .C(_05585_),
    .D(_05587_),
    .X(_05867_));
 sky130_fd_sc_hd__a31o_1 _13655_ (.A1(net67),
    .A2(_05551_),
    .A3(_05866_),
    .B1(_05867_),
    .X(_05868_));
 sky130_fd_sc_hd__and3_1 _13656_ (.A(net54),
    .B(_05520_),
    .C(_05521_),
    .X(_05869_));
 sky130_fd_sc_hd__and3_1 _13657_ (.A(net1027),
    .B(_05478_),
    .C(_05479_),
    .X(_05870_));
 sky130_fd_sc_hd__o211a_1 _13658_ (.A1(_05869_),
    .A2(_05870_),
    .B1(net57),
    .C1(_05472_),
    .X(_05871_));
 sky130_fd_sc_hd__a21o_1 _13659_ (.A1(_05869_),
    .A2(_05870_),
    .B1(_05871_),
    .X(_05872_));
 sky130_fd_sc_hd__o21a_1 _13660_ (.A1(_05865_),
    .A2(_05868_),
    .B1(_05872_),
    .X(_05873_));
 sky130_fd_sc_hd__a21oi_2 _13661_ (.A1(_05865_),
    .A2(_05868_),
    .B1(_05873_),
    .Y(_05874_));
 sky130_fd_sc_hd__nor2_1 _13662_ (.A(_05863_),
    .B(_05874_),
    .Y(_05875_));
 sky130_fd_sc_hd__xor2_1 _13663_ (.A(_05828_),
    .B(_05809_),
    .X(_05876_));
 sky130_fd_sc_hd__xnor2_2 _13664_ (.A(_05848_),
    .B(_05876_),
    .Y(_05877_));
 sky130_fd_sc_hd__xnor2_4 _13665_ (.A(_05830_),
    .B(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__or2_1 _13666_ (.A(_05863_),
    .B(_05874_),
    .X(_05879_));
 sky130_fd_sc_hd__nand2_1 _13667_ (.A(_05863_),
    .B(_05874_),
    .Y(_05880_));
 sky130_fd_sc_hd__and2_1 _13668_ (.A(_05879_),
    .B(_05880_),
    .X(_05881_));
 sky130_fd_sc_hd__xnor2_1 _13669_ (.A(_05832_),
    .B(_05844_),
    .Y(_05882_));
 sky130_fd_sc_hd__xnor2_1 _13670_ (.A(_05846_),
    .B(_05882_),
    .Y(_05883_));
 sky130_fd_sc_hd__nand2_1 _13671_ (.A(_05834_),
    .B(_05835_),
    .Y(_05884_));
 sky130_fd_sc_hd__xnor2_1 _13672_ (.A(_05837_),
    .B(_05842_),
    .Y(_05885_));
 sky130_fd_sc_hd__xnor2_2 _13673_ (.A(_05884_),
    .B(_05885_),
    .Y(_05886_));
 sky130_fd_sc_hd__nand2_1 _13674_ (.A(net50),
    .B(_05496_),
    .Y(_05887_));
 sky130_fd_sc_hd__xor2_1 _13675_ (.A(_05839_),
    .B(_05840_),
    .X(_05888_));
 sky130_fd_sc_hd__xnor2_2 _13676_ (.A(_05887_),
    .B(_05888_),
    .Y(_05889_));
 sky130_fd_sc_hd__nand2_1 _13677_ (.A(net58),
    .B(_05517_),
    .Y(_05890_));
 sky130_fd_sc_hd__xor2_2 _13678_ (.A(_05869_),
    .B(_05870_),
    .X(_05891_));
 sky130_fd_sc_hd__xnor2_2 _13679_ (.A(_05890_),
    .B(_05891_),
    .Y(_05892_));
 sky130_fd_sc_hd__and2_1 _13680_ (.A(_05488_),
    .B(_05490_),
    .X(_05893_));
 sky130_fd_sc_hd__buf_2 _13681_ (.A(_05893_),
    .X(_05894_));
 sky130_fd_sc_hd__a22o_1 _13682_ (.A1(net47),
    .A2(_05682_),
    .B1(_05894_),
    .B2(net50),
    .X(_05895_));
 sky130_fd_sc_hd__and4_1 _13683_ (.A(net50),
    .B(net47),
    .C(_05682_),
    .D(_05894_),
    .X(_05896_));
 sky130_fd_sc_hd__a31o_1 _13684_ (.A1(net1027),
    .A2(_05497_),
    .A3(_05895_),
    .B1(_05896_),
    .X(_05897_));
 sky130_fd_sc_hd__o21a_1 _13685_ (.A1(_05889_),
    .A2(_05892_),
    .B1(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__a21o_1 _13686_ (.A1(_05889_),
    .A2(_05892_),
    .B1(_05898_),
    .X(_05899_));
 sky130_fd_sc_hd__xor2_1 _13687_ (.A(_05872_),
    .B(_05868_),
    .X(_05900_));
 sky130_fd_sc_hd__xnor2_2 _13688_ (.A(_05865_),
    .B(_05900_),
    .Y(_05901_));
 sky130_fd_sc_hd__a21bo_1 _13689_ (.A1(_05886_),
    .A2(_05899_),
    .B1_N(_05901_),
    .X(_05902_));
 sky130_fd_sc_hd__o21a_1 _13690_ (.A1(_05886_),
    .A2(_05899_),
    .B1(_05902_),
    .X(_05903_));
 sky130_fd_sc_hd__or2_1 _13691_ (.A(_05883_),
    .B(_05903_),
    .X(_05904_));
 sky130_fd_sc_hd__nand2_1 _13692_ (.A(_05883_),
    .B(_05903_),
    .Y(_05905_));
 sky130_fd_sc_hd__a21bo_1 _13693_ (.A1(_05881_),
    .A2(_05904_),
    .B1_N(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__o21a_1 _13694_ (.A1(_05875_),
    .A2(_05878_),
    .B1(_05906_),
    .X(_05907_));
 sky130_fd_sc_hd__a21oi_1 _13695_ (.A1(_05875_),
    .A2(_05878_),
    .B1(_05907_),
    .Y(_05908_));
 sky130_fd_sc_hd__nor2_1 _13696_ (.A(_05805_),
    .B(_05731_),
    .Y(_05909_));
 sky130_fd_sc_hd__and3_1 _13697_ (.A(net57),
    .B(_05475_),
    .C(_05476_),
    .X(_05910_));
 sky130_fd_sc_hd__and3_1 _13698_ (.A(net54),
    .B(_05478_),
    .C(_05479_),
    .X(_05911_));
 sky130_fd_sc_hd__o211a_1 _13699_ (.A1(_05910_),
    .A2(_05911_),
    .B1(net59),
    .C1(_05517_),
    .X(_05912_));
 sky130_fd_sc_hd__a21o_1 _13700_ (.A1(_05910_),
    .A2(_05911_),
    .B1(_05912_),
    .X(_05913_));
 sky130_fd_sc_hd__nand2_1 _13701_ (.A(net67),
    .B(_05579_),
    .Y(_05914_));
 sky130_fd_sc_hd__o211a_1 _13702_ (.A1(_05657_),
    .A2(_05822_),
    .B1(_05588_),
    .C1(net64),
    .X(_05915_));
 sky130_fd_sc_hd__o311a_1 _13703_ (.A1(_05607_),
    .A2(_05543_),
    .A3(_05545_),
    .B1(net61),
    .C1(_05585_),
    .X(_05916_));
 sky130_fd_sc_hd__or2_1 _13704_ (.A(_05915_),
    .B(_05916_),
    .X(_05917_));
 sky130_fd_sc_hd__xnor2_2 _13705_ (.A(_05914_),
    .B(_05917_),
    .Y(_05918_));
 sky130_fd_sc_hd__and4_1 _13706_ (.A(net67),
    .B(net63),
    .C(_05586_),
    .D(_05588_),
    .X(_05919_));
 sky130_fd_sc_hd__o21a_1 _13707_ (.A1(_05913_),
    .A2(_05918_),
    .B1(_05919_),
    .X(_05920_));
 sky130_fd_sc_hd__a21o_1 _13708_ (.A1(_05913_),
    .A2(_05918_),
    .B1(_05920_),
    .X(_05921_));
 sky130_fd_sc_hd__nand2_1 _13709_ (.A(_05909_),
    .B(_05921_),
    .Y(_05922_));
 sky130_fd_sc_hd__or2_1 _13710_ (.A(_05909_),
    .B(_05921_),
    .X(_05923_));
 sky130_fd_sc_hd__nand2_1 _13711_ (.A(_05922_),
    .B(_05923_),
    .Y(_05924_));
 sky130_fd_sc_hd__xnor2_1 _13712_ (.A(_05901_),
    .B(_05899_),
    .Y(_05925_));
 sky130_fd_sc_hd__xnor2_2 _13713_ (.A(_05886_),
    .B(_05925_),
    .Y(_05926_));
 sky130_fd_sc_hd__xnor2_1 _13714_ (.A(_05913_),
    .B(_05919_),
    .Y(_05927_));
 sky130_fd_sc_hd__xnor2_2 _13715_ (.A(_05918_),
    .B(_05927_),
    .Y(_05928_));
 sky130_fd_sc_hd__nand2_1 _13716_ (.A(net59),
    .B(_05472_),
    .Y(_05929_));
 sky130_fd_sc_hd__xor2_1 _13717_ (.A(_05910_),
    .B(_05911_),
    .X(_05930_));
 sky130_fd_sc_hd__xnor2_1 _13718_ (.A(_05929_),
    .B(_05930_),
    .Y(_05931_));
 sky130_fd_sc_hd__and3_1 _13719_ (.A(net1027),
    .B(_05488_),
    .C(_05490_),
    .X(_05932_));
 sky130_fd_sc_hd__and3_1 _13720_ (.A(net50),
    .B(_05484_),
    .C(_05486_),
    .X(_05933_));
 sky130_fd_sc_hd__o211a_1 _13721_ (.A1(_05932_),
    .A2(_05933_),
    .B1(net54),
    .C1(_05495_),
    .X(_05934_));
 sky130_fd_sc_hd__a21o_1 _13722_ (.A1(_05932_),
    .A2(_05933_),
    .B1(_05934_),
    .X(_05935_));
 sky130_fd_sc_hd__or2_1 _13723_ (.A(_05931_),
    .B(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__nand2_1 _13724_ (.A(net1027),
    .B(_05496_),
    .Y(_05937_));
 sky130_fd_sc_hd__nand2_1 _13725_ (.A(net50),
    .B(_05894_),
    .Y(_05938_));
 sky130_fd_sc_hd__nand2_1 _13726_ (.A(net47),
    .B(_05683_),
    .Y(_05939_));
 sky130_fd_sc_hd__xor2_1 _13727_ (.A(_05938_),
    .B(_05939_),
    .X(_05940_));
 sky130_fd_sc_hd__xnor2_1 _13728_ (.A(_05937_),
    .B(_05940_),
    .Y(_05941_));
 sky130_fd_sc_hd__and2_1 _13729_ (.A(_05931_),
    .B(_05935_),
    .X(_05942_));
 sky130_fd_sc_hd__a21o_1 _13730_ (.A1(_05936_),
    .A2(_05941_),
    .B1(_05942_),
    .X(_05943_));
 sky130_fd_sc_hd__xnor2_1 _13731_ (.A(_05897_),
    .B(_05892_),
    .Y(_05944_));
 sky130_fd_sc_hd__xnor2_1 _13732_ (.A(_05889_),
    .B(_05944_),
    .Y(_05945_));
 sky130_fd_sc_hd__a21o_1 _13733_ (.A1(_05928_),
    .A2(_05943_),
    .B1(_05945_),
    .X(_05946_));
 sky130_fd_sc_hd__o21ai_1 _13734_ (.A1(_05928_),
    .A2(_05943_),
    .B1(_05946_),
    .Y(_05947_));
 sky130_fd_sc_hd__a21o_1 _13735_ (.A1(_05924_),
    .A2(_05926_),
    .B1(_05947_),
    .X(_05948_));
 sky130_fd_sc_hd__o21a_1 _13736_ (.A1(_05924_),
    .A2(_05926_),
    .B1(_05948_),
    .X(_05949_));
 sky130_fd_sc_hd__inv_2 _13737_ (.A(_05881_),
    .Y(_05950_));
 sky130_fd_sc_hd__mux2_1 _13738_ (.A0(_05905_),
    .A1(_05904_),
    .S(_05878_),
    .X(_05951_));
 sky130_fd_sc_hd__nand2_1 _13739_ (.A(_05905_),
    .B(_05904_),
    .Y(_05952_));
 sky130_fd_sc_hd__mux2_1 _13740_ (.A0(_05879_),
    .A1(_05880_),
    .S(_05878_),
    .X(_05953_));
 sky130_fd_sc_hd__o22a_1 _13741_ (.A1(_05950_),
    .A2(_05951_),
    .B1(_05952_),
    .B2(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__o22a_1 _13742_ (.A1(_05949_),
    .A2(_05954_),
    .B1(_05860_),
    .B2(_05908_),
    .X(_05955_));
 sky130_fd_sc_hd__nand2_1 _13743_ (.A(_05947_),
    .B(_05926_),
    .Y(_05956_));
 sky130_fd_sc_hd__or2_1 _13744_ (.A(_05947_),
    .B(_05926_),
    .X(_05957_));
 sky130_fd_sc_hd__nand2_1 _13745_ (.A(_05956_),
    .B(_05957_),
    .Y(_05958_));
 sky130_fd_sc_hd__xnor2_1 _13746_ (.A(_05924_),
    .B(_05958_),
    .Y(_05959_));
 sky130_fd_sc_hd__and2_1 _13747_ (.A(net62),
    .B(_05472_),
    .X(_05960_));
 sky130_fd_sc_hd__and3_1 _13748_ (.A(net59),
    .B(_05520_),
    .C(_05521_),
    .X(_05961_));
 sky130_fd_sc_hd__and3_1 _13749_ (.A(net58),
    .B(_05478_),
    .C(_05479_),
    .X(_05962_));
 sky130_fd_sc_hd__o21a_1 _13750_ (.A1(_05960_),
    .A2(_05961_),
    .B1(_05962_),
    .X(_05963_));
 sky130_fd_sc_hd__and3_1 _13751_ (.A(net62),
    .B(_05517_),
    .C(_05961_),
    .X(_05964_));
 sky130_fd_sc_hd__o211a_1 _13752_ (.A1(_05607_),
    .A2(_05534_),
    .B1(_05587_),
    .C1(net67),
    .X(_05965_));
 sky130_fd_sc_hd__a211o_1 _13753_ (.A1(net67),
    .A2(_05587_),
    .B1(_05534_),
    .C1(_05607_),
    .X(_05966_));
 sky130_fd_sc_hd__or2b_1 _13754_ (.A(_05965_),
    .B_N(_05966_),
    .X(_05967_));
 sky130_fd_sc_hd__o21ai_1 _13755_ (.A1(_05963_),
    .A2(_05964_),
    .B1(_05967_),
    .Y(_05968_));
 sky130_fd_sc_hd__or3_1 _13756_ (.A(_05967_),
    .B(_05963_),
    .C(_05964_),
    .X(_05969_));
 sky130_fd_sc_hd__nand2_1 _13757_ (.A(_05968_),
    .B(_05969_),
    .Y(_05970_));
 sky130_fd_sc_hd__nand2_1 _13758_ (.A(net54),
    .B(_05495_),
    .Y(_05971_));
 sky130_fd_sc_hd__xor2_1 _13759_ (.A(_05932_),
    .B(_05933_),
    .X(_05972_));
 sky130_fd_sc_hd__xnor2_2 _13760_ (.A(_05971_),
    .B(_05972_),
    .Y(_05973_));
 sky130_fd_sc_hd__and3_1 _13761_ (.A(net54),
    .B(_05489_),
    .C(_05491_),
    .X(_05974_));
 sky130_fd_sc_hd__and3_1 _13762_ (.A(net1027),
    .B(_05484_),
    .C(_05486_),
    .X(_05975_));
 sky130_fd_sc_hd__o211a_1 _13763_ (.A1(_05974_),
    .A2(_05975_),
    .B1(net58),
    .C1(_05495_),
    .X(_05976_));
 sky130_fd_sc_hd__a21o_1 _13764_ (.A1(_05974_),
    .A2(_05975_),
    .B1(_05976_),
    .X(_05977_));
 sky130_fd_sc_hd__xor2_1 _13765_ (.A(_05962_),
    .B(_05961_),
    .X(_05978_));
 sky130_fd_sc_hd__xnor2_2 _13766_ (.A(_05960_),
    .B(_05978_),
    .Y(_05979_));
 sky130_fd_sc_hd__a21bo_1 _13767_ (.A1(_05973_),
    .A2(_05977_),
    .B1_N(_05979_),
    .X(_05980_));
 sky130_fd_sc_hd__o21ai_2 _13768_ (.A1(_05973_),
    .A2(_05977_),
    .B1(_05980_),
    .Y(_05981_));
 sky130_fd_sc_hd__xor2_1 _13769_ (.A(_05931_),
    .B(_05935_),
    .X(_05982_));
 sky130_fd_sc_hd__xnor2_1 _13770_ (.A(_05941_),
    .B(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__a21o_1 _13771_ (.A1(_05970_),
    .A2(_05981_),
    .B1(_05983_),
    .X(_05984_));
 sky130_fd_sc_hd__or2_1 _13772_ (.A(_05968_),
    .B(_05984_),
    .X(_05985_));
 sky130_fd_sc_hd__xor2_1 _13773_ (.A(_05928_),
    .B(_05943_),
    .X(_05986_));
 sky130_fd_sc_hd__xnor2_1 _13774_ (.A(_05945_),
    .B(_05986_),
    .Y(_05987_));
 sky130_fd_sc_hd__inv_2 _13775_ (.A(_05969_),
    .Y(_05988_));
 sky130_fd_sc_hd__o211a_1 _13776_ (.A1(_05988_),
    .A2(_05981_),
    .B1(_05984_),
    .C1(_05968_),
    .X(_05989_));
 sky130_fd_sc_hd__a21o_1 _13777_ (.A1(_05985_),
    .A2(_05987_),
    .B1(_05989_),
    .X(_05990_));
 sky130_fd_sc_hd__inv_2 _13778_ (.A(_05985_),
    .Y(_05991_));
 sky130_fd_sc_hd__or3_1 _13779_ (.A(_05991_),
    .B(_05987_),
    .C(_05989_),
    .X(_05992_));
 sky130_fd_sc_hd__o21ai_1 _13780_ (.A1(_05991_),
    .A2(_05989_),
    .B1(_05987_),
    .Y(_05993_));
 sky130_fd_sc_hd__xor2_1 _13781_ (.A(_05973_),
    .B(_05977_),
    .X(_05994_));
 sky130_fd_sc_hd__xnor2_2 _13782_ (.A(_05979_),
    .B(_05994_),
    .Y(_05995_));
 sky130_fd_sc_hd__and3_1 _13783_ (.A(net58),
    .B(_05489_),
    .C(_05491_),
    .X(_05996_));
 sky130_fd_sc_hd__and3_1 _13784_ (.A(net54),
    .B(_05484_),
    .C(_05486_),
    .X(_05997_));
 sky130_fd_sc_hd__o211a_1 _13785_ (.A1(_05996_),
    .A2(_05997_),
    .B1(net59),
    .C1(_05496_),
    .X(_05998_));
 sky130_fd_sc_hd__a21o_1 _13786_ (.A1(_05996_),
    .A2(_05997_),
    .B1(_05998_),
    .X(_05999_));
 sky130_fd_sc_hd__nand2_1 _13787_ (.A(net58),
    .B(_05496_),
    .Y(_06000_));
 sky130_fd_sc_hd__xor2_1 _13788_ (.A(_05974_),
    .B(_05975_),
    .X(_06001_));
 sky130_fd_sc_hd__xnor2_2 _13789_ (.A(_06000_),
    .B(_06001_),
    .Y(_06002_));
 sky130_fd_sc_hd__nand2_1 _13790_ (.A(_05999_),
    .B(_06002_),
    .Y(_06003_));
 sky130_fd_sc_hd__nand2_1 _13791_ (.A(net68),
    .B(_05517_),
    .Y(_06004_));
 sky130_fd_sc_hd__and3_1 _13792_ (.A(\top0.periodTop_r[1] ),
    .B(_05520_),
    .C(_05521_),
    .X(_06005_));
 sky130_fd_sc_hd__and3_1 _13793_ (.A(\top0.periodTop_r[2] ),
    .B(_05523_),
    .C(_05524_),
    .X(_06006_));
 sky130_fd_sc_hd__xnor2_1 _13794_ (.A(_06005_),
    .B(_06006_),
    .Y(_06007_));
 sky130_fd_sc_hd__xnor2_1 _13795_ (.A(_06004_),
    .B(_06007_),
    .Y(_06008_));
 sky130_fd_sc_hd__o21bai_1 _13796_ (.A1(_05999_),
    .A2(_06002_),
    .B1_N(_06008_),
    .Y(_06009_));
 sky130_fd_sc_hd__and2_1 _13797_ (.A(_06005_),
    .B(_06006_),
    .X(_06010_));
 sky130_fd_sc_hd__o21a_1 _13798_ (.A1(_06005_),
    .A2(_06006_),
    .B1(_05517_),
    .X(_06011_));
 sky130_fd_sc_hd__o211ai_4 _13799_ (.A1(_06011_),
    .A2(_06010_),
    .B1(net68),
    .C1(_05586_),
    .Y(_06012_));
 sky130_fd_sc_hd__or3_1 _13800_ (.A(_05586_),
    .B(_06011_),
    .C(_06010_),
    .X(_06013_));
 sky130_fd_sc_hd__o211ai_2 _13801_ (.A1(net68),
    .A2(_06010_),
    .B1(_06012_),
    .C1(_06013_),
    .Y(_06014_));
 sky130_fd_sc_hd__nand3_1 _13802_ (.A(_06003_),
    .B(_06009_),
    .C(_06014_),
    .Y(_06015_));
 sky130_fd_sc_hd__a21o_1 _13803_ (.A1(_06003_),
    .A2(_06009_),
    .B1(_06014_),
    .X(_06016_));
 sky130_fd_sc_hd__a21bo_1 _13804_ (.A1(_05995_),
    .A2(_06015_),
    .B1_N(_06016_),
    .X(_06017_));
 sky130_fd_sc_hd__xor2_1 _13805_ (.A(_05983_),
    .B(_05970_),
    .X(_06018_));
 sky130_fd_sc_hd__xnor2_1 _13806_ (.A(_05981_),
    .B(_06018_),
    .Y(_06019_));
 sky130_fd_sc_hd__a21bo_1 _13807_ (.A1(_06003_),
    .A2(_06009_),
    .B1_N(_05995_),
    .X(_06020_));
 sky130_fd_sc_hd__and2b_1 _13808_ (.A_N(_06019_),
    .B(_06020_),
    .X(_06021_));
 sky130_fd_sc_hd__o2bb2a_1 _13809_ (.A1_N(_06017_),
    .A2_N(_06019_),
    .B1(_06021_),
    .B2(_06012_),
    .X(_06022_));
 sky130_fd_sc_hd__and2_1 _13810_ (.A(_05523_),
    .B(_05524_),
    .X(_06023_));
 sky130_fd_sc_hd__nand2_1 _13811_ (.A(net62),
    .B(_06023_),
    .Y(_06024_));
 sky130_fd_sc_hd__and2_2 _13812_ (.A(_05520_),
    .B(_05521_),
    .X(_06025_));
 sky130_fd_sc_hd__nand2_1 _13813_ (.A(net68),
    .B(_06025_),
    .Y(_06026_));
 sky130_fd_sc_hd__nand2_1 _13814_ (.A(net59),
    .B(_05496_),
    .Y(_06027_));
 sky130_fd_sc_hd__xor2_2 _13815_ (.A(_05996_),
    .B(_05997_),
    .X(_06028_));
 sky130_fd_sc_hd__xnor2_2 _13816_ (.A(_06027_),
    .B(_06028_),
    .Y(_06029_));
 sky130_fd_sc_hd__nand2_1 _13817_ (.A(net62),
    .B(_05496_),
    .Y(_06030_));
 sky130_fd_sc_hd__and3_1 _13818_ (.A(net59),
    .B(_05488_),
    .C(_05490_),
    .X(_06031_));
 sky130_fd_sc_hd__or3b_1 _13819_ (.A(_05735_),
    .B(_05501_),
    .C_N(_06031_),
    .X(_06032_));
 sky130_fd_sc_hd__a21oi_1 _13820_ (.A1(net58),
    .A2(_05683_),
    .B1(_06031_),
    .Y(_06033_));
 sky130_fd_sc_hd__a21oi_1 _13821_ (.A1(_06030_),
    .A2(_06032_),
    .B1(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__nand2_1 _13822_ (.A(_06029_),
    .B(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__or3_1 _13823_ (.A(_06024_),
    .B(_06026_),
    .C(_06035_),
    .X(_06036_));
 sky130_fd_sc_hd__and2_1 _13824_ (.A(_06016_),
    .B(_06015_),
    .X(_06037_));
 sky130_fd_sc_hd__xnor2_1 _13825_ (.A(_05995_),
    .B(_06037_),
    .Y(_06038_));
 sky130_fd_sc_hd__and3_1 _13826_ (.A(net62),
    .B(_05523_),
    .C(_05524_),
    .X(_06039_));
 sky130_fd_sc_hd__a311oi_1 _13827_ (.A1(net68),
    .A2(_06025_),
    .A3(_06039_),
    .B1(_06029_),
    .C1(_06034_),
    .Y(_06040_));
 sky130_fd_sc_hd__a31o_1 _13828_ (.A1(_06024_),
    .A2(_06026_),
    .A3(_06035_),
    .B1(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__xnor2_1 _13829_ (.A(_05999_),
    .B(_06008_),
    .Y(_06042_));
 sky130_fd_sc_hd__xnor2_1 _13830_ (.A(_06002_),
    .B(_06042_),
    .Y(_06043_));
 sky130_fd_sc_hd__o21a_1 _13831_ (.A1(_06041_),
    .A2(_06043_),
    .B1(_06036_),
    .X(_06044_));
 sky130_fd_sc_hd__xnor2_1 _13832_ (.A(net59),
    .B(_05497_),
    .Y(_06045_));
 sky130_fd_sc_hd__nand2_2 _13833_ (.A(_05489_),
    .B(_05491_),
    .Y(_06046_));
 sky130_fd_sc_hd__nor2_1 _13834_ (.A(_05501_),
    .B(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__and4_1 _13835_ (.A(net68),
    .B(net62),
    .C(_06023_),
    .D(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__a21oi_1 _13836_ (.A1(_05567_),
    .A2(_06032_),
    .B1(_06033_),
    .Y(_06049_));
 sky130_fd_sc_hd__o32a_1 _13837_ (.A1(_06023_),
    .A2(_06033_),
    .A3(_06030_),
    .B1(_06032_),
    .B2(_06039_),
    .X(_06050_));
 sky130_fd_sc_hd__o21a_1 _13838_ (.A1(_06024_),
    .A2(_06049_),
    .B1(_06050_),
    .X(_06051_));
 sky130_fd_sc_hd__xor2_1 _13839_ (.A(_06029_),
    .B(_06026_),
    .X(_06052_));
 sky130_fd_sc_hd__xnor2_1 _13840_ (.A(_06051_),
    .B(_06052_),
    .Y(_06053_));
 sky130_fd_sc_hd__a32o_1 _13841_ (.A1(net62),
    .A2(net59),
    .A3(_06047_),
    .B1(_05497_),
    .B2(net68),
    .X(_06054_));
 sky130_fd_sc_hd__a22o_1 _13842_ (.A1(net59),
    .A2(_05683_),
    .B1(_05894_),
    .B2(net62),
    .X(_06055_));
 sky130_fd_sc_hd__and2_1 _13843_ (.A(_06054_),
    .B(_06055_),
    .X(_06056_));
 sky130_fd_sc_hd__nand2_1 _13844_ (.A(net58),
    .B(_05683_),
    .Y(_06057_));
 sky130_fd_sc_hd__xnor2_1 _13845_ (.A(_06031_),
    .B(_06030_),
    .Y(_06058_));
 sky130_fd_sc_hd__xnor2_1 _13846_ (.A(_06057_),
    .B(_06058_),
    .Y(_06059_));
 sky130_fd_sc_hd__nand2_1 _13847_ (.A(_06056_),
    .B(_06059_),
    .Y(_06060_));
 sky130_fd_sc_hd__nand2_1 _13848_ (.A(_06053_),
    .B(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__a31o_1 _13849_ (.A1(net62),
    .A2(_06047_),
    .A3(_06045_),
    .B1(_06023_),
    .X(_06062_));
 sky130_fd_sc_hd__o211ai_1 _13850_ (.A1(_06056_),
    .A2(_06059_),
    .B1(_06062_),
    .C1(net68),
    .Y(_06063_));
 sky130_fd_sc_hd__a21oi_1 _13851_ (.A1(_06060_),
    .A2(_06063_),
    .B1(_06053_),
    .Y(_06064_));
 sky130_fd_sc_hd__a31o_1 _13852_ (.A1(_06045_),
    .A2(_06048_),
    .A3(_06061_),
    .B1(_06064_),
    .X(_06065_));
 sky130_fd_sc_hd__o21ba_1 _13853_ (.A1(_06038_),
    .A2(_06044_),
    .B1_N(_06065_),
    .X(_06066_));
 sky130_fd_sc_hd__o21a_1 _13854_ (.A1(_06041_),
    .A2(_06038_),
    .B1(_06043_),
    .X(_06067_));
 sky130_fd_sc_hd__mux2_1 _13855_ (.A0(_06020_),
    .A1(_06017_),
    .S(_06012_),
    .X(_06068_));
 sky130_fd_sc_hd__xnor2_1 _13856_ (.A(_06019_),
    .B(_06068_),
    .Y(_06069_));
 sky130_fd_sc_hd__a2111o_1 _13857_ (.A1(_06036_),
    .A2(_06038_),
    .B1(_06066_),
    .C1(_06067_),
    .D1(_06069_),
    .X(_06070_));
 sky130_fd_sc_hd__o2bb2a_1 _13858_ (.A1_N(_05992_),
    .A2_N(_05993_),
    .B1(_06022_),
    .B2(_06070_),
    .X(_06071_));
 sky130_fd_sc_hd__and2_1 _13859_ (.A(_06022_),
    .B(_06070_),
    .X(_06072_));
 sky130_fd_sc_hd__o22a_1 _13860_ (.A1(_05959_),
    .A2(_05990_),
    .B1(_06071_),
    .B2(_06072_),
    .X(_06073_));
 sky130_fd_sc_hd__a21o_1 _13861_ (.A1(_05959_),
    .A2(_05990_),
    .B1(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__xnor2_1 _13862_ (.A(_05950_),
    .B(_05952_),
    .Y(_06075_));
 sky130_fd_sc_hd__mux2_1 _13863_ (.A0(_05905_),
    .A1(_05906_),
    .S(_05879_),
    .X(_06076_));
 sky130_fd_sc_hd__xnor2_1 _13864_ (.A(_05878_),
    .B(_06076_),
    .Y(_06077_));
 sky130_fd_sc_hd__a211o_1 _13865_ (.A1(_05957_),
    .A2(_06075_),
    .B1(_06077_),
    .C1(_05922_),
    .X(_06078_));
 sky130_fd_sc_hd__or3_1 _13866_ (.A(_05922_),
    .B(_05949_),
    .C(_06075_),
    .X(_06079_));
 sky130_fd_sc_hd__a31o_1 _13867_ (.A1(_05922_),
    .A2(_05949_),
    .A3(_06075_),
    .B1(_06077_),
    .X(_06080_));
 sky130_fd_sc_hd__a22o_1 _13868_ (.A1(_06074_),
    .A2(_06078_),
    .B1(_06079_),
    .B2(_06080_),
    .X(_06081_));
 sky130_fd_sc_hd__a22o_1 _13869_ (.A1(_05860_),
    .A2(_05908_),
    .B1(_05955_),
    .B2(_06081_),
    .X(_06082_));
 sky130_fd_sc_hd__nor2_1 _13870_ (.A(_05801_),
    .B(_05855_),
    .Y(_06083_));
 sky130_fd_sc_hd__a22o_1 _13871_ (.A1(_05752_),
    .A2(_05753_),
    .B1(_05785_),
    .B2(_05751_),
    .X(_06084_));
 sky130_fd_sc_hd__o21a_2 _13872_ (.A1(_05751_),
    .A2(_05785_),
    .B1(_06084_),
    .X(_06085_));
 sky130_fd_sc_hd__nor2_1 _13873_ (.A(_05763_),
    .B(_05768_),
    .Y(_06086_));
 sky130_fd_sc_hd__a21oi_2 _13874_ (.A1(_05763_),
    .A2(_05768_),
    .B1(_05760_),
    .Y(_06087_));
 sky130_fd_sc_hd__and2_1 _13875_ (.A(_05765_),
    .B(_05766_),
    .X(_06088_));
 sky130_fd_sc_hd__o211a_1 _13876_ (.A1(_05765_),
    .A2(_05766_),
    .B1(net42),
    .C1(_05472_),
    .X(_06089_));
 sky130_fd_sc_hd__a41o_1 _13877_ (.A1(net47),
    .A2(net43),
    .A3(_05585_),
    .A4(_05587_),
    .B1(_05774_),
    .X(_06090_));
 sky130_fd_sc_hd__o21ai_2 _13878_ (.A1(_05565_),
    .A2(_05534_),
    .B1(_05775_),
    .Y(_06091_));
 sky130_fd_sc_hd__o211ai_4 _13879_ (.A1(_06088_),
    .A2(_06089_),
    .B1(_06090_),
    .C1(_06091_),
    .Y(_06092_));
 sky130_fd_sc_hd__a211o_2 _13880_ (.A1(_06090_),
    .A2(_06091_),
    .B1(_06088_),
    .C1(_06089_),
    .X(_06093_));
 sky130_fd_sc_hd__inv_1 _13881_ (.A(net41),
    .Y(_06094_));
 sky130_fd_sc_hd__nor2_1 _13882_ (.A(_06094_),
    .B(_05534_),
    .Y(_06095_));
 sky130_fd_sc_hd__nor3_1 _13883_ (.A(_05573_),
    .B(_05538_),
    .C(_05539_),
    .Y(_06096_));
 sky130_fd_sc_hd__or3_1 _13884_ (.A(_05565_),
    .B(_05543_),
    .C(_05545_),
    .X(_06097_));
 sky130_fd_sc_hd__xor2_1 _13885_ (.A(_06096_),
    .B(_06097_),
    .X(_06098_));
 sky130_fd_sc_hd__xnor2_2 _13886_ (.A(_06095_),
    .B(_06098_),
    .Y(_06099_));
 sky130_fd_sc_hd__a21oi_2 _13887_ (.A1(_06092_),
    .A2(_06093_),
    .B1(_06099_),
    .Y(_06100_));
 sky130_fd_sc_hd__and3_1 _13888_ (.A(_06099_),
    .B(_06092_),
    .C(_06093_),
    .X(_06101_));
 sky130_fd_sc_hd__o22ai_4 _13889_ (.A1(_06086_),
    .A2(_06087_),
    .B1(_06100_),
    .B2(_06101_),
    .Y(_06102_));
 sky130_fd_sc_hd__or4_4 _13890_ (.A(_06086_),
    .B(_06087_),
    .C(_06100_),
    .D(_06101_),
    .X(_06103_));
 sky130_fd_sc_hd__nand2_2 _13891_ (.A(net22),
    .B(_05683_),
    .Y(_06104_));
 sky130_fd_sc_hd__nand2_1 _13892_ (.A(net1030),
    .B(_05893_),
    .Y(_06105_));
 sky130_fd_sc_hd__inv_2 _13893_ (.A(net30),
    .Y(_06106_));
 sky130_fd_sc_hd__nor2_1 _13894_ (.A(_06106_),
    .B(_05567_),
    .Y(_06107_));
 sky130_fd_sc_hd__xor2_2 _13895_ (.A(_06105_),
    .B(_06107_),
    .X(_06108_));
 sky130_fd_sc_hd__xnor2_4 _13896_ (.A(_06104_),
    .B(_06108_),
    .Y(_06109_));
 sky130_fd_sc_hd__a21bo_1 _13897_ (.A1(_05756_),
    .A2(_05757_),
    .B1_N(_05758_),
    .X(_06110_));
 sky130_fd_sc_hd__o21a_1 _13898_ (.A1(_05756_),
    .A2(_05757_),
    .B1(_06110_),
    .X(_06111_));
 sky130_fd_sc_hd__nand2_1 _13899_ (.A(net40),
    .B(_05472_),
    .Y(_06112_));
 sky130_fd_sc_hd__and3_1 _13900_ (.A(net33),
    .B(_05478_),
    .C(_05479_),
    .X(_06113_));
 sky130_fd_sc_hd__and3_1 _13901_ (.A(net37),
    .B(_05475_),
    .C(_05476_),
    .X(_06114_));
 sky130_fd_sc_hd__xor2_1 _13902_ (.A(_06113_),
    .B(_06114_),
    .X(_06115_));
 sky130_fd_sc_hd__xnor2_2 _13903_ (.A(_06112_),
    .B(_06115_),
    .Y(_06116_));
 sky130_fd_sc_hd__xor2_2 _13904_ (.A(_06111_),
    .B(_06116_),
    .X(_06117_));
 sky130_fd_sc_hd__xnor2_4 _13905_ (.A(_06109_),
    .B(_06117_),
    .Y(_06118_));
 sky130_fd_sc_hd__a21oi_2 _13906_ (.A1(_06102_),
    .A2(_06103_),
    .B1(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__and3_1 _13907_ (.A(_06118_),
    .B(_06102_),
    .C(_06103_),
    .X(_06120_));
 sky130_fd_sc_hd__a21o_1 _13908_ (.A1(_05772_),
    .A2(_05783_),
    .B1(_05770_),
    .X(_06121_));
 sky130_fd_sc_hd__or2_1 _13909_ (.A(_05772_),
    .B(_05783_),
    .X(_06122_));
 sky130_fd_sc_hd__o211a_1 _13910_ (.A1(_06119_),
    .A2(_06120_),
    .B1(_06121_),
    .C1(_06122_),
    .X(_06123_));
 sky130_fd_sc_hd__a21oi_2 _13911_ (.A1(_05772_),
    .A2(_05783_),
    .B1(_05770_),
    .Y(_06124_));
 sky130_fd_sc_hd__nor2_1 _13912_ (.A(_05772_),
    .B(_05783_),
    .Y(_06125_));
 sky130_fd_sc_hd__a21o_1 _13913_ (.A1(_06102_),
    .A2(_06103_),
    .B1(_06118_),
    .X(_06126_));
 sky130_fd_sc_hd__nand3_1 _13914_ (.A(_06118_),
    .B(_06102_),
    .C(_06103_),
    .Y(_06127_));
 sky130_fd_sc_hd__o211a_1 _13915_ (.A1(_06124_),
    .A2(_06125_),
    .B1(_06126_),
    .C1(_06127_),
    .X(_06128_));
 sky130_fd_sc_hd__a2bb2oi_1 _13916_ (.A1_N(_05743_),
    .A2_N(_05744_),
    .B1(_05745_),
    .B2(_05746_),
    .Y(_06129_));
 sky130_fd_sc_hd__o21ai_4 _13917_ (.A1(_05742_),
    .A2(_06129_),
    .B1(_05748_),
    .Y(_06130_));
 sky130_fd_sc_hd__buf_4 _13918_ (.A(_05721_),
    .X(_06131_));
 sky130_fd_sc_hd__o211a_1 _13919_ (.A1(_05725_),
    .A2(_05728_),
    .B1(\top0.periodTop_r[0] ),
    .C1(_06131_),
    .X(_06132_));
 sky130_fd_sc_hd__a21o_2 _13920_ (.A1(_05725_),
    .A2(_05728_),
    .B1(_06132_),
    .X(_06133_));
 sky130_fd_sc_hd__a32o_1 _13921_ (.A1(\top0.matmul0.beta_pass[15] ),
    .A2(_05436_),
    .A3(_05719_),
    .B1(_05465_),
    .B2(\top0.c_out_calc[15] ),
    .X(_06134_));
 sky130_fd_sc_hd__a31o_4 _13922_ (.A1(\top0.matmul0.alpha_pass[15] ),
    .A2(_05436_),
    .A3(_05717_),
    .B1(_06134_),
    .X(_06135_));
 sky130_fd_sc_hd__and2_2 _13923_ (.A(net65),
    .B(_06135_),
    .X(_06136_));
 sky130_fd_sc_hd__xnor2_1 _13924_ (.A(_06133_),
    .B(_06136_),
    .Y(_06137_));
 sky130_fd_sc_hd__xnor2_2 _13925_ (.A(_06130_),
    .B(_06137_),
    .Y(_06138_));
 sky130_fd_sc_hd__and3_2 _13926_ (.A(net51),
    .B(_05602_),
    .C(_05603_),
    .X(_06139_));
 sky130_fd_sc_hd__nand2_1 _13927_ (.A(net1025),
    .B(_05624_),
    .Y(_06140_));
 sky130_fd_sc_hd__nand2_2 _13928_ (.A(net48),
    .B(_05639_),
    .Y(_06141_));
 sky130_fd_sc_hd__xnor2_2 _13929_ (.A(_06140_),
    .B(_06141_),
    .Y(_06142_));
 sky130_fd_sc_hd__xnor2_4 _13930_ (.A(_06139_),
    .B(_06142_),
    .Y(_06143_));
 sky130_fd_sc_hd__or2b_1 _13931_ (.A(_05737_),
    .B_N(_05738_),
    .X(_06144_));
 sky130_fd_sc_hd__a32o_1 _13932_ (.A1(net51),
    .A2(_05639_),
    .A3(_05737_),
    .B1(_05624_),
    .B2(net56),
    .X(_06145_));
 sky130_fd_sc_hd__nand2_1 _13933_ (.A(_06144_),
    .B(_06145_),
    .Y(_06146_));
 sky130_fd_sc_hd__nand2_1 _13934_ (.A(net64),
    .B(_05721_),
    .Y(_06147_));
 sky130_fd_sc_hd__and3_1 _13935_ (.A(net56),
    .B(_05723_),
    .C(_05724_),
    .X(_06148_));
 sky130_fd_sc_hd__and3_1 _13936_ (.A(net60),
    .B(_05726_),
    .C(_05727_),
    .X(_06149_));
 sky130_fd_sc_hd__xnor2_1 _13937_ (.A(_06148_),
    .B(_06149_),
    .Y(_06150_));
 sky130_fd_sc_hd__xnor2_1 _13938_ (.A(_06147_),
    .B(_06150_),
    .Y(_06151_));
 sky130_fd_sc_hd__nor2_1 _13939_ (.A(_06146_),
    .B(_06151_),
    .Y(_06152_));
 sky130_fd_sc_hd__nand2_1 _13940_ (.A(_06146_),
    .B(_06151_),
    .Y(_06153_));
 sky130_fd_sc_hd__and2b_1 _13941_ (.A_N(_06152_),
    .B(_06153_),
    .X(_06154_));
 sky130_fd_sc_hd__xnor2_4 _13942_ (.A(_06143_),
    .B(_06154_),
    .Y(_06155_));
 sky130_fd_sc_hd__a21bo_1 _13943_ (.A1(_05779_),
    .A2(_05781_),
    .B1_N(_05777_),
    .X(_06156_));
 sky130_fd_sc_hd__o21a_1 _13944_ (.A1(_05779_),
    .A2(_05781_),
    .B1(_06156_),
    .X(_06157_));
 sky130_fd_sc_hd__a21bo_1 _13945_ (.A1(_05734_),
    .A2(_05740_),
    .B1_N(_05730_),
    .X(_06158_));
 sky130_fd_sc_hd__o21a_1 _13946_ (.A1(_05734_),
    .A2(_05740_),
    .B1(_06158_),
    .X(_06159_));
 sky130_fd_sc_hd__xnor2_2 _13947_ (.A(_06157_),
    .B(_06159_),
    .Y(_06160_));
 sky130_fd_sc_hd__xor2_2 _13948_ (.A(_06155_),
    .B(_06160_),
    .X(_06161_));
 sky130_fd_sc_hd__o211a_1 _13949_ (.A1(_06123_),
    .A2(_06128_),
    .B1(_06138_),
    .C1(_06161_),
    .X(_06162_));
 sky130_fd_sc_hd__xnor2_1 _13950_ (.A(_06155_),
    .B(_06160_),
    .Y(_06163_));
 sky130_fd_sc_hd__a211o_1 _13951_ (.A1(_06126_),
    .A2(_06127_),
    .B1(_06124_),
    .C1(_06125_),
    .X(_06164_));
 sky130_fd_sc_hd__a211o_1 _13952_ (.A1(_06121_),
    .A2(_06122_),
    .B1(_06119_),
    .C1(_06120_),
    .X(_06165_));
 sky130_fd_sc_hd__and4_1 _13953_ (.A(_06163_),
    .B(_06164_),
    .C(_06165_),
    .D(_06138_),
    .X(_06166_));
 sky130_fd_sc_hd__or4_1 _13954_ (.A(_06163_),
    .B(_06123_),
    .C(_06128_),
    .D(_06138_),
    .X(_06167_));
 sky130_fd_sc_hd__a211o_1 _13955_ (.A1(_06164_),
    .A2(_06165_),
    .B1(_06138_),
    .C1(_06161_),
    .X(_06168_));
 sky130_fd_sc_hd__and4bb_1 _13956_ (.A_N(_06162_),
    .B_N(_06166_),
    .C(_06167_),
    .D(_06168_),
    .X(_06169_));
 sky130_fd_sc_hd__xor2_2 _13957_ (.A(_06085_),
    .B(_06169_),
    .X(_06170_));
 sky130_fd_sc_hd__nor2_2 _13958_ (.A(_05790_),
    .B(_05792_),
    .Y(_06171_));
 sky130_fd_sc_hd__o32a_1 _13959_ (.A1(_05786_),
    .A2(_05787_),
    .A3(_05796_),
    .B1(_05794_),
    .B2(_05789_),
    .X(_06172_));
 sky130_fd_sc_hd__or2_1 _13960_ (.A(_05795_),
    .B(_05789_),
    .X(_06173_));
 sky130_fd_sc_hd__o211a_1 _13961_ (.A1(_05786_),
    .A2(_05787_),
    .B1(_06173_),
    .C1(_06171_),
    .X(_06174_));
 sky130_fd_sc_hd__o21bai_1 _13962_ (.A1(_06171_),
    .A2(_06172_),
    .B1_N(_06174_),
    .Y(_06175_));
 sky130_fd_sc_hd__xor2_1 _13963_ (.A(_06170_),
    .B(_06175_),
    .X(_06176_));
 sky130_fd_sc_hd__a211o_1 _13964_ (.A1(_05799_),
    .A2(_06083_),
    .B1(_05857_),
    .C1(_06176_),
    .X(_06177_));
 sky130_fd_sc_hd__a21o_2 _13965_ (.A1(_05858_),
    .A2(_06082_),
    .B1(_06177_),
    .X(_06178_));
 sky130_fd_sc_hd__o22ai_4 _13966_ (.A1(_06171_),
    .A2(_06172_),
    .B1(_06174_),
    .B2(_06170_),
    .Y(_06179_));
 sky130_fd_sc_hd__inv_2 _13967_ (.A(_06103_),
    .Y(_06180_));
 sky130_fd_sc_hd__o21ai_4 _13968_ (.A1(_06118_),
    .A2(_06180_),
    .B1(_06102_),
    .Y(_06181_));
 sky130_fd_sc_hd__nand2_1 _13969_ (.A(net48),
    .B(_05605_),
    .Y(_06182_));
 sky130_fd_sc_hd__or3_1 _13970_ (.A(_05541_),
    .B(_05608_),
    .C(_05609_),
    .X(_06183_));
 sky130_fd_sc_hd__and3_1 _13971_ (.A(net45),
    .B(_05611_),
    .C(_05612_),
    .X(_06184_));
 sky130_fd_sc_hd__xnor2_1 _13972_ (.A(_06183_),
    .B(_06184_),
    .Y(_06185_));
 sky130_fd_sc_hd__xnor2_2 _13973_ (.A(_06182_),
    .B(_06185_),
    .Y(_06186_));
 sky130_fd_sc_hd__nand2_1 _13974_ (.A(net51),
    .B(_05605_),
    .Y(_06187_));
 sky130_fd_sc_hd__a32oi_2 _13975_ (.A1(net48),
    .A2(_05639_),
    .A3(_06139_),
    .B1(_05625_),
    .B2(net1025),
    .Y(_06188_));
 sky130_fd_sc_hd__a21oi_2 _13976_ (.A1(_06187_),
    .A2(_06141_),
    .B1(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__and3_1 _13977_ (.A(net1025),
    .B(_05723_),
    .C(_05724_),
    .X(_06190_));
 sky130_fd_sc_hd__clkbuf_2 _13978_ (.A(_06190_),
    .X(_06191_));
 sky130_fd_sc_hd__and3_1 _13979_ (.A(net56),
    .B(_05663_),
    .C(_05664_),
    .X(_06192_));
 sky130_fd_sc_hd__clkbuf_2 _13980_ (.A(_06192_),
    .X(_06193_));
 sky130_fd_sc_hd__or3_1 _13981_ (.A(_05657_),
    .B(_05718_),
    .C(_05720_),
    .X(_06194_));
 sky130_fd_sc_hd__xor2_1 _13982_ (.A(_06193_),
    .B(_06194_),
    .X(_06195_));
 sky130_fd_sc_hd__xnor2_1 _13983_ (.A(_06191_),
    .B(_06195_),
    .Y(_06196_));
 sky130_fd_sc_hd__xnor2_1 _13984_ (.A(_06189_),
    .B(_06196_),
    .Y(_06197_));
 sky130_fd_sc_hd__xnor2_2 _13985_ (.A(_06186_),
    .B(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__inv_2 _13986_ (.A(_06092_),
    .Y(_06199_));
 sky130_fd_sc_hd__o21ai_4 _13987_ (.A1(_06099_),
    .A2(_06199_),
    .B1(_06093_),
    .Y(_06200_));
 sky130_fd_sc_hd__o21ai_2 _13988_ (.A1(_06143_),
    .A2(_06152_),
    .B1(_06153_),
    .Y(_06201_));
 sky130_fd_sc_hd__xor2_1 _13989_ (.A(_06200_),
    .B(_06201_),
    .X(_06202_));
 sky130_fd_sc_hd__xnor2_2 _13990_ (.A(_06198_),
    .B(_06202_),
    .Y(_06203_));
 sky130_fd_sc_hd__xnor2_2 _13991_ (.A(_06181_),
    .B(_06203_),
    .Y(_06204_));
 sky130_fd_sc_hd__nand2_2 _13992_ (.A(net37),
    .B(net1015),
    .Y(_06205_));
 sky130_fd_sc_hd__and3_1 _13993_ (.A(net30),
    .B(_05478_),
    .C(_05479_),
    .X(_06206_));
 sky130_fd_sc_hd__and3_1 _13994_ (.A(net33),
    .B(_05475_),
    .C(_05476_),
    .X(_06207_));
 sky130_fd_sc_hd__xor2_2 _13995_ (.A(_06206_),
    .B(_06207_),
    .X(_06208_));
 sky130_fd_sc_hd__xnor2_4 _13996_ (.A(_06205_),
    .B(_06208_),
    .Y(_06209_));
 sky130_fd_sc_hd__and3_1 _13997_ (.A(\top0.matmul0.alpha_pass[1] ),
    .B(_05435_),
    .C(_05474_),
    .X(_06210_));
 sky130_fd_sc_hd__or4b_1 _13998_ (.A(_06210_),
    .B(_05493_),
    .C(_05494_),
    .D_N(_05490_),
    .X(_06211_));
 sky130_fd_sc_hd__nand2_4 _13999_ (.A(net27),
    .B(net22),
    .Y(_06212_));
 sky130_fd_sc_hd__o32a_1 _14000_ (.A1(_05683_),
    .A2(_06211_),
    .A3(_06212_),
    .B1(_05894_),
    .B2(net1030),
    .X(_06213_));
 sky130_fd_sc_hd__o21a_1 _14001_ (.A1(_05683_),
    .A2(_05894_),
    .B1(net24),
    .X(_06214_));
 sky130_fd_sc_hd__o22a_1 _14002_ (.A1(net32),
    .A2(_06213_),
    .B1(_06214_),
    .B2(net1030),
    .X(_06215_));
 sky130_fd_sc_hd__o21bai_1 _14003_ (.A1(_05567_),
    .A2(_05757_),
    .B1_N(net24),
    .Y(_06216_));
 sky130_fd_sc_hd__inv_2 _14004_ (.A(net1030),
    .Y(_06217_));
 sky130_fd_sc_hd__o22a_1 _14005_ (.A1(net1030),
    .A2(_06211_),
    .B1(_06212_),
    .B2(_05894_),
    .X(_06218_));
 sky130_fd_sc_hd__o32a_1 _14006_ (.A1(_06217_),
    .A2(_05501_),
    .A3(_05497_),
    .B1(_05686_),
    .B2(_06218_),
    .X(_06219_));
 sky130_fd_sc_hd__o2111a_2 _14007_ (.A1(_05894_),
    .A2(_05497_),
    .B1(_06215_),
    .C1(_06216_),
    .D1(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__xnor2_4 _14008_ (.A(_06209_),
    .B(_06220_),
    .Y(_06221_));
 sky130_fd_sc_hd__or3_2 _14009_ (.A(_05504_),
    .B(_05531_),
    .C(_05532_),
    .X(_06222_));
 sky130_fd_sc_hd__or3_1 _14010_ (.A(_05565_),
    .B(_05538_),
    .C(_05539_),
    .X(_06223_));
 sky130_fd_sc_hd__or3_1 _14011_ (.A(_06094_),
    .B(_05543_),
    .C(_05545_),
    .X(_06224_));
 sky130_fd_sc_hd__xor2_1 _14012_ (.A(_06223_),
    .B(_06224_),
    .X(_06225_));
 sky130_fd_sc_hd__xnor2_2 _14013_ (.A(_06222_),
    .B(_06225_),
    .Y(_06226_));
 sky130_fd_sc_hd__nor3_1 _14014_ (.A(_06094_),
    .B(_05822_),
    .C(_06097_),
    .Y(_06227_));
 sky130_fd_sc_hd__o21ai_1 _14015_ (.A1(_06094_),
    .A2(_05822_),
    .B1(_06097_),
    .Y(_06228_));
 sky130_fd_sc_hd__o21a_1 _14016_ (.A1(_06096_),
    .A2(_06227_),
    .B1(_06228_),
    .X(_06229_));
 sky130_fd_sc_hd__a22o_1 _14017_ (.A1(net39),
    .A2(_05517_),
    .B1(_06113_),
    .B2(_06114_),
    .X(_06230_));
 sky130_fd_sc_hd__o21a_1 _14018_ (.A1(_06113_),
    .A2(_06114_),
    .B1(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__xnor2_1 _14019_ (.A(_06229_),
    .B(_06231_),
    .Y(_06232_));
 sky130_fd_sc_hd__xnor2_2 _14020_ (.A(_06226_),
    .B(_06232_),
    .Y(_06233_));
 sky130_fd_sc_hd__nor2_1 _14021_ (.A(_06111_),
    .B(_06116_),
    .Y(_06234_));
 sky130_fd_sc_hd__nand2_1 _14022_ (.A(_06111_),
    .B(_06116_),
    .Y(_06235_));
 sky130_fd_sc_hd__o21ai_4 _14023_ (.A1(_06109_),
    .A2(_06234_),
    .B1(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__xnor2_2 _14024_ (.A(_06233_),
    .B(_06236_),
    .Y(_06237_));
 sky130_fd_sc_hd__xnor2_4 _14025_ (.A(_06221_),
    .B(_06237_),
    .Y(_06238_));
 sky130_fd_sc_hd__xnor2_4 _14026_ (.A(_06204_),
    .B(_06238_),
    .Y(_06239_));
 sky130_fd_sc_hd__or4_1 _14027_ (.A(_06124_),
    .B(_06125_),
    .C(_06119_),
    .D(_06120_),
    .X(_06240_));
 sky130_fd_sc_hd__o22a_1 _14028_ (.A1(_06124_),
    .A2(_06125_),
    .B1(_06119_),
    .B2(_06120_),
    .X(_06241_));
 sky130_fd_sc_hd__a21oi_1 _14029_ (.A1(_06161_),
    .A2(_06240_),
    .B1(_06241_),
    .Y(_06242_));
 sky130_fd_sc_hd__a22o_1 _14030_ (.A1(net64),
    .A2(_06131_),
    .B1(_06148_),
    .B2(_06149_),
    .X(_06243_));
 sky130_fd_sc_hd__o21a_1 _14031_ (.A1(_06148_),
    .A2(_06149_),
    .B1(_06243_),
    .X(_06244_));
 sky130_fd_sc_hd__nand2_1 _14032_ (.A(net64),
    .B(_06135_),
    .Y(_06245_));
 sky130_fd_sc_hd__xor2_1 _14033_ (.A(_06244_),
    .B(_06245_),
    .X(_06246_));
 sky130_fd_sc_hd__and2b_1 _14034_ (.A_N(_06159_),
    .B(_06157_),
    .X(_06247_));
 sky130_fd_sc_hd__or2b_1 _14035_ (.A(_06157_),
    .B_N(_06159_),
    .X(_06248_));
 sky130_fd_sc_hd__o21ai_2 _14036_ (.A1(_06155_),
    .A2(_06247_),
    .B1(_06248_),
    .Y(_06249_));
 sky130_fd_sc_hd__xnor2_1 _14037_ (.A(_06246_),
    .B(_06249_),
    .Y(_06250_));
 sky130_fd_sc_hd__nor2_1 _14038_ (.A(_06242_),
    .B(_06250_),
    .Y(_06251_));
 sky130_fd_sc_hd__nand2_1 _14039_ (.A(_06242_),
    .B(_06250_),
    .Y(_06252_));
 sky130_fd_sc_hd__and2b_1 _14040_ (.A_N(_06251_),
    .B(_06252_),
    .X(_06253_));
 sky130_fd_sc_hd__xor2_2 _14041_ (.A(_06239_),
    .B(_06253_),
    .X(_06254_));
 sky130_fd_sc_hd__or2_1 _14042_ (.A(_06179_),
    .B(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__nand2_2 _14043_ (.A(_06179_),
    .B(_06254_),
    .Y(_06256_));
 sky130_fd_sc_hd__nand2_1 _14044_ (.A(_06255_),
    .B(_06256_),
    .Y(_06257_));
 sky130_fd_sc_hd__nor2_1 _14045_ (.A(_06085_),
    .B(_06130_),
    .Y(_06258_));
 sky130_fd_sc_hd__a21oi_1 _14046_ (.A1(_06085_),
    .A2(_06130_),
    .B1(_06136_),
    .Y(_06259_));
 sky130_fd_sc_hd__or2_2 _14047_ (.A(_06258_),
    .B(_06259_),
    .X(_06260_));
 sky130_fd_sc_hd__and3_1 _14048_ (.A(_06161_),
    .B(_06164_),
    .C(_06165_),
    .X(_06261_));
 sky130_fd_sc_hd__a21oi_1 _14049_ (.A1(_06164_),
    .A2(_06165_),
    .B1(_06161_),
    .Y(_06262_));
 sky130_fd_sc_hd__nor2_2 _14050_ (.A(_06261_),
    .B(_06262_),
    .Y(_06263_));
 sky130_fd_sc_hd__nand2_1 _14051_ (.A(_06263_),
    .B(_06133_),
    .Y(_06264_));
 sky130_fd_sc_hd__o2111ai_4 _14052_ (.A1(_06263_),
    .A2(_06133_),
    .B1(_06136_),
    .C1(_06130_),
    .D1(_06085_),
    .Y(_06265_));
 sky130_fd_sc_hd__o21ai_4 _14053_ (.A1(_06260_),
    .A2(_06264_),
    .B1(_06265_),
    .Y(_06266_));
 sky130_fd_sc_hd__nor2_1 _14054_ (.A(_06263_),
    .B(_06133_),
    .Y(_06267_));
 sky130_fd_sc_hd__buf_4 _14055_ (.A(_06135_),
    .X(_06268_));
 sky130_fd_sc_hd__nand2_1 _14056_ (.A(net65),
    .B(_06268_),
    .Y(_06269_));
 sky130_fd_sc_hd__and3b_1 _14057_ (.A_N(_06133_),
    .B(_06269_),
    .C(_06258_),
    .X(_06270_));
 sky130_fd_sc_hd__and3b_1 _14058_ (.A_N(_06263_),
    .B(_06269_),
    .C(_06258_),
    .X(_06271_));
 sky130_fd_sc_hd__a211o_1 _14059_ (.A1(_06260_),
    .A2(_06267_),
    .B1(_06270_),
    .C1(_06271_),
    .X(_06272_));
 sky130_fd_sc_hd__or2_1 _14060_ (.A(_06266_),
    .B(_06272_),
    .X(_06273_));
 sky130_fd_sc_hd__xor2_1 _14061_ (.A(_06257_),
    .B(_06273_),
    .X(_06274_));
 sky130_fd_sc_hd__xnor2_2 _14062_ (.A(_06178_),
    .B(_06274_),
    .Y(_06275_));
 sky130_fd_sc_hd__or2_1 _14063_ (.A(\top0.svm0.state[1] ),
    .B(\top0.svm0.state[0] ),
    .X(_06276_));
 sky130_fd_sc_hd__clkbuf_4 _14064_ (.A(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__a21o_1 _14065_ (.A1(\top0.svm0.state[1] ),
    .A2(\top0.svm0.state[0] ),
    .B1(net171),
    .X(_06278_));
 sky130_fd_sc_hd__nand2_4 _14066_ (.A(_06277_),
    .B(_06278_),
    .Y(_06279_));
 sky130_fd_sc_hd__clkbuf_4 _14067_ (.A(_06279_),
    .X(_06280_));
 sky130_fd_sc_hd__a22o_1 _14068_ (.A1(_05465_),
    .A2(_06275_),
    .B1(_06280_),
    .B2(net736),
    .X(_00019_));
 sky130_fd_sc_hd__nand2_2 _14069_ (.A(net56),
    .B(_05721_),
    .Y(_06281_));
 sky130_fd_sc_hd__and3_1 _14070_ (.A(net51),
    .B(_05723_),
    .C(_05724_),
    .X(_06282_));
 sky130_fd_sc_hd__and3_1 _14071_ (.A(net1025),
    .B(_05726_),
    .C(_05727_),
    .X(_06283_));
 sky130_fd_sc_hd__xnor2_2 _14072_ (.A(_06282_),
    .B(_06283_),
    .Y(_06284_));
 sky130_fd_sc_hd__xnor2_4 _14073_ (.A(_06281_),
    .B(_06284_),
    .Y(_06285_));
 sky130_fd_sc_hd__a32o_1 _14074_ (.A1(net48),
    .A2(_05604_),
    .A3(_06184_),
    .B1(_05624_),
    .B2(net51),
    .X(_06286_));
 sky130_fd_sc_hd__a21o_1 _14075_ (.A1(net48),
    .A2(_05605_),
    .B1(_06184_),
    .X(_06287_));
 sky130_fd_sc_hd__nand2_2 _14076_ (.A(_06286_),
    .B(_06287_),
    .Y(_06288_));
 sky130_fd_sc_hd__and3_1 _14077_ (.A(net45),
    .B(_05602_),
    .C(_05603_),
    .X(_06289_));
 sky130_fd_sc_hd__or3_1 _14078_ (.A(_05530_),
    .B(_05608_),
    .C(_05609_),
    .X(_06290_));
 sky130_fd_sc_hd__or3_1 _14079_ (.A(_05565_),
    .B(_05637_),
    .C(_05638_),
    .X(_06291_));
 sky130_fd_sc_hd__xor2_1 _14080_ (.A(_06290_),
    .B(_06291_),
    .X(_06292_));
 sky130_fd_sc_hd__xnor2_2 _14081_ (.A(_06289_),
    .B(_06292_),
    .Y(_06293_));
 sky130_fd_sc_hd__xnor2_2 _14082_ (.A(_06288_),
    .B(_06293_),
    .Y(_06294_));
 sky130_fd_sc_hd__xnor2_4 _14083_ (.A(_06285_),
    .B(_06294_),
    .Y(_06295_));
 sky130_fd_sc_hd__nor2_1 _14084_ (.A(_06229_),
    .B(_06231_),
    .Y(_06296_));
 sky130_fd_sc_hd__a21oi_1 _14085_ (.A1(_06229_),
    .A2(_06231_),
    .B1(_06226_),
    .Y(_06297_));
 sky130_fd_sc_hd__a21oi_1 _14086_ (.A1(_06189_),
    .A2(_06196_),
    .B1(_06186_),
    .Y(_06298_));
 sky130_fd_sc_hd__nor2_1 _14087_ (.A(_06189_),
    .B(_06196_),
    .Y(_06299_));
 sky130_fd_sc_hd__nor4_1 _14088_ (.A(_06296_),
    .B(_06297_),
    .C(_06298_),
    .D(_06299_),
    .Y(_06300_));
 sky130_fd_sc_hd__o22a_1 _14089_ (.A1(_06296_),
    .A2(_06297_),
    .B1(_06298_),
    .B2(_06299_),
    .X(_06301_));
 sky130_fd_sc_hd__nor2_2 _14090_ (.A(_06300_),
    .B(_06301_),
    .Y(_06302_));
 sky130_fd_sc_hd__xnor2_4 _14091_ (.A(_06295_),
    .B(_06302_),
    .Y(_06303_));
 sky130_fd_sc_hd__nand2_1 _14092_ (.A(_06233_),
    .B(_06236_),
    .Y(_06304_));
 sky130_fd_sc_hd__o21bai_1 _14093_ (.A1(_06233_),
    .A2(_06236_),
    .B1_N(_06221_),
    .Y(_06305_));
 sky130_fd_sc_hd__nor3_1 _14094_ (.A(_05688_),
    .B(_05531_),
    .C(_05532_),
    .Y(_06306_));
 sky130_fd_sc_hd__or3_1 _14095_ (.A(_06094_),
    .B(_05538_),
    .C(_05539_),
    .X(_06307_));
 sky130_fd_sc_hd__or3_1 _14096_ (.A(_05504_),
    .B(_05543_),
    .C(_05545_),
    .X(_06308_));
 sky130_fd_sc_hd__xnor2_1 _14097_ (.A(_06307_),
    .B(_06308_),
    .Y(_06309_));
 sky130_fd_sc_hd__xor2_1 _14098_ (.A(_06306_),
    .B(_06309_),
    .X(_06310_));
 sky130_fd_sc_hd__or2_1 _14099_ (.A(_06222_),
    .B(_06224_),
    .X(_06311_));
 sky130_fd_sc_hd__a21o_1 _14100_ (.A1(_06222_),
    .A2(_06224_),
    .B1(_06223_),
    .X(_06312_));
 sky130_fd_sc_hd__and2_1 _14101_ (.A(_06206_),
    .B(_06207_),
    .X(_06313_));
 sky130_fd_sc_hd__o211a_1 _14102_ (.A1(_06206_),
    .A2(_06207_),
    .B1(net37),
    .C1(_05472_),
    .X(_06314_));
 sky130_fd_sc_hd__a211o_1 _14103_ (.A1(_06311_),
    .A2(_06312_),
    .B1(_06313_),
    .C1(_06314_),
    .X(_06315_));
 sky130_fd_sc_hd__o211ai_1 _14104_ (.A1(_06313_),
    .A2(_06314_),
    .B1(_06311_),
    .C1(_06312_),
    .Y(_06316_));
 sky130_fd_sc_hd__and3_1 _14105_ (.A(_06310_),
    .B(_06315_),
    .C(_06316_),
    .X(_06317_));
 sky130_fd_sc_hd__a21oi_1 _14106_ (.A1(_06315_),
    .A2(_06316_),
    .B1(_06310_),
    .Y(_06318_));
 sky130_fd_sc_hd__or2_1 _14107_ (.A(_06317_),
    .B(_06318_),
    .X(_06319_));
 sky130_fd_sc_hd__and2_2 _14108_ (.A(net25),
    .B(net20),
    .X(_06320_));
 sky130_fd_sc_hd__and4b_1 _14109_ (.A_N(net24),
    .B(_05489_),
    .C(_05491_),
    .D(net1030),
    .X(_06321_));
 sky130_fd_sc_hd__a41o_1 _14110_ (.A1(_05484_),
    .A2(_05486_),
    .A3(_06046_),
    .A4(_06320_),
    .B1(_06321_),
    .X(_06322_));
 sky130_fd_sc_hd__and2_2 _14111_ (.A(_06217_),
    .B(net22),
    .X(_06323_));
 sky130_fd_sc_hd__and3_1 _14112_ (.A(net32),
    .B(_05496_),
    .C(_06323_),
    .X(_06324_));
 sky130_fd_sc_hd__and4_1 _14113_ (.A(_05683_),
    .B(_05894_),
    .C(_05567_),
    .D(_06320_),
    .X(_06325_));
 sky130_fd_sc_hd__a221o_1 _14114_ (.A1(_06107_),
    .A2(_06322_),
    .B1(_06324_),
    .B2(_06047_),
    .C1(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__a21o_1 _14115_ (.A1(net24),
    .A2(_05894_),
    .B1(_05497_),
    .X(_06327_));
 sky130_fd_sc_hd__o211ai_4 _14116_ (.A1(_06209_),
    .A2(_06326_),
    .B1(_06327_),
    .C1(_06215_),
    .Y(_06328_));
 sky130_fd_sc_hd__nor3_2 _14117_ (.A(_05500_),
    .B(_05468_),
    .C(_05471_),
    .Y(_06329_));
 sky130_fd_sc_hd__and3_2 _14118_ (.A(net30),
    .B(_05520_),
    .C(_05521_),
    .X(_06330_));
 sky130_fd_sc_hd__xor2_2 _14119_ (.A(_06329_),
    .B(_06330_),
    .X(_06331_));
 sky130_fd_sc_hd__nand2_1 _14120_ (.A(net22),
    .B(_05497_),
    .Y(_06332_));
 sky130_fd_sc_hd__a22o_1 _14121_ (.A1(_05523_),
    .A2(_05524_),
    .B1(_05489_),
    .B2(_05491_),
    .X(_06333_));
 sky130_fd_sc_hd__and2_1 _14122_ (.A(net27),
    .B(_06333_),
    .X(_06334_));
 sky130_fd_sc_hd__nand2_1 _14123_ (.A(net1030),
    .B(_06023_),
    .Y(_06335_));
 sky130_fd_sc_hd__and3_1 _14124_ (.A(net22),
    .B(_06046_),
    .C(_05496_),
    .X(_06336_));
 sky130_fd_sc_hd__o22a_1 _14125_ (.A1(_06332_),
    .A2(_06334_),
    .B1(_06335_),
    .B2(_06336_),
    .X(_06337_));
 sky130_fd_sc_hd__xor2_2 _14126_ (.A(_06331_),
    .B(_06337_),
    .X(_06338_));
 sky130_fd_sc_hd__xnor2_1 _14127_ (.A(_06328_),
    .B(_06338_),
    .Y(_06339_));
 sky130_fd_sc_hd__xnor2_1 _14128_ (.A(_06319_),
    .B(_06339_),
    .Y(_06340_));
 sky130_fd_sc_hd__a21oi_1 _14129_ (.A1(_06304_),
    .A2(_06305_),
    .B1(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__and3_1 _14130_ (.A(_06304_),
    .B(_06305_),
    .C(_06340_),
    .X(_06342_));
 sky130_fd_sc_hd__nor2_2 _14131_ (.A(_06341_),
    .B(_06342_),
    .Y(_06343_));
 sky130_fd_sc_hd__xnor2_4 _14132_ (.A(_06303_),
    .B(_06343_),
    .Y(_06344_));
 sky130_fd_sc_hd__o21a_1 _14133_ (.A1(_06181_),
    .A2(_06203_),
    .B1(_06238_),
    .X(_06345_));
 sky130_fd_sc_hd__a21o_1 _14134_ (.A1(_06181_),
    .A2(_06203_),
    .B1(_06345_),
    .X(_06346_));
 sky130_fd_sc_hd__o21ba_1 _14135_ (.A1(_06200_),
    .A2(_06201_),
    .B1_N(_06198_),
    .X(_06347_));
 sky130_fd_sc_hd__a21oi_2 _14136_ (.A1(_06200_),
    .A2(_06201_),
    .B1(_06347_),
    .Y(_06348_));
 sky130_fd_sc_hd__nand2_1 _14137_ (.A(net60),
    .B(_06135_),
    .Y(_06349_));
 sky130_fd_sc_hd__o21a_1 _14138_ (.A1(_06191_),
    .A2(_06193_),
    .B1(_06131_),
    .X(_06350_));
 sky130_fd_sc_hd__buf_4 _14139_ (.A(_06131_),
    .X(_06351_));
 sky130_fd_sc_hd__a21oi_1 _14140_ (.A1(_06351_),
    .A2(_06193_),
    .B1(_06191_),
    .Y(_06352_));
 sky130_fd_sc_hd__o21ai_1 _14141_ (.A1(_06351_),
    .A2(_06193_),
    .B1(_06135_),
    .Y(_06353_));
 sky130_fd_sc_hd__o221a_1 _14142_ (.A1(_06135_),
    .A2(_06350_),
    .B1(_06352_),
    .B2(_06353_),
    .C1(net60),
    .X(_06354_));
 sky130_fd_sc_hd__a31o_1 _14143_ (.A1(_06191_),
    .A2(_06193_),
    .A3(_06349_),
    .B1(_06354_),
    .X(_06355_));
 sky130_fd_sc_hd__xor2_2 _14144_ (.A(_06348_),
    .B(_06355_),
    .X(_06356_));
 sky130_fd_sc_hd__xnor2_2 _14145_ (.A(_06346_),
    .B(_06356_),
    .Y(_06357_));
 sky130_fd_sc_hd__xnor2_4 _14146_ (.A(_06344_),
    .B(_06357_),
    .Y(_06358_));
 sky130_fd_sc_hd__or2b_1 _14147_ (.A(_06244_),
    .B_N(_06245_),
    .X(_06359_));
 sky130_fd_sc_hd__nor2_1 _14148_ (.A(_06124_),
    .B(_06125_),
    .Y(_06360_));
 sky130_fd_sc_hd__nand2_1 _14149_ (.A(_06155_),
    .B(_06247_),
    .Y(_06361_));
 sky130_fd_sc_hd__o21a_1 _14150_ (.A1(_06360_),
    .A2(_06249_),
    .B1(_06361_),
    .X(_06362_));
 sky130_fd_sc_hd__nor2_1 _14151_ (.A(_06119_),
    .B(_06120_),
    .Y(_06363_));
 sky130_fd_sc_hd__o22a_1 _14152_ (.A1(_06360_),
    .A2(_06361_),
    .B1(_06362_),
    .B2(_06363_),
    .X(_06364_));
 sky130_fd_sc_hd__and3_1 _14153_ (.A(net64),
    .B(_06268_),
    .C(_06244_),
    .X(_06365_));
 sky130_fd_sc_hd__a21o_1 _14154_ (.A1(_06249_),
    .A2(_06359_),
    .B1(_06365_),
    .X(_06366_));
 sky130_fd_sc_hd__a21oi_1 _14155_ (.A1(_06239_),
    .A2(_06252_),
    .B1(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__o211a_1 _14156_ (.A1(_06239_),
    .A2(_06251_),
    .B1(_06252_),
    .C1(_06366_),
    .X(_06368_));
 sky130_fd_sc_hd__o22a_2 _14157_ (.A1(_06359_),
    .A2(_06364_),
    .B1(_06367_),
    .B2(_06368_),
    .X(_06369_));
 sky130_fd_sc_hd__xor2_4 _14158_ (.A(_06358_),
    .B(_06369_),
    .X(_06370_));
 sky130_fd_sc_hd__nand2_1 _14159_ (.A(_06255_),
    .B(_06272_),
    .Y(_06371_));
 sky130_fd_sc_hd__o21ai_1 _14160_ (.A1(_06256_),
    .A2(_06266_),
    .B1(_06371_),
    .Y(_06372_));
 sky130_fd_sc_hd__inv_2 _14161_ (.A(_06266_),
    .Y(_06373_));
 sky130_fd_sc_hd__nor2_1 _14162_ (.A(_06179_),
    .B(_06254_),
    .Y(_06374_));
 sky130_fd_sc_hd__a21oi_1 _14163_ (.A1(_06256_),
    .A2(_06266_),
    .B1(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__o22a_1 _14164_ (.A1(_06255_),
    .A2(_06373_),
    .B1(_06375_),
    .B2(_06178_),
    .X(_06376_));
 sky130_fd_sc_hd__a211oi_1 _14165_ (.A1(_06260_),
    .A2(_06267_),
    .B1(_06270_),
    .C1(_06271_),
    .Y(_06377_));
 sky130_fd_sc_hd__mux2_1 _14166_ (.A0(_06256_),
    .A1(_06376_),
    .S(_06377_),
    .X(_06378_));
 sky130_fd_sc_hd__a21bo_1 _14167_ (.A1(_06178_),
    .A2(_06372_),
    .B1_N(_06378_),
    .X(_06379_));
 sky130_fd_sc_hd__xnor2_2 _14168_ (.A(_06370_),
    .B(_06379_),
    .Y(_06380_));
 sky130_fd_sc_hd__clkbuf_4 _14169_ (.A(_05465_),
    .X(_06381_));
 sky130_fd_sc_hd__a22o_1 _14170_ (.A1(net852),
    .A2(_06280_),
    .B1(_06380_),
    .B2(_06381_),
    .X(_00020_));
 sky130_fd_sc_hd__mux2_1 _14171_ (.A0(_06255_),
    .A1(_06256_),
    .S(_06370_),
    .X(_06382_));
 sky130_fd_sc_hd__mux2_1 _14172_ (.A0(_06373_),
    .A1(_06377_),
    .S(_06370_),
    .X(_06383_));
 sky130_fd_sc_hd__o22a_1 _14173_ (.A1(_06273_),
    .A2(_06382_),
    .B1(_06383_),
    .B2(_06257_),
    .X(_06384_));
 sky130_fd_sc_hd__o21a_1 _14174_ (.A1(_06374_),
    .A2(_06370_),
    .B1(_06266_),
    .X(_06385_));
 sky130_fd_sc_hd__a31o_1 _14175_ (.A1(_06256_),
    .A2(_06370_),
    .A3(_06371_),
    .B1(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__o21ba_1 _14176_ (.A1(_06178_),
    .A2(_06384_),
    .B1_N(_06386_),
    .X(_06387_));
 sky130_fd_sc_hd__o21ai_1 _14177_ (.A1(_06239_),
    .A2(_06251_),
    .B1(_06252_),
    .Y(_06388_));
 sky130_fd_sc_hd__o21ai_1 _14178_ (.A1(_06358_),
    .A2(_06366_),
    .B1(_06388_),
    .Y(_06389_));
 sky130_fd_sc_hd__nand2_1 _14179_ (.A(_06358_),
    .B(_06366_),
    .Y(_06390_));
 sky130_fd_sc_hd__inv_2 _14180_ (.A(_06356_),
    .Y(_06391_));
 sky130_fd_sc_hd__o21a_1 _14181_ (.A1(_06344_),
    .A2(_06391_),
    .B1(_06346_),
    .X(_06392_));
 sky130_fd_sc_hd__a21o_1 _14182_ (.A1(_06344_),
    .A2(_06391_),
    .B1(_06392_),
    .X(_06393_));
 sky130_fd_sc_hd__nand2_1 _14183_ (.A(net45),
    .B(_05625_),
    .Y(_06394_));
 sky130_fd_sc_hd__and3_1 _14184_ (.A(net44),
    .B(_05602_),
    .C(_05603_),
    .X(_06395_));
 sky130_fd_sc_hd__and3_1 _14185_ (.A(net41),
    .B(_05611_),
    .C(_05612_),
    .X(_06396_));
 sky130_fd_sc_hd__xor2_1 _14186_ (.A(_06395_),
    .B(_06396_),
    .X(_06397_));
 sky130_fd_sc_hd__xnor2_2 _14187_ (.A(_06394_),
    .B(_06397_),
    .Y(_06398_));
 sky130_fd_sc_hd__nor2_1 _14188_ (.A(_05565_),
    .B(_05731_),
    .Y(_06399_));
 sky130_fd_sc_hd__a32o_1 _14189_ (.A1(net44),
    .A2(_05639_),
    .A3(_06289_),
    .B1(_05625_),
    .B2(net48),
    .X(_06400_));
 sky130_fd_sc_hd__o21a_1 _14190_ (.A1(_06289_),
    .A2(_06399_),
    .B1(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__nand2_1 _14191_ (.A(net1025),
    .B(_05721_),
    .Y(_06402_));
 sky130_fd_sc_hd__and3_1 _14192_ (.A(net48),
    .B(_05723_),
    .C(_05724_),
    .X(_06403_));
 sky130_fd_sc_hd__and3_1 _14193_ (.A(net51),
    .B(_05726_),
    .C(_05727_),
    .X(_06404_));
 sky130_fd_sc_hd__xor2_1 _14194_ (.A(_06403_),
    .B(_06404_),
    .X(_06405_));
 sky130_fd_sc_hd__xnor2_1 _14195_ (.A(_06402_),
    .B(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__xor2_1 _14196_ (.A(_06401_),
    .B(_06406_),
    .X(_06407_));
 sky130_fd_sc_hd__xnor2_2 _14197_ (.A(_06398_),
    .B(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__nand2_1 _14198_ (.A(_06311_),
    .B(_06312_),
    .Y(_06409_));
 sky130_fd_sc_hd__or2_1 _14199_ (.A(_06313_),
    .B(_06314_),
    .X(_06410_));
 sky130_fd_sc_hd__nor2_1 _14200_ (.A(_06409_),
    .B(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__a21boi_1 _14201_ (.A1(_06409_),
    .A2(_06410_),
    .B1_N(_06310_),
    .Y(_06412_));
 sky130_fd_sc_hd__and2_1 _14202_ (.A(_06288_),
    .B(_06293_),
    .X(_06413_));
 sky130_fd_sc_hd__o21a_1 _14203_ (.A1(_06288_),
    .A2(_06293_),
    .B1(_06285_),
    .X(_06414_));
 sky130_fd_sc_hd__or4_4 _14204_ (.A(_06411_),
    .B(_06412_),
    .C(_06413_),
    .D(_06414_),
    .X(_06415_));
 sky130_fd_sc_hd__o22ai_2 _14205_ (.A1(_06411_),
    .A2(_06412_),
    .B1(_06413_),
    .B2(_06414_),
    .Y(_06416_));
 sky130_fd_sc_hd__nand3_2 _14206_ (.A(_06408_),
    .B(_06415_),
    .C(_06416_),
    .Y(_06417_));
 sky130_fd_sc_hd__a21o_1 _14207_ (.A1(_06415_),
    .A2(_06416_),
    .B1(_06408_),
    .X(_06418_));
 sky130_fd_sc_hd__and2_1 _14208_ (.A(_06328_),
    .B(_06338_),
    .X(_06419_));
 sky130_fd_sc_hd__o22a_1 _14209_ (.A1(_06317_),
    .A2(_06318_),
    .B1(_06338_),
    .B2(_06328_),
    .X(_06420_));
 sky130_fd_sc_hd__or3_2 _14210_ (.A(_05500_),
    .B(_05531_),
    .C(_05532_),
    .X(_06421_));
 sky130_fd_sc_hd__nor3_1 _14211_ (.A(_05504_),
    .B(_05538_),
    .C(_05539_),
    .Y(_06422_));
 sky130_fd_sc_hd__or3_2 _14212_ (.A(_05688_),
    .B(_05543_),
    .C(_05545_),
    .X(_06423_));
 sky130_fd_sc_hd__xor2_1 _14213_ (.A(_06422_),
    .B(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__xor2_2 _14214_ (.A(_06421_),
    .B(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__and3_2 _14215_ (.A(net27),
    .B(_05523_),
    .C(_05524_),
    .X(_06426_));
 sky130_fd_sc_hd__a21oi_2 _14216_ (.A1(_06330_),
    .A2(_06426_),
    .B1(_06329_),
    .Y(_06427_));
 sky130_fd_sc_hd__nor2_2 _14217_ (.A(_06330_),
    .B(_06426_),
    .Y(_06428_));
 sky130_fd_sc_hd__o31a_1 _14218_ (.A1(_05688_),
    .A2(_05822_),
    .A3(_06308_),
    .B1(_06307_),
    .X(_06429_));
 sky130_fd_sc_hd__and2b_1 _14219_ (.A_N(_06306_),
    .B(_06308_),
    .X(_06430_));
 sky130_fd_sc_hd__or4_1 _14220_ (.A(_06427_),
    .B(_06428_),
    .C(_06429_),
    .D(_06430_),
    .X(_06431_));
 sky130_fd_sc_hd__o22ai_2 _14221_ (.A1(_06427_),
    .A2(_06428_),
    .B1(_06429_),
    .B2(_06430_),
    .Y(_06432_));
 sky130_fd_sc_hd__and3_2 _14222_ (.A(_06425_),
    .B(_06431_),
    .C(_06432_),
    .X(_06433_));
 sky130_fd_sc_hd__a21oi_2 _14223_ (.A1(_06431_),
    .A2(_06432_),
    .B1(_06425_),
    .Y(_06434_));
 sky130_fd_sc_hd__nand2_2 _14224_ (.A(net30),
    .B(net1015),
    .Y(_06435_));
 sky130_fd_sc_hd__and3_1 _14225_ (.A(net28),
    .B(_05520_),
    .C(_05521_),
    .X(_06436_));
 sky130_fd_sc_hd__buf_2 _14226_ (.A(_06436_),
    .X(_06437_));
 sky130_fd_sc_hd__and3_2 _14227_ (.A(net22),
    .B(_05523_),
    .C(_05524_),
    .X(_06438_));
 sky130_fd_sc_hd__xnor2_2 _14228_ (.A(_06437_),
    .B(_06438_),
    .Y(_06439_));
 sky130_fd_sc_hd__xnor2_4 _14229_ (.A(_06435_),
    .B(_06439_),
    .Y(_06440_));
 sky130_fd_sc_hd__nand2_1 _14230_ (.A(_06046_),
    .B(_06426_),
    .Y(_06441_));
 sky130_fd_sc_hd__mux2_1 _14231_ (.A0(_06333_),
    .A1(_06441_),
    .S(_06331_),
    .X(_06442_));
 sky130_fd_sc_hd__o21ba_1 _14232_ (.A1(net28),
    .A2(_06331_),
    .B1_N(_06332_),
    .X(_06443_));
 sky130_fd_sc_hd__nand3_2 _14233_ (.A(_06440_),
    .B(_06442_),
    .C(_06443_),
    .Y(_06444_));
 sky130_fd_sc_hd__a21o_1 _14234_ (.A1(_06442_),
    .A2(_06443_),
    .B1(_06440_),
    .X(_06445_));
 sky130_fd_sc_hd__o211ai_2 _14235_ (.A1(_06433_),
    .A2(_06434_),
    .B1(_06444_),
    .C1(_06445_),
    .Y(_06446_));
 sky130_fd_sc_hd__a211o_1 _14236_ (.A1(_06444_),
    .A2(_06445_),
    .B1(_06433_),
    .C1(_06434_),
    .X(_06447_));
 sky130_fd_sc_hd__o211a_1 _14237_ (.A1(_06419_),
    .A2(_06420_),
    .B1(_06446_),
    .C1(_06447_),
    .X(_06448_));
 sky130_fd_sc_hd__a211oi_2 _14238_ (.A1(_06446_),
    .A2(_06447_),
    .B1(_06419_),
    .C1(_06420_),
    .Y(_06449_));
 sky130_fd_sc_hd__a211o_1 _14239_ (.A1(_06417_),
    .A2(_06418_),
    .B1(_06448_),
    .C1(_06449_),
    .X(_06450_));
 sky130_fd_sc_hd__o211ai_2 _14240_ (.A1(_06448_),
    .A2(_06449_),
    .B1(_06417_),
    .C1(_06418_),
    .Y(_06451_));
 sky130_fd_sc_hd__or4_1 _14241_ (.A(_06296_),
    .B(_06297_),
    .C(_06298_),
    .D(_06299_),
    .X(_06452_));
 sky130_fd_sc_hd__a21o_1 _14242_ (.A1(_06295_),
    .A2(_06452_),
    .B1(_06301_),
    .X(_06453_));
 sky130_fd_sc_hd__a22o_1 _14243_ (.A1(net56),
    .A2(_06131_),
    .B1(_06282_),
    .B2(_06283_),
    .X(_06454_));
 sky130_fd_sc_hd__o21a_1 _14244_ (.A1(_06282_),
    .A2(_06283_),
    .B1(_06454_),
    .X(_06455_));
 sky130_fd_sc_hd__nand2_1 _14245_ (.A(net56),
    .B(_06135_),
    .Y(_06456_));
 sky130_fd_sc_hd__xor2_1 _14246_ (.A(_06455_),
    .B(_06456_),
    .X(_06457_));
 sky130_fd_sc_hd__xor2_1 _14247_ (.A(_06453_),
    .B(_06457_),
    .X(_06458_));
 sky130_fd_sc_hd__a21o_1 _14248_ (.A1(_06450_),
    .A2(_06451_),
    .B1(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__nand3_1 _14249_ (.A(_06450_),
    .B(_06451_),
    .C(_06458_),
    .Y(_06460_));
 sky130_fd_sc_hd__o21bai_2 _14250_ (.A1(_06303_),
    .A2(_06341_),
    .B1_N(_06342_),
    .Y(_06461_));
 sky130_fd_sc_hd__a21oi_1 _14251_ (.A1(_06459_),
    .A2(_06460_),
    .B1(_06461_),
    .Y(_06462_));
 sky130_fd_sc_hd__and3_1 _14252_ (.A(_06461_),
    .B(_06459_),
    .C(_06460_),
    .X(_06463_));
 sky130_fd_sc_hd__or2_2 _14253_ (.A(_06462_),
    .B(_06463_),
    .X(_06464_));
 sky130_fd_sc_hd__a22oi_2 _14254_ (.A1(_06191_),
    .A2(_06193_),
    .B1(_06350_),
    .B2(net60),
    .Y(_06465_));
 sky130_fd_sc_hd__a21bo_1 _14255_ (.A1(_06349_),
    .A2(_06465_),
    .B1_N(_06348_),
    .X(_06466_));
 sky130_fd_sc_hd__o21a_1 _14256_ (.A1(_06349_),
    .A2(_06465_),
    .B1(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__xnor2_1 _14257_ (.A(_06464_),
    .B(_06467_),
    .Y(_06468_));
 sky130_fd_sc_hd__xnor2_2 _14258_ (.A(_06393_),
    .B(_06468_),
    .Y(_06469_));
 sky130_fd_sc_hd__a21oi_2 _14259_ (.A1(_06389_),
    .A2(_06390_),
    .B1(_06469_),
    .Y(_06470_));
 sky130_fd_sc_hd__and3_1 _14260_ (.A(_06389_),
    .B(_06390_),
    .C(_06469_),
    .X(_06471_));
 sky130_fd_sc_hd__nor2_2 _14261_ (.A(_06470_),
    .B(_06471_),
    .Y(_06472_));
 sky130_fd_sc_hd__xnor2_2 _14262_ (.A(_06387_),
    .B(_06472_),
    .Y(_06473_));
 sky130_fd_sc_hd__a22o_1 _14263_ (.A1(net853),
    .A2(_06280_),
    .B1(_06473_),
    .B2(_06381_),
    .X(_00021_));
 sky130_fd_sc_hd__o21ba_2 _14264_ (.A1(_06387_),
    .A2(_06471_),
    .B1_N(_06470_),
    .X(_06474_));
 sky130_fd_sc_hd__a21o_1 _14265_ (.A1(_06464_),
    .A2(_06467_),
    .B1(_06393_),
    .X(_06475_));
 sky130_fd_sc_hd__o21a_1 _14266_ (.A1(_06464_),
    .A2(_06467_),
    .B1(_06475_),
    .X(_06476_));
 sky130_fd_sc_hd__o211a_1 _14267_ (.A1(_06433_),
    .A2(_06434_),
    .B1(_06444_),
    .C1(_06445_),
    .X(_06477_));
 sky130_fd_sc_hd__a211oi_1 _14268_ (.A1(_06444_),
    .A2(_06445_),
    .B1(_06433_),
    .C1(_06434_),
    .Y(_06478_));
 sky130_fd_sc_hd__or4_2 _14269_ (.A(_06419_),
    .B(_06420_),
    .C(_06477_),
    .D(_06478_),
    .X(_06479_));
 sky130_fd_sc_hd__o22a_1 _14270_ (.A1(_06419_),
    .A2(_06420_),
    .B1(_06477_),
    .B2(_06478_),
    .X(_06480_));
 sky130_fd_sc_hd__a31oi_4 _14271_ (.A1(_06417_),
    .A2(_06418_),
    .A3(_06479_),
    .B1(_06480_),
    .Y(_06481_));
 sky130_fd_sc_hd__a21boi_4 _14272_ (.A1(_06408_),
    .A2(_06415_),
    .B1_N(_06416_),
    .Y(_06482_));
 sky130_fd_sc_hd__a22o_1 _14273_ (.A1(net1025),
    .A2(_06351_),
    .B1(_06403_),
    .B2(_06404_),
    .X(_06483_));
 sky130_fd_sc_hd__o21a_2 _14274_ (.A1(_06403_),
    .A2(_06404_),
    .B1(_06483_),
    .X(_06484_));
 sky130_fd_sc_hd__and2_2 _14275_ (.A(net55),
    .B(_06135_),
    .X(_06485_));
 sky130_fd_sc_hd__xnor2_2 _14276_ (.A(_06484_),
    .B(_06485_),
    .Y(_06486_));
 sky130_fd_sc_hd__xnor2_4 _14277_ (.A(_06482_),
    .B(_06486_),
    .Y(_06487_));
 sky130_fd_sc_hd__nand2_2 _14278_ (.A(net51),
    .B(_05721_),
    .Y(_06488_));
 sky130_fd_sc_hd__and3_1 _14279_ (.A(net45),
    .B(_05723_),
    .C(_05724_),
    .X(_06489_));
 sky130_fd_sc_hd__and3_1 _14280_ (.A(net48),
    .B(_05726_),
    .C(_05727_),
    .X(_06490_));
 sky130_fd_sc_hd__xnor2_2 _14281_ (.A(_06489_),
    .B(_06490_),
    .Y(_06491_));
 sky130_fd_sc_hd__xnor2_4 _14282_ (.A(_06488_),
    .B(_06491_),
    .Y(_06492_));
 sky130_fd_sc_hd__a22o_1 _14283_ (.A1(net45),
    .A2(_05625_),
    .B1(_06395_),
    .B2(_06396_),
    .X(_06493_));
 sky130_fd_sc_hd__o21a_2 _14284_ (.A1(_06395_),
    .A2(_06396_),
    .B1(_06493_),
    .X(_06494_));
 sky130_fd_sc_hd__and3_2 _14285_ (.A(net41),
    .B(_05602_),
    .C(_05603_),
    .X(_06495_));
 sky130_fd_sc_hd__or3_2 _14286_ (.A(_05565_),
    .B(_05608_),
    .C(_05609_),
    .X(_06496_));
 sky130_fd_sc_hd__and3_1 _14287_ (.A(net39),
    .B(_05611_),
    .C(_05612_),
    .X(_06497_));
 sky130_fd_sc_hd__xnor2_2 _14288_ (.A(_06496_),
    .B(_06497_),
    .Y(_06498_));
 sky130_fd_sc_hd__xor2_4 _14289_ (.A(_06495_),
    .B(_06498_),
    .X(_06499_));
 sky130_fd_sc_hd__xnor2_2 _14290_ (.A(_06494_),
    .B(_06499_),
    .Y(_06500_));
 sky130_fd_sc_hd__xnor2_4 _14291_ (.A(_06492_),
    .B(_06500_),
    .Y(_06501_));
 sky130_fd_sc_hd__and2_1 _14292_ (.A(_06401_),
    .B(_06406_),
    .X(_06502_));
 sky130_fd_sc_hd__or2_1 _14293_ (.A(_06401_),
    .B(_06406_),
    .X(_06503_));
 sky130_fd_sc_hd__o21ai_2 _14294_ (.A1(_06398_),
    .A2(_06502_),
    .B1(_06503_),
    .Y(_06504_));
 sky130_fd_sc_hd__nor2_1 _14295_ (.A(_06429_),
    .B(_06430_),
    .Y(_06505_));
 sky130_fd_sc_hd__nor2_1 _14296_ (.A(_06425_),
    .B(_06505_),
    .Y(_06506_));
 sky130_fd_sc_hd__nand2_1 _14297_ (.A(_06425_),
    .B(_06505_),
    .Y(_06507_));
 sky130_fd_sc_hd__o31ai_4 _14298_ (.A1(_06427_),
    .A2(_06428_),
    .A3(_06506_),
    .B1(_06507_),
    .Y(_06508_));
 sky130_fd_sc_hd__xor2_2 _14299_ (.A(_06504_),
    .B(_06508_),
    .X(_06509_));
 sky130_fd_sc_hd__xnor2_4 _14300_ (.A(_06501_),
    .B(_06509_),
    .Y(_06510_));
 sky130_fd_sc_hd__nand2_1 _14301_ (.A(_06442_),
    .B(_06443_),
    .Y(_06511_));
 sky130_fd_sc_hd__o22a_1 _14302_ (.A1(_06433_),
    .A2(_06434_),
    .B1(_06511_),
    .B2(_06440_),
    .X(_06512_));
 sky130_fd_sc_hd__a21oi_4 _14303_ (.A1(_06440_),
    .A2(_06511_),
    .B1(_06512_),
    .Y(_06513_));
 sky130_fd_sc_hd__nand2_1 _14304_ (.A(net23),
    .B(_06025_),
    .Y(_06514_));
 sky130_fd_sc_hd__nand2_1 _14305_ (.A(net28),
    .B(net1015),
    .Y(_06515_));
 sky130_fd_sc_hd__xnor2_2 _14306_ (.A(_06514_),
    .B(_06515_),
    .Y(_06516_));
 sky130_fd_sc_hd__nand2_2 _14307_ (.A(net31),
    .B(_05586_),
    .Y(_06517_));
 sky130_fd_sc_hd__nand2_1 _14308_ (.A(net36),
    .B(_05551_),
    .Y(_06518_));
 sky130_fd_sc_hd__nand2_2 _14309_ (.A(net33),
    .B(_05588_),
    .Y(_06519_));
 sky130_fd_sc_hd__xnor2_1 _14310_ (.A(_06518_),
    .B(_06519_),
    .Y(_06520_));
 sky130_fd_sc_hd__xnor2_2 _14311_ (.A(_06517_),
    .B(_06520_),
    .Y(_06521_));
 sky130_fd_sc_hd__o211a_1 _14312_ (.A1(_06437_),
    .A2(_06438_),
    .B1(net30),
    .C1(net1015),
    .X(_06522_));
 sky130_fd_sc_hd__a21o_1 _14313_ (.A1(_06437_),
    .A2(_06438_),
    .B1(_06522_),
    .X(_06523_));
 sky130_fd_sc_hd__o21ba_1 _14314_ (.A1(_06421_),
    .A2(_06423_),
    .B1_N(_06422_),
    .X(_06524_));
 sky130_fd_sc_hd__a21oi_2 _14315_ (.A1(_06421_),
    .A2(_06423_),
    .B1(_06524_),
    .Y(_06525_));
 sky130_fd_sc_hd__xnor2_1 _14316_ (.A(_06523_),
    .B(_06525_),
    .Y(_06526_));
 sky130_fd_sc_hd__xnor2_2 _14317_ (.A(_06521_),
    .B(_06526_),
    .Y(_06527_));
 sky130_fd_sc_hd__xor2_2 _14318_ (.A(_06516_),
    .B(_06527_),
    .X(_06528_));
 sky130_fd_sc_hd__xor2_2 _14319_ (.A(_06513_),
    .B(_06528_),
    .X(_06529_));
 sky130_fd_sc_hd__xnor2_4 _14320_ (.A(_06510_),
    .B(_06529_),
    .Y(_06530_));
 sky130_fd_sc_hd__xor2_1 _14321_ (.A(_06487_),
    .B(_06530_),
    .X(_06531_));
 sky130_fd_sc_hd__xnor2_1 _14322_ (.A(_06481_),
    .B(_06531_),
    .Y(_06532_));
 sky130_fd_sc_hd__nand3_1 _14323_ (.A(net56),
    .B(_06268_),
    .C(_06455_),
    .Y(_06533_));
 sky130_fd_sc_hd__and2b_1 _14324_ (.A_N(_06455_),
    .B(_06456_),
    .X(_06534_));
 sky130_fd_sc_hd__a21o_1 _14325_ (.A1(_06453_),
    .A2(_06533_),
    .B1(_06534_),
    .X(_06535_));
 sky130_fd_sc_hd__clkinvlp_2 _14326_ (.A(_06535_),
    .Y(_06536_));
 sky130_fd_sc_hd__xnor2_1 _14327_ (.A(_06453_),
    .B(_06457_),
    .Y(_06537_));
 sky130_fd_sc_hd__a21o_1 _14328_ (.A1(_06450_),
    .A2(_06451_),
    .B1(_06537_),
    .X(_06538_));
 sky130_fd_sc_hd__and3_1 _14329_ (.A(_06450_),
    .B(_06451_),
    .C(_06537_),
    .X(_06539_));
 sky130_fd_sc_hd__a21oi_1 _14330_ (.A1(_06461_),
    .A2(_06538_),
    .B1(_06539_),
    .Y(_06540_));
 sky130_fd_sc_hd__xnor2_1 _14331_ (.A(_06536_),
    .B(_06540_),
    .Y(_06541_));
 sky130_fd_sc_hd__xnor2_1 _14332_ (.A(_06532_),
    .B(_06541_),
    .Y(_06542_));
 sky130_fd_sc_hd__nor2_1 _14333_ (.A(_06476_),
    .B(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__and2_1 _14334_ (.A(_06476_),
    .B(_06542_),
    .X(_06544_));
 sky130_fd_sc_hd__nor2_4 _14335_ (.A(_06543_),
    .B(_06544_),
    .Y(_06545_));
 sky130_fd_sc_hd__xnor2_4 _14336_ (.A(_06474_),
    .B(_06545_),
    .Y(_06546_));
 sky130_fd_sc_hd__a22o_1 _14337_ (.A1(net855),
    .A2(_06280_),
    .B1(_06546_),
    .B2(_06381_),
    .X(_00022_));
 sky130_fd_sc_hd__nand4bb_4 _14338_ (.A_N(_06178_),
    .B_N(_06384_),
    .C(_06472_),
    .D(_06545_),
    .Y(_06547_));
 sky130_fd_sc_hd__inv_2 _14339_ (.A(_06471_),
    .Y(_06548_));
 sky130_fd_sc_hd__a21oi_1 _14340_ (.A1(_06386_),
    .A2(_06548_),
    .B1(_06470_),
    .Y(_06549_));
 sky130_fd_sc_hd__o21ba_1 _14341_ (.A1(_06549_),
    .A2(_06544_),
    .B1_N(_06543_),
    .X(_06550_));
 sky130_fd_sc_hd__nand2_4 _14342_ (.A(_06547_),
    .B(_06550_),
    .Y(_06551_));
 sky130_fd_sc_hd__a21o_1 _14343_ (.A1(_06484_),
    .A2(_06485_),
    .B1(_06482_),
    .X(_06552_));
 sky130_fd_sc_hd__o21ai_2 _14344_ (.A1(_06484_),
    .A2(_06485_),
    .B1(_06552_),
    .Y(_06553_));
 sky130_fd_sc_hd__inv_1 _14345_ (.A(_06553_),
    .Y(_06554_));
 sky130_fd_sc_hd__a21o_1 _14346_ (.A1(_06487_),
    .A2(_06530_),
    .B1(_06481_),
    .X(_06555_));
 sky130_fd_sc_hd__o21ai_4 _14347_ (.A1(_06487_),
    .A2(_06530_),
    .B1(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__xnor2_2 _14348_ (.A(_06554_),
    .B(_06556_),
    .Y(_06557_));
 sky130_fd_sc_hd__nand2_1 _14349_ (.A(_06513_),
    .B(_06528_),
    .Y(_06558_));
 sky130_fd_sc_hd__nor2_1 _14350_ (.A(_06513_),
    .B(_06528_),
    .Y(_06559_));
 sky130_fd_sc_hd__a21oi_2 _14351_ (.A1(_06510_),
    .A2(_06558_),
    .B1(_06559_),
    .Y(_06560_));
 sky130_fd_sc_hd__nand2_2 _14352_ (.A(net48),
    .B(_06131_),
    .Y(_06561_));
 sky130_fd_sc_hd__and3_1 _14353_ (.A(net44),
    .B(_05723_),
    .C(_05724_),
    .X(_06562_));
 sky130_fd_sc_hd__and3_1 _14354_ (.A(net45),
    .B(_05726_),
    .C(_05727_),
    .X(_06563_));
 sky130_fd_sc_hd__xnor2_2 _14355_ (.A(_06562_),
    .B(_06563_),
    .Y(_06564_));
 sky130_fd_sc_hd__xnor2_4 _14356_ (.A(_06561_),
    .B(_06564_),
    .Y(_06565_));
 sky130_fd_sc_hd__a21bo_1 _14357_ (.A1(_06495_),
    .A2(_06497_),
    .B1_N(_06496_),
    .X(_06566_));
 sky130_fd_sc_hd__o21a_1 _14358_ (.A1(_06495_),
    .A2(_06497_),
    .B1(_06566_),
    .X(_06567_));
 sky130_fd_sc_hd__nand2_2 _14359_ (.A(net39),
    .B(_05605_),
    .Y(_06568_));
 sky130_fd_sc_hd__nand2_1 _14360_ (.A(net41),
    .B(_05625_),
    .Y(_06569_));
 sky130_fd_sc_hd__nand2_1 _14361_ (.A(net36),
    .B(_05639_),
    .Y(_06570_));
 sky130_fd_sc_hd__xor2_1 _14362_ (.A(_06569_),
    .B(_06570_),
    .X(_06571_));
 sky130_fd_sc_hd__xnor2_2 _14363_ (.A(_06568_),
    .B(_06571_),
    .Y(_06572_));
 sky130_fd_sc_hd__xnor2_2 _14364_ (.A(_06567_),
    .B(_06572_),
    .Y(_06573_));
 sky130_fd_sc_hd__xnor2_4 _14365_ (.A(_06565_),
    .B(_06573_),
    .Y(_06574_));
 sky130_fd_sc_hd__a21bo_1 _14366_ (.A1(_06494_),
    .A2(_06499_),
    .B1_N(_06492_),
    .X(_06575_));
 sky130_fd_sc_hd__o21ai_2 _14367_ (.A1(_06494_),
    .A2(_06499_),
    .B1(_06575_),
    .Y(_06576_));
 sky130_fd_sc_hd__nand2_1 _14368_ (.A(_06523_),
    .B(_06525_),
    .Y(_06577_));
 sky130_fd_sc_hd__nor2_1 _14369_ (.A(_06523_),
    .B(_06525_),
    .Y(_06578_));
 sky130_fd_sc_hd__a21o_1 _14370_ (.A1(_06521_),
    .A2(_06577_),
    .B1(_06578_),
    .X(_06579_));
 sky130_fd_sc_hd__xnor2_2 _14371_ (.A(_06576_),
    .B(_06579_),
    .Y(_06580_));
 sky130_fd_sc_hd__xnor2_4 _14372_ (.A(_06574_),
    .B(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__nor2_1 _14373_ (.A(_06516_),
    .B(_06527_),
    .Y(_06582_));
 sky130_fd_sc_hd__nor2_2 _14374_ (.A(_06217_),
    .B(_05822_),
    .Y(_06583_));
 sky130_fd_sc_hd__nand2_1 _14375_ (.A(net33),
    .B(_05551_),
    .Y(_06584_));
 sky130_fd_sc_hd__nand2_1 _14376_ (.A(net30),
    .B(_05588_),
    .Y(_06585_));
 sky130_fd_sc_hd__xnor2_2 _14377_ (.A(_06584_),
    .B(_06585_),
    .Y(_06586_));
 sky130_fd_sc_hd__xnor2_4 _14378_ (.A(_06583_),
    .B(_06586_),
    .Y(_06587_));
 sky130_fd_sc_hd__o21a_1 _14379_ (.A1(_06517_),
    .A2(_06519_),
    .B1(_06518_),
    .X(_06588_));
 sky130_fd_sc_hd__a21oi_4 _14380_ (.A1(_06517_),
    .A2(_06519_),
    .B1(_06588_),
    .Y(_06589_));
 sky130_fd_sc_hd__xnor2_4 _14381_ (.A(_06587_),
    .B(_06589_),
    .Y(_06590_));
 sky130_fd_sc_hd__and3b_1 _14382_ (.A_N(_06437_),
    .B(net1015),
    .C(net23),
    .X(_06591_));
 sky130_fd_sc_hd__xor2_4 _14383_ (.A(_06590_),
    .B(_06591_),
    .X(_06592_));
 sky130_fd_sc_hd__xnor2_1 _14384_ (.A(_06582_),
    .B(_06592_),
    .Y(_06593_));
 sky130_fd_sc_hd__xnor2_2 _14385_ (.A(_06581_),
    .B(_06593_),
    .Y(_06594_));
 sky130_fd_sc_hd__a22o_1 _14386_ (.A1(net51),
    .A2(_06351_),
    .B1(_06489_),
    .B2(_06490_),
    .X(_06595_));
 sky130_fd_sc_hd__o21a_1 _14387_ (.A1(_06489_),
    .A2(_06490_),
    .B1(_06595_),
    .X(_06596_));
 sky130_fd_sc_hd__nand2_1 _14388_ (.A(net51),
    .B(_06268_),
    .Y(_06597_));
 sky130_fd_sc_hd__xnor2_1 _14389_ (.A(_06596_),
    .B(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__a21boi_1 _14390_ (.A1(_06501_),
    .A2(_06504_),
    .B1_N(_06508_),
    .Y(_06599_));
 sky130_fd_sc_hd__o21ba_1 _14391_ (.A1(_06501_),
    .A2(_06504_),
    .B1_N(_06599_),
    .X(_06600_));
 sky130_fd_sc_hd__xnor2_1 _14392_ (.A(_06598_),
    .B(_06600_),
    .Y(_06601_));
 sky130_fd_sc_hd__xnor2_1 _14393_ (.A(_06594_),
    .B(_06601_),
    .Y(_06602_));
 sky130_fd_sc_hd__xnor2_1 _14394_ (.A(_06560_),
    .B(_06602_),
    .Y(_06603_));
 sky130_fd_sc_hd__xnor2_1 _14395_ (.A(_06481_),
    .B(_06487_),
    .Y(_06604_));
 sky130_fd_sc_hd__nor3_1 _14396_ (.A(_06535_),
    .B(_06530_),
    .C(_06604_),
    .Y(_06605_));
 sky130_fd_sc_hd__a311o_1 _14397_ (.A1(_06536_),
    .A2(_06530_),
    .A3(_06604_),
    .B1(_06605_),
    .C1(_06540_),
    .X(_06606_));
 sky130_fd_sc_hd__a21boi_1 _14398_ (.A1(_06535_),
    .A2(_06532_),
    .B1_N(_06606_),
    .Y(_06607_));
 sky130_fd_sc_hd__and2_1 _14399_ (.A(_06603_),
    .B(_06607_),
    .X(_06608_));
 sky130_fd_sc_hd__nor2_1 _14400_ (.A(_06603_),
    .B(_06607_),
    .Y(_06609_));
 sky130_fd_sc_hd__or2_1 _14401_ (.A(_06608_),
    .B(_06609_),
    .X(_06610_));
 sky130_fd_sc_hd__xor2_2 _14402_ (.A(_06557_),
    .B(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__xnor2_4 _14403_ (.A(_06551_),
    .B(_06611_),
    .Y(_06612_));
 sky130_fd_sc_hd__a22o_1 _14404_ (.A1(net869),
    .A2(_06280_),
    .B1(_06612_),
    .B2(_06381_),
    .X(_00023_));
 sky130_fd_sc_hd__o21ba_1 _14405_ (.A1(_06581_),
    .A2(_06592_),
    .B1_N(_06582_),
    .X(_06613_));
 sky130_fd_sc_hd__a21oi_4 _14406_ (.A1(_06581_),
    .A2(_06592_),
    .B1(_06613_),
    .Y(_06614_));
 sky130_fd_sc_hd__nand2_2 _14407_ (.A(net45),
    .B(_06131_),
    .Y(_06615_));
 sky130_fd_sc_hd__nand2_2 _14408_ (.A(net41),
    .B(_05619_),
    .Y(_06616_));
 sky130_fd_sc_hd__nand2_2 _14409_ (.A(net44),
    .B(_05666_),
    .Y(_06617_));
 sky130_fd_sc_hd__xnor2_2 _14410_ (.A(_06616_),
    .B(_06617_),
    .Y(_06618_));
 sky130_fd_sc_hd__xnor2_4 _14411_ (.A(_06615_),
    .B(_06618_),
    .Y(_06619_));
 sky130_fd_sc_hd__nand2_1 _14412_ (.A(_06568_),
    .B(_06570_),
    .Y(_06620_));
 sky130_fd_sc_hd__nor2_1 _14413_ (.A(_06568_),
    .B(_06570_),
    .Y(_06621_));
 sky130_fd_sc_hd__a31o_1 _14414_ (.A1(net41),
    .A2(_05625_),
    .A3(_06620_),
    .B1(_06621_),
    .X(_06622_));
 sky130_fd_sc_hd__and3_2 _14415_ (.A(net36),
    .B(_05602_),
    .C(_05603_),
    .X(_06623_));
 sky130_fd_sc_hd__nand2_1 _14416_ (.A(net39),
    .B(_05625_),
    .Y(_06624_));
 sky130_fd_sc_hd__nor2_1 _14417_ (.A(_05500_),
    .B(_05731_),
    .Y(_06625_));
 sky130_fd_sc_hd__xor2_1 _14418_ (.A(_06624_),
    .B(_06625_),
    .X(_06626_));
 sky130_fd_sc_hd__xnor2_2 _14419_ (.A(_06623_),
    .B(_06626_),
    .Y(_06627_));
 sky130_fd_sc_hd__xnor2_2 _14420_ (.A(_06622_),
    .B(_06627_),
    .Y(_06628_));
 sky130_fd_sc_hd__xnor2_4 _14421_ (.A(_06619_),
    .B(_06628_),
    .Y(_06629_));
 sky130_fd_sc_hd__nor2_1 _14422_ (.A(_06567_),
    .B(_06572_),
    .Y(_06630_));
 sky130_fd_sc_hd__nand2_1 _14423_ (.A(_06567_),
    .B(_06572_),
    .Y(_06631_));
 sky130_fd_sc_hd__o21a_2 _14424_ (.A1(_06565_),
    .A2(_06630_),
    .B1(_06631_),
    .X(_06632_));
 sky130_fd_sc_hd__a32o_1 _14425_ (.A1(_06025_),
    .A2(net1015),
    .A3(_06320_),
    .B1(_06587_),
    .B2(_06589_),
    .X(_06633_));
 sky130_fd_sc_hd__o21a_1 _14426_ (.A1(_06587_),
    .A2(_06589_),
    .B1(_06633_),
    .X(_06634_));
 sky130_fd_sc_hd__xor2_2 _14427_ (.A(_06632_),
    .B(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__xnor2_4 _14428_ (.A(_06629_),
    .B(_06635_),
    .Y(_06636_));
 sky130_fd_sc_hd__xnor2_1 _14429_ (.A(_06437_),
    .B(_06590_),
    .Y(_06637_));
 sky130_fd_sc_hd__nand3_2 _14430_ (.A(net23),
    .B(net1015),
    .C(_06637_),
    .Y(_06638_));
 sky130_fd_sc_hd__or2b_1 _14431_ (.A(_06583_),
    .B_N(_06585_),
    .X(_06639_));
 sky130_fd_sc_hd__buf_2 _14432_ (.A(_05588_),
    .X(_06640_));
 sky130_fd_sc_hd__a32o_1 _14433_ (.A1(net30),
    .A2(_06640_),
    .A3(_06583_),
    .B1(_05579_),
    .B2(net33),
    .X(_06641_));
 sky130_fd_sc_hd__nand2_1 _14434_ (.A(_06639_),
    .B(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__nand2_1 _14435_ (.A(net28),
    .B(_06640_),
    .Y(_06643_));
 sky130_fd_sc_hd__nand2_1 _14436_ (.A(net23),
    .B(_05586_),
    .Y(_06644_));
 sky130_fd_sc_hd__nand2_1 _14437_ (.A(net30),
    .B(_05579_),
    .Y(_06645_));
 sky130_fd_sc_hd__xnor2_1 _14438_ (.A(_06644_),
    .B(_06645_),
    .Y(_06646_));
 sky130_fd_sc_hd__xnor2_1 _14439_ (.A(_06643_),
    .B(_06646_),
    .Y(_06647_));
 sky130_fd_sc_hd__and2_1 _14440_ (.A(_06642_),
    .B(_06647_),
    .X(_06648_));
 sky130_fd_sc_hd__nor2_1 _14441_ (.A(_06642_),
    .B(_06647_),
    .Y(_06649_));
 sky130_fd_sc_hd__or2_2 _14442_ (.A(_06648_),
    .B(_06649_),
    .X(_06650_));
 sky130_fd_sc_hd__xor2_2 _14443_ (.A(_06638_),
    .B(_06650_),
    .X(_06651_));
 sky130_fd_sc_hd__xnor2_4 _14444_ (.A(_06636_),
    .B(_06651_),
    .Y(_06652_));
 sky130_fd_sc_hd__a21o_1 _14445_ (.A1(_06574_),
    .A2(_06579_),
    .B1(_06576_),
    .X(_06653_));
 sky130_fd_sc_hd__o21ai_2 _14446_ (.A1(_06574_),
    .A2(_06579_),
    .B1(_06653_),
    .Y(_06654_));
 sky130_fd_sc_hd__a22o_1 _14447_ (.A1(net49),
    .A2(_06131_),
    .B1(_06562_),
    .B2(_06563_),
    .X(_06655_));
 sky130_fd_sc_hd__o21a_1 _14448_ (.A1(_06562_),
    .A2(_06563_),
    .B1(_06655_),
    .X(_06656_));
 sky130_fd_sc_hd__and2_1 _14449_ (.A(net49),
    .B(_06135_),
    .X(_06657_));
 sky130_fd_sc_hd__xor2_1 _14450_ (.A(_06656_),
    .B(_06657_),
    .X(_06658_));
 sky130_fd_sc_hd__xnor2_2 _14451_ (.A(_06654_),
    .B(_06658_),
    .Y(_06659_));
 sky130_fd_sc_hd__xor2_2 _14452_ (.A(_06652_),
    .B(_06659_),
    .X(_06660_));
 sky130_fd_sc_hd__xnor2_4 _14453_ (.A(_06614_),
    .B(_06660_),
    .Y(_06661_));
 sky130_fd_sc_hd__nand2_2 _14454_ (.A(_06597_),
    .B(_06600_),
    .Y(_06662_));
 sky130_fd_sc_hd__or2_1 _14455_ (.A(_06596_),
    .B(_06594_),
    .X(_06663_));
 sky130_fd_sc_hd__nor2_1 _14456_ (.A(_06597_),
    .B(_06600_),
    .Y(_06664_));
 sky130_fd_sc_hd__and2_1 _14457_ (.A(_06596_),
    .B(_06594_),
    .X(_06665_));
 sky130_fd_sc_hd__o22a_1 _14458_ (.A1(_06663_),
    .A2(_06664_),
    .B1(_06665_),
    .B2(_06662_),
    .X(_06666_));
 sky130_fd_sc_hd__o211a_1 _14459_ (.A1(_06596_),
    .A2(_06664_),
    .B1(_06662_),
    .C1(_06560_),
    .X(_06667_));
 sky130_fd_sc_hd__and3_1 _14460_ (.A(_06596_),
    .B(_06594_),
    .C(_06664_),
    .X(_06668_));
 sky130_fd_sc_hd__a21o_1 _14461_ (.A1(_06596_),
    .A2(_06664_),
    .B1(_06594_),
    .X(_06669_));
 sky130_fd_sc_hd__o21ai_1 _14462_ (.A1(_06667_),
    .A2(_06668_),
    .B1(_06669_),
    .Y(_06670_));
 sky130_fd_sc_hd__o221a_2 _14463_ (.A1(_06662_),
    .A2(_06663_),
    .B1(_06666_),
    .B2(_06560_),
    .C1(_06670_),
    .X(_06671_));
 sky130_fd_sc_hd__xor2_4 _14464_ (.A(_06661_),
    .B(_06671_),
    .X(_06672_));
 sky130_fd_sc_hd__nor2_2 _14465_ (.A(_06553_),
    .B(_06556_),
    .Y(_06673_));
 sky130_fd_sc_hd__nand2_1 _14466_ (.A(_06553_),
    .B(_06556_),
    .Y(_06674_));
 sky130_fd_sc_hd__inv_2 _14467_ (.A(_06674_),
    .Y(_06675_));
 sky130_fd_sc_hd__o21ba_1 _14468_ (.A1(_06554_),
    .A2(_06608_),
    .B1_N(_06609_),
    .X(_06676_));
 sky130_fd_sc_hd__clkinvlp_2 _14469_ (.A(_06556_),
    .Y(_06677_));
 sky130_fd_sc_hd__a2bb2o_1 _14470_ (.A1_N(_06676_),
    .A2_N(_06677_),
    .B1(_06553_),
    .B2(_06609_),
    .X(_06678_));
 sky130_fd_sc_hd__a22o_1 _14471_ (.A1(_06554_),
    .A2(_06608_),
    .B1(_06676_),
    .B2(_06677_),
    .X(_06679_));
 sky130_fd_sc_hd__mux2_1 _14472_ (.A0(_06678_),
    .A1(_06679_),
    .S(_06551_),
    .X(_06680_));
 sky130_fd_sc_hd__a221o_2 _14473_ (.A1(_06608_),
    .A2(_06673_),
    .B1(_06675_),
    .B2(_06609_),
    .C1(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__xnor2_4 _14474_ (.A(_06672_),
    .B(_06681_),
    .Y(_06682_));
 sky130_fd_sc_hd__a22o_1 _14475_ (.A1(net864),
    .A2(_06280_),
    .B1(_06682_),
    .B2(_06381_),
    .X(_00024_));
 sky130_fd_sc_hd__o221a_1 _14476_ (.A1(_06554_),
    .A2(_06677_),
    .B1(_06603_),
    .B2(_06607_),
    .C1(_06672_),
    .X(_06683_));
 sky130_fd_sc_hd__o21a_1 _14477_ (.A1(_06672_),
    .A2(_06673_),
    .B1(_06608_),
    .X(_06684_));
 sky130_fd_sc_hd__a211oi_2 _14478_ (.A1(_06672_),
    .A2(_06673_),
    .B1(_06683_),
    .C1(_06684_),
    .Y(_06685_));
 sky130_fd_sc_hd__mux2_1 _14479_ (.A0(_06608_),
    .A1(_06609_),
    .S(_06672_),
    .X(_06686_));
 sky130_fd_sc_hd__inv_2 _14480_ (.A(_06673_),
    .Y(_06687_));
 sky130_fd_sc_hd__mux2_1 _14481_ (.A0(_06687_),
    .A1(_06674_),
    .S(_06672_),
    .X(_06688_));
 sky130_fd_sc_hd__o2bb2a_1 _14482_ (.A1_N(_06557_),
    .A2_N(_06686_),
    .B1(_06688_),
    .B2(_06610_),
    .X(_06689_));
 sky130_fd_sc_hd__a21o_1 _14483_ (.A1(_06547_),
    .A2(_06550_),
    .B1(_06689_),
    .X(_06690_));
 sky130_fd_sc_hd__and2_2 _14484_ (.A(_06685_),
    .B(_06690_),
    .X(_06691_));
 sky130_fd_sc_hd__a21o_1 _14485_ (.A1(_06560_),
    .A2(_06663_),
    .B1(_06665_),
    .X(_06692_));
 sky130_fd_sc_hd__a21oi_1 _14486_ (.A1(_06661_),
    .A2(_06692_),
    .B1(_06664_),
    .Y(_06693_));
 sky130_fd_sc_hd__nor2_1 _14487_ (.A(_06661_),
    .B(_06692_),
    .Y(_06694_));
 sky130_fd_sc_hd__o211a_1 _14488_ (.A1(_06661_),
    .A2(_06665_),
    .B1(_06662_),
    .C1(_06560_),
    .X(_06695_));
 sky130_fd_sc_hd__a31oi_2 _14489_ (.A1(_06661_),
    .A2(_06662_),
    .A3(_06663_),
    .B1(_06695_),
    .Y(_06696_));
 sky130_fd_sc_hd__o21ai_4 _14490_ (.A1(_06693_),
    .A2(_06694_),
    .B1(_06696_),
    .Y(_06697_));
 sky130_fd_sc_hd__o21a_1 _14491_ (.A1(_06636_),
    .A2(_06650_),
    .B1(_06638_),
    .X(_06698_));
 sky130_fd_sc_hd__a21oi_4 _14492_ (.A1(_06636_),
    .A2(_06650_),
    .B1(_06698_),
    .Y(_06699_));
 sky130_fd_sc_hd__nand2_1 _14493_ (.A(net44),
    .B(_06131_),
    .Y(_06700_));
 sky130_fd_sc_hd__and3_1 _14494_ (.A(net39),
    .B(_05723_),
    .C(_05724_),
    .X(_06701_));
 sky130_fd_sc_hd__and3_1 _14495_ (.A(net41),
    .B(_05726_),
    .C(_05727_),
    .X(_06702_));
 sky130_fd_sc_hd__xnor2_1 _14496_ (.A(_06701_),
    .B(_06702_),
    .Y(_06703_));
 sky130_fd_sc_hd__xnor2_1 _14497_ (.A(_06700_),
    .B(_06703_),
    .Y(_06704_));
 sky130_fd_sc_hd__a21bo_1 _14498_ (.A1(_06623_),
    .A2(_06625_),
    .B1_N(_06624_),
    .X(_06705_));
 sky130_fd_sc_hd__o21a_1 _14499_ (.A1(_06623_),
    .A2(_06625_),
    .B1(_06705_),
    .X(_06706_));
 sky130_fd_sc_hd__nand2_2 _14500_ (.A(net33),
    .B(_05605_),
    .Y(_06707_));
 sky130_fd_sc_hd__nand2_1 _14501_ (.A(net36),
    .B(_05625_),
    .Y(_06708_));
 sky130_fd_sc_hd__nand2_2 _14502_ (.A(net31),
    .B(_05639_),
    .Y(_06709_));
 sky130_fd_sc_hd__xor2_2 _14503_ (.A(_06708_),
    .B(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__xnor2_2 _14504_ (.A(_06707_),
    .B(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__xnor2_1 _14505_ (.A(_06706_),
    .B(_06711_),
    .Y(_06712_));
 sky130_fd_sc_hd__xnor2_1 _14506_ (.A(_06704_),
    .B(_06712_),
    .Y(_06713_));
 sky130_fd_sc_hd__xnor2_1 _14507_ (.A(_06649_),
    .B(_06713_),
    .Y(_06714_));
 sky130_fd_sc_hd__nand2_1 _14508_ (.A(_05579_),
    .B(_06640_),
    .Y(_06715_));
 sky130_fd_sc_hd__nor2_1 _14509_ (.A(_06212_),
    .B(_06715_),
    .Y(_06716_));
 sky130_fd_sc_hd__o2bb2a_1 _14510_ (.A1_N(_05822_),
    .A2_N(_06716_),
    .B1(_06640_),
    .B2(net28),
    .X(_06717_));
 sky130_fd_sc_hd__o22a_1 _14511_ (.A1(_06640_),
    .A2(_06212_),
    .B1(_06715_),
    .B2(net25),
    .X(_06718_));
 sky130_fd_sc_hd__o22a_1 _14512_ (.A1(_06217_),
    .A2(_05579_),
    .B1(_06718_),
    .B2(_06106_),
    .X(_06719_));
 sky130_fd_sc_hd__o21a_1 _14513_ (.A1(_05586_),
    .A2(_06640_),
    .B1(net23),
    .X(_06720_));
 sky130_fd_sc_hd__a21o_1 _14514_ (.A1(_05579_),
    .A2(_06585_),
    .B1(net23),
    .X(_06721_));
 sky130_fd_sc_hd__o221a_1 _14515_ (.A1(_05579_),
    .A2(_06640_),
    .B1(_06720_),
    .B2(net28),
    .C1(_06721_),
    .X(_06722_));
 sky130_fd_sc_hd__o221a_1 _14516_ (.A1(net30),
    .A2(_06717_),
    .B1(_06719_),
    .B2(_05822_),
    .C1(_06722_),
    .X(_06723_));
 sky130_fd_sc_hd__a21bo_1 _14517_ (.A1(_06622_),
    .A2(_06627_),
    .B1_N(_06619_),
    .X(_06724_));
 sky130_fd_sc_hd__o21a_1 _14518_ (.A1(_06622_),
    .A2(_06627_),
    .B1(_06724_),
    .X(_06725_));
 sky130_fd_sc_hd__xor2_1 _14519_ (.A(_06723_),
    .B(_06725_),
    .X(_06726_));
 sky130_fd_sc_hd__xnor2_1 _14520_ (.A(_06714_),
    .B(_06726_),
    .Y(_06727_));
 sky130_fd_sc_hd__a21bo_1 _14521_ (.A1(_06629_),
    .A2(_06632_),
    .B1_N(_06634_),
    .X(_06728_));
 sky130_fd_sc_hd__o21ai_2 _14522_ (.A1(_06629_),
    .A2(_06632_),
    .B1(_06728_),
    .Y(_06729_));
 sky130_fd_sc_hd__nand2_1 _14523_ (.A(_06616_),
    .B(_06617_),
    .Y(_06730_));
 sky130_fd_sc_hd__nor2_1 _14524_ (.A(_06616_),
    .B(_06617_),
    .Y(_06731_));
 sky130_fd_sc_hd__a31o_1 _14525_ (.A1(net45),
    .A2(_06351_),
    .A3(_06730_),
    .B1(_06731_),
    .X(_06732_));
 sky130_fd_sc_hd__nand2_1 _14526_ (.A(net45),
    .B(_06268_),
    .Y(_06733_));
 sky130_fd_sc_hd__xnor2_1 _14527_ (.A(_06732_),
    .B(_06733_),
    .Y(_06734_));
 sky130_fd_sc_hd__xnor2_1 _14528_ (.A(_06729_),
    .B(_06734_),
    .Y(_06735_));
 sky130_fd_sc_hd__nand2_1 _14529_ (.A(_06727_),
    .B(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__inv_2 _14530_ (.A(_06736_),
    .Y(_06737_));
 sky130_fd_sc_hd__nor2_1 _14531_ (.A(_06727_),
    .B(_06735_),
    .Y(_06738_));
 sky130_fd_sc_hd__nor2_2 _14532_ (.A(_06737_),
    .B(_06738_),
    .Y(_06739_));
 sky130_fd_sc_hd__xnor2_4 _14533_ (.A(_06699_),
    .B(_06739_),
    .Y(_06740_));
 sky130_fd_sc_hd__a21o_1 _14534_ (.A1(_06656_),
    .A2(_06657_),
    .B1(_06654_),
    .X(_06741_));
 sky130_fd_sc_hd__o21ai_4 _14535_ (.A1(_06656_),
    .A2(_06657_),
    .B1(_06741_),
    .Y(_06742_));
 sky130_fd_sc_hd__a21bo_1 _14536_ (.A1(_06652_),
    .A2(_06614_),
    .B1_N(_06659_),
    .X(_06743_));
 sky130_fd_sc_hd__o21ai_4 _14537_ (.A1(_06652_),
    .A2(_06614_),
    .B1(_06743_),
    .Y(_06744_));
 sky130_fd_sc_hd__xnor2_2 _14538_ (.A(_06742_),
    .B(_06744_),
    .Y(_06745_));
 sky130_fd_sc_hd__xor2_2 _14539_ (.A(_06740_),
    .B(_06745_),
    .X(_06746_));
 sky130_fd_sc_hd__xor2_2 _14540_ (.A(_06697_),
    .B(_06746_),
    .X(_06747_));
 sky130_fd_sc_hd__xnor2_4 _14541_ (.A(_06691_),
    .B(_06747_),
    .Y(_06748_));
 sky130_fd_sc_hd__a22o_1 _14542_ (.A1(net861),
    .A2(_06280_),
    .B1(_06748_),
    .B2(_06381_),
    .X(_00025_));
 sky130_fd_sc_hd__a21o_2 _14543_ (.A1(_06699_),
    .A2(_06736_),
    .B1(_06738_),
    .X(_06749_));
 sky130_fd_sc_hd__a21bo_1 _14544_ (.A1(_06729_),
    .A2(_06732_),
    .B1_N(_06733_),
    .X(_06750_));
 sky130_fd_sc_hd__o21a_2 _14545_ (.A1(_06729_),
    .A2(_06732_),
    .B1(_06750_),
    .X(_06751_));
 sky130_fd_sc_hd__a21bo_1 _14546_ (.A1(_06649_),
    .A2(_06725_),
    .B1_N(_06713_),
    .X(_06752_));
 sky130_fd_sc_hd__o21a_2 _14547_ (.A1(_06649_),
    .A2(_06725_),
    .B1(_06752_),
    .X(_06753_));
 sky130_fd_sc_hd__a22o_1 _14548_ (.A1(net44),
    .A2(_06351_),
    .B1(_06701_),
    .B2(_06702_),
    .X(_06754_));
 sky130_fd_sc_hd__o21a_1 _14549_ (.A1(_06701_),
    .A2(_06702_),
    .B1(_06754_),
    .X(_06755_));
 sky130_fd_sc_hd__and2_1 _14550_ (.A(net44),
    .B(_06268_),
    .X(_06756_));
 sky130_fd_sc_hd__xnor2_2 _14551_ (.A(_06755_),
    .B(_06756_),
    .Y(_06757_));
 sky130_fd_sc_hd__xnor2_4 _14552_ (.A(_06753_),
    .B(_06757_),
    .Y(_06758_));
 sky130_fd_sc_hd__and3_1 _14553_ (.A(net23),
    .B(_05579_),
    .C(_06643_),
    .X(_06759_));
 sky130_fd_sc_hd__nand2_2 _14554_ (.A(net30),
    .B(_05605_),
    .Y(_06760_));
 sky130_fd_sc_hd__nand2_1 _14555_ (.A(net33),
    .B(_05626_),
    .Y(_06761_));
 sky130_fd_sc_hd__nand2_1 _14556_ (.A(net25),
    .B(_05640_),
    .Y(_06762_));
 sky130_fd_sc_hd__xor2_1 _14557_ (.A(_06761_),
    .B(_06762_),
    .X(_06763_));
 sky130_fd_sc_hd__xnor2_2 _14558_ (.A(_06760_),
    .B(_06763_),
    .Y(_06764_));
 sky130_fd_sc_hd__o21a_1 _14559_ (.A1(_06707_),
    .A2(_06709_),
    .B1(_06708_),
    .X(_06765_));
 sky130_fd_sc_hd__a21o_1 _14560_ (.A1(_06707_),
    .A2(_06709_),
    .B1(_06765_),
    .X(_06766_));
 sky130_fd_sc_hd__nand2_1 _14561_ (.A(net41),
    .B(_06131_),
    .Y(_06767_));
 sky130_fd_sc_hd__and3_1 _14562_ (.A(net36),
    .B(_05723_),
    .C(_05724_),
    .X(_06768_));
 sky130_fd_sc_hd__and3_1 _14563_ (.A(net39),
    .B(_05726_),
    .C(_05727_),
    .X(_06769_));
 sky130_fd_sc_hd__xnor2_1 _14564_ (.A(_06768_),
    .B(_06769_),
    .Y(_06770_));
 sky130_fd_sc_hd__xnor2_2 _14565_ (.A(_06767_),
    .B(_06770_),
    .Y(_06771_));
 sky130_fd_sc_hd__xor2_1 _14566_ (.A(_06766_),
    .B(_06771_),
    .X(_06772_));
 sky130_fd_sc_hd__xnor2_2 _14567_ (.A(_06764_),
    .B(_06772_),
    .Y(_06773_));
 sky130_fd_sc_hd__a21bo_1 _14568_ (.A1(_06706_),
    .A2(_06711_),
    .B1_N(_06704_),
    .X(_06774_));
 sky130_fd_sc_hd__o21a_1 _14569_ (.A1(_06706_),
    .A2(_06711_),
    .B1(_06774_),
    .X(_06775_));
 sky130_fd_sc_hd__nand2_1 _14570_ (.A(_05586_),
    .B(_06640_),
    .Y(_06776_));
 sky130_fd_sc_hd__inv_2 _14571_ (.A(_06323_),
    .Y(_06777_));
 sky130_fd_sc_hd__nor2_1 _14572_ (.A(_05822_),
    .B(_06640_),
    .Y(_06778_));
 sky130_fd_sc_hd__mux2_1 _14573_ (.A0(_06640_),
    .A1(_06778_),
    .S(net23),
    .X(_06779_));
 sky130_fd_sc_hd__a2bb2o_1 _14574_ (.A1_N(_06776_),
    .A2_N(_06777_),
    .B1(_06779_),
    .B2(net28),
    .X(_06780_));
 sky130_fd_sc_hd__inv_2 _14575_ (.A(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__o32a_1 _14576_ (.A1(_05579_),
    .A2(_06776_),
    .A3(_06212_),
    .B1(_06645_),
    .B2(_06781_),
    .X(_06782_));
 sky130_fd_sc_hd__xnor2_1 _14577_ (.A(_06775_),
    .B(_06782_),
    .Y(_06783_));
 sky130_fd_sc_hd__xnor2_2 _14578_ (.A(_06773_),
    .B(_06783_),
    .Y(_06784_));
 sky130_fd_sc_hd__xor2_2 _14579_ (.A(_06759_),
    .B(_06784_),
    .X(_06785_));
 sky130_fd_sc_hd__nand2_1 _14580_ (.A(_06714_),
    .B(_06725_),
    .Y(_06786_));
 sky130_fd_sc_hd__or2_1 _14581_ (.A(_06714_),
    .B(_06725_),
    .X(_06787_));
 sky130_fd_sc_hd__and3_1 _14582_ (.A(_06723_),
    .B(_06786_),
    .C(_06787_),
    .X(_06788_));
 sky130_fd_sc_hd__xnor2_2 _14583_ (.A(_06785_),
    .B(_06788_),
    .Y(_06789_));
 sky130_fd_sc_hd__xnor2_4 _14584_ (.A(_06758_),
    .B(_06789_),
    .Y(_06790_));
 sky130_fd_sc_hd__xnor2_4 _14585_ (.A(_06751_),
    .B(_06790_),
    .Y(_06791_));
 sky130_fd_sc_hd__xor2_4 _14586_ (.A(_06749_),
    .B(_06791_),
    .X(_06792_));
 sky130_fd_sc_hd__or2_1 _14587_ (.A(_06742_),
    .B(_06744_),
    .X(_06793_));
 sky130_fd_sc_hd__and2_1 _14588_ (.A(_06742_),
    .B(_06744_),
    .X(_06794_));
 sky130_fd_sc_hd__a21o_1 _14589_ (.A1(_06740_),
    .A2(_06793_),
    .B1(_06794_),
    .X(_06795_));
 sky130_fd_sc_hd__xnor2_2 _14590_ (.A(_06792_),
    .B(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__o21ba_1 _14591_ (.A1(_06697_),
    .A2(_06746_),
    .B1_N(_06691_),
    .X(_06797_));
 sky130_fd_sc_hd__a21o_1 _14592_ (.A1(_06697_),
    .A2(_06746_),
    .B1(_06797_),
    .X(_06798_));
 sky130_fd_sc_hd__xnor2_4 _14593_ (.A(_06796_),
    .B(_06798_),
    .Y(_06799_));
 sky130_fd_sc_hd__a22o_1 _14594_ (.A1(net810),
    .A2(_06280_),
    .B1(_06799_),
    .B2(_06381_),
    .X(_00026_));
 sky130_fd_sc_hd__xnor2_2 _14595_ (.A(_06749_),
    .B(_06791_),
    .Y(_06800_));
 sky130_fd_sc_hd__nor2_1 _14596_ (.A(_06800_),
    .B(_06793_),
    .Y(_06801_));
 sky130_fd_sc_hd__a21oi_1 _14597_ (.A1(_06800_),
    .A2(_06794_),
    .B1(_06801_),
    .Y(_06802_));
 sky130_fd_sc_hd__xor2_1 _14598_ (.A(_06697_),
    .B(_06740_),
    .X(_06803_));
 sky130_fd_sc_hd__or4b_1 _14599_ (.A(_06740_),
    .B(_06745_),
    .C(_06800_),
    .D_N(_06697_),
    .X(_06804_));
 sky130_fd_sc_hd__or4b_1 _14600_ (.A(_06697_),
    .B(_06792_),
    .C(_06745_),
    .D_N(_06740_),
    .X(_06805_));
 sky130_fd_sc_hd__o211a_1 _14601_ (.A1(_06802_),
    .A2(_06803_),
    .B1(_06804_),
    .C1(_06805_),
    .X(_06806_));
 sky130_fd_sc_hd__nor2_1 _14602_ (.A(_06689_),
    .B(_06806_),
    .Y(_06807_));
 sky130_fd_sc_hd__and2_1 _14603_ (.A(_06685_),
    .B(_06744_),
    .X(_06808_));
 sky130_fd_sc_hd__nor2_1 _14604_ (.A(_06740_),
    .B(_06742_),
    .Y(_06809_));
 sky130_fd_sc_hd__nand2_1 _14605_ (.A(_06740_),
    .B(_06742_),
    .Y(_06810_));
 sky130_fd_sc_hd__o21ai_1 _14606_ (.A1(_06697_),
    .A2(_06809_),
    .B1(_06810_),
    .Y(_06811_));
 sky130_fd_sc_hd__o21a_1 _14607_ (.A1(_06792_),
    .A2(_06808_),
    .B1(_06811_),
    .X(_06812_));
 sky130_fd_sc_hd__a21oi_1 _14608_ (.A1(_06800_),
    .A2(_06810_),
    .B1(_06697_),
    .Y(_06813_));
 sky130_fd_sc_hd__nor2_1 _14609_ (.A(_06800_),
    .B(_06809_),
    .Y(_06814_));
 sky130_fd_sc_hd__o22a_1 _14610_ (.A1(_06685_),
    .A2(_06744_),
    .B1(_06813_),
    .B2(_06814_),
    .X(_06815_));
 sky130_fd_sc_hd__a211oi_1 _14611_ (.A1(_06792_),
    .A2(_06808_),
    .B1(_06812_),
    .C1(_06815_),
    .Y(_06816_));
 sky130_fd_sc_hd__a21o_1 _14612_ (.A1(_06551_),
    .A2(_06807_),
    .B1(_06816_),
    .X(_06817_));
 sky130_fd_sc_hd__o21a_1 _14613_ (.A1(_06751_),
    .A2(_06790_),
    .B1(_06749_),
    .X(_06818_));
 sky130_fd_sc_hd__a21o_1 _14614_ (.A1(_06751_),
    .A2(_06790_),
    .B1(_06818_),
    .X(_06819_));
 sky130_fd_sc_hd__and2_1 _14615_ (.A(_06759_),
    .B(_06784_),
    .X(_06820_));
 sky130_fd_sc_hd__and2b_1 _14616_ (.A_N(_06775_),
    .B(_06782_),
    .X(_06821_));
 sky130_fd_sc_hd__or2b_1 _14617_ (.A(_06782_),
    .B_N(_06775_),
    .X(_06822_));
 sky130_fd_sc_hd__o21ai_2 _14618_ (.A1(_06773_),
    .A2(_06821_),
    .B1(_06822_),
    .Y(_06823_));
 sky130_fd_sc_hd__buf_6 _14619_ (.A(_06351_),
    .X(_06824_));
 sky130_fd_sc_hd__a22o_1 _14620_ (.A1(net41),
    .A2(_06824_),
    .B1(_06768_),
    .B2(_06769_),
    .X(_06825_));
 sky130_fd_sc_hd__o21a_1 _14621_ (.A1(_06768_),
    .A2(_06769_),
    .B1(_06825_),
    .X(_06826_));
 sky130_fd_sc_hd__nand2_1 _14622_ (.A(net41),
    .B(_06268_),
    .Y(_06827_));
 sky130_fd_sc_hd__xnor2_1 _14623_ (.A(_06826_),
    .B(_06827_),
    .Y(_06828_));
 sky130_fd_sc_hd__xnor2_1 _14624_ (.A(_06823_),
    .B(_06828_),
    .Y(_06829_));
 sky130_fd_sc_hd__o21ba_1 _14625_ (.A1(_06766_),
    .A2(_06771_),
    .B1_N(_06764_),
    .X(_06830_));
 sky130_fd_sc_hd__a21o_1 _14626_ (.A1(_06766_),
    .A2(_06771_),
    .B1(_06830_),
    .X(_06831_));
 sky130_fd_sc_hd__buf_2 _14627_ (.A(_05605_),
    .X(_06832_));
 sky130_fd_sc_hd__nand2_2 _14628_ (.A(net25),
    .B(_06832_),
    .Y(_06833_));
 sky130_fd_sc_hd__o211a_1 _14629_ (.A1(_06106_),
    .A2(_05629_),
    .B1(_05640_),
    .C1(net20),
    .X(_06834_));
 sky130_fd_sc_hd__a211o_1 _14630_ (.A1(net20),
    .A2(_05640_),
    .B1(_05629_),
    .C1(_06106_),
    .X(_06835_));
 sky130_fd_sc_hd__or2b_1 _14631_ (.A(_06834_),
    .B_N(_06835_),
    .X(_06836_));
 sky130_fd_sc_hd__xnor2_2 _14632_ (.A(_06833_),
    .B(_06836_),
    .Y(_06837_));
 sky130_fd_sc_hd__o21a_1 _14633_ (.A1(_06760_),
    .A2(_06762_),
    .B1(_06761_),
    .X(_06838_));
 sky130_fd_sc_hd__a21o_1 _14634_ (.A1(_06760_),
    .A2(_06762_),
    .B1(_06838_),
    .X(_06839_));
 sky130_fd_sc_hd__nand2_1 _14635_ (.A(net40),
    .B(_06351_),
    .Y(_06840_));
 sky130_fd_sc_hd__nand2_1 _14636_ (.A(net34),
    .B(_05619_),
    .Y(_06841_));
 sky130_fd_sc_hd__nand2_1 _14637_ (.A(net36),
    .B(_05666_),
    .Y(_06842_));
 sky130_fd_sc_hd__xnor2_1 _14638_ (.A(_06841_),
    .B(_06842_),
    .Y(_06843_));
 sky130_fd_sc_hd__xnor2_2 _14639_ (.A(_06840_),
    .B(_06843_),
    .Y(_06844_));
 sky130_fd_sc_hd__xor2_1 _14640_ (.A(_06839_),
    .B(_06844_),
    .X(_06845_));
 sky130_fd_sc_hd__xnor2_2 _14641_ (.A(_06837_),
    .B(_06845_),
    .Y(_06846_));
 sky130_fd_sc_hd__xor2_1 _14642_ (.A(_06716_),
    .B(_06846_),
    .X(_06847_));
 sky130_fd_sc_hd__xnor2_1 _14643_ (.A(_06831_),
    .B(_06847_),
    .Y(_06848_));
 sky130_fd_sc_hd__nor2_1 _14644_ (.A(_06829_),
    .B(_06848_),
    .Y(_06849_));
 sky130_fd_sc_hd__nand2_1 _14645_ (.A(_06829_),
    .B(_06848_),
    .Y(_06850_));
 sky130_fd_sc_hd__and2b_1 _14646_ (.A_N(_06849_),
    .B(_06850_),
    .X(_06851_));
 sky130_fd_sc_hd__xor2_2 _14647_ (.A(_06820_),
    .B(_06851_),
    .X(_06852_));
 sky130_fd_sc_hd__a21o_1 _14648_ (.A1(_06758_),
    .A2(_06788_),
    .B1(_06785_),
    .X(_06853_));
 sky130_fd_sc_hd__o21ai_1 _14649_ (.A1(_06758_),
    .A2(_06788_),
    .B1(_06853_),
    .Y(_06854_));
 sky130_fd_sc_hd__a21o_1 _14650_ (.A1(_06755_),
    .A2(_06756_),
    .B1(_06753_),
    .X(_06855_));
 sky130_fd_sc_hd__o21a_1 _14651_ (.A1(_06755_),
    .A2(_06756_),
    .B1(_06855_),
    .X(_06856_));
 sky130_fd_sc_hd__xor2_1 _14652_ (.A(_06854_),
    .B(_06856_),
    .X(_06857_));
 sky130_fd_sc_hd__xnor2_2 _14653_ (.A(_06852_),
    .B(_06857_),
    .Y(_06858_));
 sky130_fd_sc_hd__xnor2_2 _14654_ (.A(_06819_),
    .B(_06858_),
    .Y(_06859_));
 sky130_fd_sc_hd__xnor2_4 _14655_ (.A(_06817_),
    .B(_06859_),
    .Y(_06860_));
 sky130_fd_sc_hd__a22o_1 _14656_ (.A1(net848),
    .A2(_06280_),
    .B1(_06860_),
    .B2(_06381_),
    .X(_00027_));
 sky130_fd_sc_hd__or2_1 _14657_ (.A(_06819_),
    .B(_06858_),
    .X(_06861_));
 sky130_fd_sc_hd__a221o_1 _14658_ (.A1(_06551_),
    .A2(_06807_),
    .B1(_06819_),
    .B2(_06858_),
    .C1(_06816_),
    .X(_06862_));
 sky130_fd_sc_hd__nand2_2 _14659_ (.A(_06861_),
    .B(_06862_),
    .Y(_06863_));
 sky130_fd_sc_hd__a21bo_1 _14660_ (.A1(_06852_),
    .A2(_06856_),
    .B1_N(_06854_),
    .X(_06864_));
 sky130_fd_sc_hd__o21ai_1 _14661_ (.A1(_06852_),
    .A2(_06856_),
    .B1(_06864_),
    .Y(_06865_));
 sky130_fd_sc_hd__o21ai_1 _14662_ (.A1(_06820_),
    .A2(_06849_),
    .B1(_06850_),
    .Y(_06866_));
 sky130_fd_sc_hd__buf_6 _14663_ (.A(_06268_),
    .X(_06867_));
 sky130_fd_sc_hd__or2_1 _14664_ (.A(_06823_),
    .B(_06826_),
    .X(_06868_));
 sky130_fd_sc_hd__and2_1 _14665_ (.A(_06823_),
    .B(_06826_),
    .X(_06869_));
 sky130_fd_sc_hd__a31o_1 _14666_ (.A1(\top0.periodTop_r[9] ),
    .A2(_06867_),
    .A3(_06868_),
    .B1(_06869_),
    .X(_06870_));
 sky130_fd_sc_hd__nand2_1 _14667_ (.A(_06831_),
    .B(_06846_),
    .Y(_06871_));
 sky130_fd_sc_hd__nor2_1 _14668_ (.A(_06831_),
    .B(_06846_),
    .Y(_06872_));
 sky130_fd_sc_hd__a21oi_2 _14669_ (.A1(_06716_),
    .A2(_06871_),
    .B1(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__nand2_1 _14670_ (.A(_06841_),
    .B(_06842_),
    .Y(_06874_));
 sky130_fd_sc_hd__nor2_1 _14671_ (.A(_06841_),
    .B(_06842_),
    .Y(_06875_));
 sky130_fd_sc_hd__a31o_1 _14672_ (.A1(net39),
    .A2(_06824_),
    .A3(_06874_),
    .B1(_06875_),
    .X(_06876_));
 sky130_fd_sc_hd__nand2_1 _14673_ (.A(net39),
    .B(_06268_),
    .Y(_06877_));
 sky130_fd_sc_hd__xor2_1 _14674_ (.A(_06876_),
    .B(_06877_),
    .X(_06878_));
 sky130_fd_sc_hd__xnor2_1 _14675_ (.A(_06873_),
    .B(_06878_),
    .Y(_06879_));
 sky130_fd_sc_hd__nand2_1 _14676_ (.A(_05626_),
    .B(_06832_),
    .Y(_06880_));
 sky130_fd_sc_hd__o32a_1 _14677_ (.A1(_05640_),
    .A2(_06212_),
    .A3(_06880_),
    .B1(_06832_),
    .B2(net25),
    .X(_06881_));
 sky130_fd_sc_hd__o22a_1 _14678_ (.A1(_06832_),
    .A2(_06212_),
    .B1(_06880_),
    .B2(net25),
    .X(_06882_));
 sky130_fd_sc_hd__o22a_1 _14679_ (.A1(_06217_),
    .A2(_05626_),
    .B1(_06882_),
    .B2(_06106_),
    .X(_06883_));
 sky130_fd_sc_hd__o21a_1 _14680_ (.A1(_06832_),
    .A2(_05640_),
    .B1(net20),
    .X(_06884_));
 sky130_fd_sc_hd__a21o_1 _14681_ (.A1(_05626_),
    .A2(_06760_),
    .B1(net20),
    .X(_06885_));
 sky130_fd_sc_hd__o221a_1 _14682_ (.A1(_05626_),
    .A2(_06832_),
    .B1(_06884_),
    .B2(net25),
    .C1(_06885_),
    .X(_06886_));
 sky130_fd_sc_hd__o221a_1 _14683_ (.A1(net31),
    .A2(_06881_),
    .B1(_06883_),
    .B2(_05731_),
    .C1(_06886_),
    .X(_06887_));
 sky130_fd_sc_hd__nand2_1 _14684_ (.A(net37),
    .B(_06351_),
    .Y(_06888_));
 sky130_fd_sc_hd__nand2_1 _14685_ (.A(net31),
    .B(_05619_),
    .Y(_06889_));
 sky130_fd_sc_hd__nand2_1 _14686_ (.A(net33),
    .B(_05666_),
    .Y(_06890_));
 sky130_fd_sc_hd__xnor2_1 _14687_ (.A(_06889_),
    .B(_06890_),
    .Y(_06891_));
 sky130_fd_sc_hd__xnor2_1 _14688_ (.A(_06888_),
    .B(_06891_),
    .Y(_06892_));
 sky130_fd_sc_hd__xor2_1 _14689_ (.A(_06887_),
    .B(_06892_),
    .X(_06893_));
 sky130_fd_sc_hd__o21ba_1 _14690_ (.A1(_06839_),
    .A2(_06844_),
    .B1_N(_06837_),
    .X(_06894_));
 sky130_fd_sc_hd__a21o_1 _14691_ (.A1(_06839_),
    .A2(_06844_),
    .B1(_06894_),
    .X(_06895_));
 sky130_fd_sc_hd__nor2_1 _14692_ (.A(_06893_),
    .B(_06895_),
    .Y(_06896_));
 sky130_fd_sc_hd__and2_1 _14693_ (.A(_06893_),
    .B(_06895_),
    .X(_06897_));
 sky130_fd_sc_hd__or2_1 _14694_ (.A(_06896_),
    .B(_06897_),
    .X(_06898_));
 sky130_fd_sc_hd__nand2_1 _14695_ (.A(_06879_),
    .B(_06898_),
    .Y(_06899_));
 sky130_fd_sc_hd__or2_1 _14696_ (.A(_06879_),
    .B(_06898_),
    .X(_06900_));
 sky130_fd_sc_hd__and2_1 _14697_ (.A(_06899_),
    .B(_06900_),
    .X(_06901_));
 sky130_fd_sc_hd__xnor2_1 _14698_ (.A(_06870_),
    .B(_06901_),
    .Y(_06902_));
 sky130_fd_sc_hd__xnor2_1 _14699_ (.A(_06866_),
    .B(_06902_),
    .Y(_06903_));
 sky130_fd_sc_hd__and2_1 _14700_ (.A(_06865_),
    .B(_06903_),
    .X(_06904_));
 sky130_fd_sc_hd__nor2_1 _14701_ (.A(_06865_),
    .B(_06903_),
    .Y(_06905_));
 sky130_fd_sc_hd__nor2_2 _14702_ (.A(_06904_),
    .B(_06905_),
    .Y(_06906_));
 sky130_fd_sc_hd__xnor2_4 _14703_ (.A(_06863_),
    .B(_06906_),
    .Y(_06907_));
 sky130_fd_sc_hd__a22o_1 _14704_ (.A1(net817),
    .A2(_06280_),
    .B1(_06907_),
    .B2(_05465_),
    .X(_00028_));
 sky130_fd_sc_hd__or2_1 _14705_ (.A(_06861_),
    .B(_06905_),
    .X(_06908_));
 sky130_fd_sc_hd__nand2_1 _14706_ (.A(_06865_),
    .B(_06903_),
    .Y(_06909_));
 sky130_fd_sc_hd__o211a_2 _14707_ (.A1(_06862_),
    .A2(_06905_),
    .B1(_06908_),
    .C1(_06909_),
    .X(_06910_));
 sky130_fd_sc_hd__inv_2 _14708_ (.A(_06876_),
    .Y(_06911_));
 sky130_fd_sc_hd__o21a_1 _14709_ (.A1(_06873_),
    .A2(_06911_),
    .B1(_06877_),
    .X(_06912_));
 sky130_fd_sc_hd__a21oi_2 _14710_ (.A1(_06873_),
    .A2(_06911_),
    .B1(_06912_),
    .Y(_06913_));
 sky130_fd_sc_hd__nand2_1 _14711_ (.A(_06889_),
    .B(_06890_),
    .Y(_06914_));
 sky130_fd_sc_hd__nor2_1 _14712_ (.A(_06889_),
    .B(_06890_),
    .Y(_06915_));
 sky130_fd_sc_hd__a31o_1 _14713_ (.A1(net36),
    .A2(_06824_),
    .A3(_06914_),
    .B1(_06915_),
    .X(_06916_));
 sky130_fd_sc_hd__nand2_1 _14714_ (.A(net37),
    .B(_06268_),
    .Y(_06917_));
 sky130_fd_sc_hd__xor2_1 _14715_ (.A(_06916_),
    .B(_06917_),
    .X(_06918_));
 sky130_fd_sc_hd__xnor2_1 _14716_ (.A(_06896_),
    .B(_06918_),
    .Y(_06919_));
 sky130_fd_sc_hd__nand2_1 _14717_ (.A(net34),
    .B(_06351_),
    .Y(_06920_));
 sky130_fd_sc_hd__nand2_1 _14718_ (.A(net25),
    .B(_05619_),
    .Y(_06921_));
 sky130_fd_sc_hd__nand2_1 _14719_ (.A(net31),
    .B(_05666_),
    .Y(_06922_));
 sky130_fd_sc_hd__xor2_1 _14720_ (.A(_06921_),
    .B(_06922_),
    .X(_06923_));
 sky130_fd_sc_hd__xnor2_2 _14721_ (.A(_06920_),
    .B(_06923_),
    .Y(_06924_));
 sky130_fd_sc_hd__and3_1 _14722_ (.A(net20),
    .B(_05626_),
    .C(_06833_),
    .X(_06925_));
 sky130_fd_sc_hd__xor2_2 _14723_ (.A(_06924_),
    .B(_06925_),
    .X(_06926_));
 sky130_fd_sc_hd__nor2_1 _14724_ (.A(_06832_),
    .B(_05731_),
    .Y(_06927_));
 sky130_fd_sc_hd__mux2_1 _14725_ (.A0(_06832_),
    .A1(_06927_),
    .S(net20),
    .X(_06928_));
 sky130_fd_sc_hd__a32o_1 _14726_ (.A1(_06832_),
    .A2(_05640_),
    .A3(_06323_),
    .B1(_06928_),
    .B2(net25),
    .X(_06929_));
 sky130_fd_sc_hd__and4_1 _14727_ (.A(_05629_),
    .B(_06832_),
    .C(_05640_),
    .D(_06320_),
    .X(_06930_));
 sky130_fd_sc_hd__and2b_1 _14728_ (.A_N(_06892_),
    .B(_06887_),
    .X(_06931_));
 sky130_fd_sc_hd__a311o_1 _14729_ (.A1(net31),
    .A2(_05626_),
    .A3(_06929_),
    .B1(_06930_),
    .C1(_06931_),
    .X(_06932_));
 sky130_fd_sc_hd__xor2_1 _14730_ (.A(_06926_),
    .B(_06932_),
    .X(_06933_));
 sky130_fd_sc_hd__and2_1 _14731_ (.A(_06919_),
    .B(_06933_),
    .X(_06934_));
 sky130_fd_sc_hd__buf_6 _14732_ (.A(_06934_),
    .X(_06935_));
 sky130_fd_sc_hd__nor2_1 _14733_ (.A(_06919_),
    .B(_06933_),
    .Y(_06936_));
 sky130_fd_sc_hd__nor2_1 _14734_ (.A(_06935_),
    .B(_06936_),
    .Y(_06937_));
 sky130_fd_sc_hd__xor2_1 _14735_ (.A(_06913_),
    .B(_06937_),
    .X(_06938_));
 sky130_fd_sc_hd__xnor2_1 _14736_ (.A(_06900_),
    .B(_06938_),
    .Y(_06939_));
 sky130_fd_sc_hd__o21ba_1 _14737_ (.A1(_06870_),
    .A2(_06901_),
    .B1_N(_06866_),
    .X(_06940_));
 sky130_fd_sc_hd__a21o_1 _14738_ (.A1(_06870_),
    .A2(_06901_),
    .B1(_06940_),
    .X(_06941_));
 sky130_fd_sc_hd__nor2_1 _14739_ (.A(_06939_),
    .B(_06941_),
    .Y(_06942_));
 sky130_fd_sc_hd__and2_1 _14740_ (.A(_06939_),
    .B(_06941_),
    .X(_06943_));
 sky130_fd_sc_hd__or2_1 _14741_ (.A(_06942_),
    .B(_06943_),
    .X(_06944_));
 sky130_fd_sc_hd__xnor2_2 _14742_ (.A(_06910_),
    .B(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__a22o_1 _14743_ (.A1(net807),
    .A2(_06279_),
    .B1(_06945_),
    .B2(_05465_),
    .X(_00029_));
 sky130_fd_sc_hd__nor2_1 _14744_ (.A(_06910_),
    .B(_06943_),
    .Y(_06946_));
 sky130_fd_sc_hd__nor2_1 _14745_ (.A(_06942_),
    .B(_06946_),
    .Y(_06947_));
 sky130_fd_sc_hd__a21bo_1 _14746_ (.A1(_06913_),
    .A2(_06937_),
    .B1_N(_06900_),
    .X(_06948_));
 sky130_fd_sc_hd__o21a_2 _14747_ (.A1(_06913_),
    .A2(_06937_),
    .B1(_06948_),
    .X(_06949_));
 sky130_fd_sc_hd__a21bo_1 _14748_ (.A1(_06896_),
    .A2(_06916_),
    .B1_N(_06917_),
    .X(_06950_));
 sky130_fd_sc_hd__o21ai_2 _14749_ (.A1(_06896_),
    .A2(_06916_),
    .B1(_06950_),
    .Y(_06951_));
 sky130_fd_sc_hd__nand2_2 _14750_ (.A(_06926_),
    .B(_06932_),
    .Y(_06952_));
 sky130_fd_sc_hd__nand2_1 _14751_ (.A(net31),
    .B(_06824_),
    .Y(_06953_));
 sky130_fd_sc_hd__and3_1 _14752_ (.A(net23),
    .B(_05723_),
    .C(_05724_),
    .X(_06954_));
 sky130_fd_sc_hd__and3_2 _14753_ (.A(net25),
    .B(_05726_),
    .C(_05727_),
    .X(_06955_));
 sky130_fd_sc_hd__xnor2_1 _14754_ (.A(_06954_),
    .B(_06955_),
    .Y(_06956_));
 sky130_fd_sc_hd__xnor2_2 _14755_ (.A(_06953_),
    .B(_06956_),
    .Y(_06957_));
 sky130_fd_sc_hd__and2b_1 _14756_ (.A_N(_06924_),
    .B(_06833_),
    .X(_06958_));
 sky130_fd_sc_hd__or3b_1 _14757_ (.A(_06958_),
    .B(_05629_),
    .C_N(net20),
    .X(_06959_));
 sky130_fd_sc_hd__xor2_2 _14758_ (.A(_06957_),
    .B(_06959_),
    .X(_06960_));
 sky130_fd_sc_hd__nand2_1 _14759_ (.A(_06921_),
    .B(_06922_),
    .Y(_06961_));
 sky130_fd_sc_hd__nor2_1 _14760_ (.A(_06921_),
    .B(_06922_),
    .Y(_06962_));
 sky130_fd_sc_hd__a31o_1 _14761_ (.A1(net33),
    .A2(_06824_),
    .A3(_06961_),
    .B1(_06962_),
    .X(_06963_));
 sky130_fd_sc_hd__nand2_1 _14762_ (.A(net34),
    .B(_06867_),
    .Y(_06964_));
 sky130_fd_sc_hd__xnor2_1 _14763_ (.A(_06963_),
    .B(_06964_),
    .Y(_06965_));
 sky130_fd_sc_hd__xnor2_1 _14764_ (.A(_06960_),
    .B(_06965_),
    .Y(_06966_));
 sky130_fd_sc_hd__xnor2_2 _14765_ (.A(_06952_),
    .B(_06966_),
    .Y(_06967_));
 sky130_fd_sc_hd__xnor2_1 _14766_ (.A(_06951_),
    .B(_06967_),
    .Y(_06968_));
 sky130_fd_sc_hd__xnor2_1 _14767_ (.A(_06935_),
    .B(_06968_),
    .Y(_06969_));
 sky130_fd_sc_hd__xnor2_2 _14768_ (.A(_06949_),
    .B(_06969_),
    .Y(_06970_));
 sky130_fd_sc_hd__xnor2_2 _14769_ (.A(_06947_),
    .B(_06970_),
    .Y(_06971_));
 sky130_fd_sc_hd__a22o_1 _14770_ (.A1(net857),
    .A2(_06279_),
    .B1(_06971_),
    .B2(_05465_),
    .X(_00030_));
 sky130_fd_sc_hd__or2_1 _14771_ (.A(_06957_),
    .B(_06959_),
    .X(_06972_));
 sky130_fd_sc_hd__a22o_1 _14772_ (.A1(net31),
    .A2(_06824_),
    .B1(_06954_),
    .B2(_06955_),
    .X(_06973_));
 sky130_fd_sc_hd__o21a_1 _14773_ (.A1(_06954_),
    .A2(_06955_),
    .B1(_06973_),
    .X(_06974_));
 sky130_fd_sc_hd__nand2_1 _14774_ (.A(net26),
    .B(_06824_),
    .Y(_06975_));
 sky130_fd_sc_hd__nand2_1 _14775_ (.A(net21),
    .B(_05666_),
    .Y(_06976_));
 sky130_fd_sc_hd__xor2_2 _14776_ (.A(_06975_),
    .B(_06976_),
    .X(_06977_));
 sky130_fd_sc_hd__nand2_1 _14777_ (.A(net31),
    .B(_06867_),
    .Y(_06978_));
 sky130_fd_sc_hd__xor2_1 _14778_ (.A(_06977_),
    .B(_06978_),
    .X(_06979_));
 sky130_fd_sc_hd__xnor2_1 _14779_ (.A(_06974_),
    .B(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__xnor2_1 _14780_ (.A(_06972_),
    .B(_06980_),
    .Y(_06981_));
 sky130_fd_sc_hd__inv_2 _14781_ (.A(_06981_),
    .Y(_06982_));
 sky130_fd_sc_hd__nor2_1 _14782_ (.A(_06960_),
    .B(_06963_),
    .Y(_06983_));
 sky130_fd_sc_hd__and2_1 _14783_ (.A(_06960_),
    .B(_06963_),
    .X(_06984_));
 sky130_fd_sc_hd__o21ba_1 _14784_ (.A1(_06952_),
    .A2(_06983_),
    .B1_N(_06984_),
    .X(_06985_));
 sky130_fd_sc_hd__and3_1 _14785_ (.A(net34),
    .B(_06867_),
    .C(_06984_),
    .X(_06986_));
 sky130_fd_sc_hd__mux2_1 _14786_ (.A0(_06986_),
    .A1(_06983_),
    .S(_06952_),
    .X(_06987_));
 sky130_fd_sc_hd__a21oi_2 _14787_ (.A1(_06964_),
    .A2(_06985_),
    .B1(_06987_),
    .Y(_06988_));
 sky130_fd_sc_hd__xnor2_4 _14788_ (.A(_06982_),
    .B(_06988_),
    .Y(_06989_));
 sky130_fd_sc_hd__nand2_1 _14789_ (.A(_06951_),
    .B(_06967_),
    .Y(_06990_));
 sky130_fd_sc_hd__or2_1 _14790_ (.A(_06949_),
    .B(_06990_),
    .X(_06991_));
 sky130_fd_sc_hd__clkinvlp_2 _14791_ (.A(_06942_),
    .Y(_06992_));
 sky130_fd_sc_hd__nor2_1 _14792_ (.A(_06951_),
    .B(_06967_),
    .Y(_06993_));
 sky130_fd_sc_hd__o21a_1 _14793_ (.A1(_06949_),
    .A2(_06993_),
    .B1(_06990_),
    .X(_06994_));
 sky130_fd_sc_hd__or2_1 _14794_ (.A(_06943_),
    .B(_06994_),
    .X(_06995_));
 sky130_fd_sc_hd__o221a_1 _14795_ (.A1(_06992_),
    .A2(_06994_),
    .B1(_06995_),
    .B2(_06910_),
    .C1(_06991_),
    .X(_06996_));
 sky130_fd_sc_hd__a22o_1 _14796_ (.A1(_06949_),
    .A2(_06993_),
    .B1(_06994_),
    .B2(_06935_),
    .X(_06997_));
 sky130_fd_sc_hd__or3b_1 _14797_ (.A(_06942_),
    .B(_06946_),
    .C_N(_06997_),
    .X(_06998_));
 sky130_fd_sc_hd__o221a_1 _14798_ (.A1(_06947_),
    .A2(_06991_),
    .B1(_06996_),
    .B2(_06935_),
    .C1(_06998_),
    .X(_06999_));
 sky130_fd_sc_hd__xor2_2 _14799_ (.A(_06989_),
    .B(_06999_),
    .X(_07000_));
 sky130_fd_sc_hd__a22o_1 _14800_ (.A1(net868),
    .A2(_06279_),
    .B1(_07000_),
    .B2(_05465_),
    .X(_00031_));
 sky130_fd_sc_hd__and2_1 _14801_ (.A(_06989_),
    .B(_06990_),
    .X(_07001_));
 sky130_fd_sc_hd__o22a_1 _14802_ (.A1(_06989_),
    .A2(_06993_),
    .B1(_07001_),
    .B2(_06949_),
    .X(_07002_));
 sky130_fd_sc_hd__o22a_1 _14803_ (.A1(_06989_),
    .A2(_06994_),
    .B1(_07002_),
    .B2(_06935_),
    .X(_07003_));
 sky130_fd_sc_hd__or2_1 _14804_ (.A(_06943_),
    .B(_06949_),
    .X(_07004_));
 sky130_fd_sc_hd__o21a_1 _14805_ (.A1(_06935_),
    .A2(_07004_),
    .B1(_06989_),
    .X(_07005_));
 sky130_fd_sc_hd__a21o_1 _14806_ (.A1(_06935_),
    .A2(_07004_),
    .B1(_07001_),
    .X(_07006_));
 sky130_fd_sc_hd__o221a_1 _14807_ (.A1(_06989_),
    .A2(_06990_),
    .B1(_07005_),
    .B2(_06993_),
    .C1(_07006_),
    .X(_07007_));
 sky130_fd_sc_hd__a31o_1 _14808_ (.A1(_06910_),
    .A2(_06992_),
    .A3(_07003_),
    .B1(_07007_),
    .X(_07008_));
 sky130_fd_sc_hd__inv_2 _14809_ (.A(_06972_),
    .Y(_07009_));
 sky130_fd_sc_hd__or2_1 _14810_ (.A(_06974_),
    .B(_06977_),
    .X(_07010_));
 sky130_fd_sc_hd__a21o_1 _14811_ (.A1(_06974_),
    .A2(_06977_),
    .B1(_07009_),
    .X(_07011_));
 sky130_fd_sc_hd__a21bo_1 _14812_ (.A1(_07010_),
    .A2(_07011_),
    .B1_N(_06978_),
    .X(_07012_));
 sky130_fd_sc_hd__o21a_1 _14813_ (.A1(_07009_),
    .A2(_07010_),
    .B1(_07012_),
    .X(_07013_));
 sky130_fd_sc_hd__and2_1 _14814_ (.A(net21),
    .B(_06824_),
    .X(_07014_));
 sky130_fd_sc_hd__o21ai_1 _14815_ (.A1(_05666_),
    .A2(_06867_),
    .B1(net26),
    .Y(_07015_));
 sky130_fd_sc_hd__nand2_1 _14816_ (.A(net21),
    .B(_06824_),
    .Y(_07016_));
 sky130_fd_sc_hd__o211a_1 _14817_ (.A1(_05666_),
    .A2(_07016_),
    .B1(_06867_),
    .C1(net26),
    .X(_07017_));
 sky130_fd_sc_hd__a21oi_1 _14818_ (.A1(_07014_),
    .A2(_07015_),
    .B1(_07017_),
    .Y(_07018_));
 sky130_fd_sc_hd__or2b_1 _14819_ (.A(_07013_),
    .B_N(_07018_),
    .X(_07019_));
 sky130_fd_sc_hd__or2b_1 _14820_ (.A(_07018_),
    .B_N(_07013_),
    .X(_07020_));
 sky130_fd_sc_hd__nand2_1 _14821_ (.A(_07019_),
    .B(_07020_),
    .Y(_07021_));
 sky130_fd_sc_hd__nor2_1 _14822_ (.A(_06981_),
    .B(_06984_),
    .Y(_07022_));
 sky130_fd_sc_hd__o22a_1 _14823_ (.A1(_06982_),
    .A2(_06983_),
    .B1(_07022_),
    .B2(_06952_),
    .X(_07023_));
 sky130_fd_sc_hd__o22a_1 _14824_ (.A1(_06982_),
    .A2(_06985_),
    .B1(_07023_),
    .B2(_06964_),
    .X(_07024_));
 sky130_fd_sc_hd__nor2_1 _14825_ (.A(_07021_),
    .B(_07024_),
    .Y(_07025_));
 sky130_fd_sc_hd__nand2_1 _14826_ (.A(_07021_),
    .B(_07024_),
    .Y(_07026_));
 sky130_fd_sc_hd__or2b_1 _14827_ (.A(_07025_),
    .B_N(_07026_),
    .X(_07027_));
 sky130_fd_sc_hd__xnor2_2 _14828_ (.A(_07008_),
    .B(_07027_),
    .Y(_07028_));
 sky130_fd_sc_hd__a22o_1 _14829_ (.A1(net851),
    .A2(_06279_),
    .B1(_07028_),
    .B2(_05465_),
    .X(_00032_));
 sky130_fd_sc_hd__and3b_1 _14830_ (.A_N(_06867_),
    .B(_05726_),
    .C(_05727_),
    .X(_07029_));
 sky130_fd_sc_hd__mux2_1 _14831_ (.A0(_07029_),
    .A1(_06867_),
    .S(_06975_),
    .X(_07030_));
 sky130_fd_sc_hd__nand2_1 _14832_ (.A(net21),
    .B(_07030_),
    .Y(_07031_));
 sky130_fd_sc_hd__xnor2_1 _14833_ (.A(_07020_),
    .B(_07031_),
    .Y(_07032_));
 sky130_fd_sc_hd__o21a_1 _14834_ (.A1(_07008_),
    .A2(_07025_),
    .B1(_07026_),
    .X(_07033_));
 sky130_fd_sc_hd__xnor2_1 _14835_ (.A(_07032_),
    .B(_07033_),
    .Y(_07034_));
 sky130_fd_sc_hd__a22o_1 _14836_ (.A1(net824),
    .A2(_06279_),
    .B1(_07034_),
    .B2(_05465_),
    .X(_00033_));
 sky130_fd_sc_hd__and3b_1 _14837_ (.A_N(_06955_),
    .B(_07013_),
    .C(_07014_),
    .X(_07035_));
 sky130_fd_sc_hd__o211a_1 _14838_ (.A1(_07013_),
    .A2(_07014_),
    .B1(net26),
    .C1(_06867_),
    .X(_07036_));
 sky130_fd_sc_hd__a21o_1 _14839_ (.A1(_06824_),
    .A2(_06955_),
    .B1(_06867_),
    .X(_07037_));
 sky130_fd_sc_hd__o311a_1 _14840_ (.A1(_07033_),
    .A2(_07035_),
    .A3(_07036_),
    .B1(_07037_),
    .C1(net20),
    .X(_07038_));
 sky130_fd_sc_hd__a22o_1 _14841_ (.A1(net858),
    .A2(_06279_),
    .B1(_07038_),
    .B2(_05465_),
    .X(_00034_));
 sky130_fd_sc_hd__a21oi_1 _14842_ (.A1(\state[0] ),
    .A2(_05425_),
    .B1(_05422_),
    .Y(_07039_));
 sky130_fd_sc_hd__a21boi_1 _14843_ (.A1(\state[0] ),
    .A2(_05426_),
    .B1_N(net7),
    .Y(_07040_));
 sky130_fd_sc_hd__o22a_1 _14844_ (.A1(net7),
    .A2(_07039_),
    .B1(_07040_),
    .B2(net744),
    .X(_00035_));
 sky130_fd_sc_hd__nand2_4 _14845_ (.A(\state[0] ),
    .B(net17),
    .Y(_07041_));
 sky130_fd_sc_hd__buf_4 _14846_ (.A(_07041_),
    .X(_07042_));
 sky130_fd_sc_hd__mux2_1 _14847_ (.A0(\spi0.data_packed[64] ),
    .A1(\top0.kpd[0] ),
    .S(_07042_),
    .X(_07043_));
 sky130_fd_sc_hd__clkbuf_1 _14848_ (.A(_07043_),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _14849_ (.A0(\spi0.data_packed[65] ),
    .A1(\top0.kpd[1] ),
    .S(_07042_),
    .X(_07044_));
 sky130_fd_sc_hd__clkbuf_1 _14850_ (.A(_07044_),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_1 _14851_ (.A0(\spi0.data_packed[66] ),
    .A1(\top0.kpd[2] ),
    .S(_07042_),
    .X(_07045_));
 sky130_fd_sc_hd__clkbuf_1 _14852_ (.A(_07045_),
    .X(_00038_));
 sky130_fd_sc_hd__mux2_1 _14853_ (.A0(\spi0.data_packed[67] ),
    .A1(\top0.kpd[3] ),
    .S(_07042_),
    .X(_07046_));
 sky130_fd_sc_hd__clkbuf_1 _14854_ (.A(_07046_),
    .X(_00039_));
 sky130_fd_sc_hd__mux2_1 _14855_ (.A0(\spi0.data_packed[68] ),
    .A1(\top0.kpd[4] ),
    .S(_07042_),
    .X(_07047_));
 sky130_fd_sc_hd__clkbuf_1 _14856_ (.A(_07047_),
    .X(_00040_));
 sky130_fd_sc_hd__mux2_1 _14857_ (.A0(\spi0.data_packed[69] ),
    .A1(\top0.kpd[5] ),
    .S(_07042_),
    .X(_07048_));
 sky130_fd_sc_hd__clkbuf_1 _14858_ (.A(_07048_),
    .X(_00041_));
 sky130_fd_sc_hd__mux2_1 _14859_ (.A0(\spi0.data_packed[70] ),
    .A1(\top0.kpd[6] ),
    .S(_07042_),
    .X(_07049_));
 sky130_fd_sc_hd__clkbuf_1 _14860_ (.A(_07049_),
    .X(_00042_));
 sky130_fd_sc_hd__mux2_1 _14861_ (.A0(\spi0.data_packed[71] ),
    .A1(\top0.kpd[7] ),
    .S(_07042_),
    .X(_07050_));
 sky130_fd_sc_hd__clkbuf_1 _14862_ (.A(_07050_),
    .X(_00043_));
 sky130_fd_sc_hd__mux2_1 _14863_ (.A0(\spi0.data_packed[72] ),
    .A1(\top0.kpd[8] ),
    .S(_07042_),
    .X(_07051_));
 sky130_fd_sc_hd__clkbuf_1 _14864_ (.A(_07051_),
    .X(_00044_));
 sky130_fd_sc_hd__mux2_1 _14865_ (.A0(\spi0.data_packed[73] ),
    .A1(\top0.kpd[9] ),
    .S(_07042_),
    .X(_07052_));
 sky130_fd_sc_hd__clkbuf_1 _14866_ (.A(_07052_),
    .X(_00045_));
 sky130_fd_sc_hd__buf_4 _14867_ (.A(_07041_),
    .X(_07053_));
 sky130_fd_sc_hd__mux2_1 _14868_ (.A0(\spi0.data_packed[74] ),
    .A1(\top0.kpd[10] ),
    .S(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__clkbuf_1 _14869_ (.A(_07054_),
    .X(_00046_));
 sky130_fd_sc_hd__mux2_1 _14870_ (.A0(\spi0.data_packed[75] ),
    .A1(\top0.kpd[11] ),
    .S(_07053_),
    .X(_07055_));
 sky130_fd_sc_hd__clkbuf_1 _14871_ (.A(_07055_),
    .X(_00047_));
 sky130_fd_sc_hd__mux2_1 _14872_ (.A0(\spi0.data_packed[76] ),
    .A1(\top0.kpd[12] ),
    .S(_07053_),
    .X(_07056_));
 sky130_fd_sc_hd__clkbuf_1 _14873_ (.A(_07056_),
    .X(_00048_));
 sky130_fd_sc_hd__mux2_1 _14874_ (.A0(\spi0.data_packed[77] ),
    .A1(\top0.kpd[13] ),
    .S(_07053_),
    .X(_07057_));
 sky130_fd_sc_hd__clkbuf_1 _14875_ (.A(_07057_),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_1 _14876_ (.A0(\spi0.data_packed[78] ),
    .A1(\top0.kpd[14] ),
    .S(_07053_),
    .X(_07058_));
 sky130_fd_sc_hd__clkbuf_1 _14877_ (.A(_07058_),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _14878_ (.A0(\spi0.data_packed[79] ),
    .A1(\top0.kpd[15] ),
    .S(_07053_),
    .X(_07059_));
 sky130_fd_sc_hd__clkbuf_1 _14879_ (.A(_07059_),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _14880_ (.A0(\spi0.data_packed[48] ),
    .A1(\top0.kpq[0] ),
    .S(_07053_),
    .X(_07060_));
 sky130_fd_sc_hd__clkbuf_1 _14881_ (.A(_07060_),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _14882_ (.A0(\spi0.data_packed[49] ),
    .A1(\top0.kpq[1] ),
    .S(_07053_),
    .X(_07061_));
 sky130_fd_sc_hd__clkbuf_1 _14883_ (.A(_07061_),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _14884_ (.A0(\spi0.data_packed[50] ),
    .A1(\top0.kpq[2] ),
    .S(_07053_),
    .X(_07062_));
 sky130_fd_sc_hd__clkbuf_1 _14885_ (.A(_07062_),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _14886_ (.A0(\spi0.data_packed[51] ),
    .A1(\top0.kpq[3] ),
    .S(_07053_),
    .X(_07063_));
 sky130_fd_sc_hd__clkbuf_1 _14887_ (.A(_07063_),
    .X(_00055_));
 sky130_fd_sc_hd__clkbuf_4 _14888_ (.A(_07041_),
    .X(_07064_));
 sky130_fd_sc_hd__mux2_1 _14889_ (.A0(\spi0.data_packed[52] ),
    .A1(\top0.kpq[4] ),
    .S(_07064_),
    .X(_07065_));
 sky130_fd_sc_hd__clkbuf_1 _14890_ (.A(_07065_),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _14891_ (.A0(\spi0.data_packed[53] ),
    .A1(\top0.kpq[5] ),
    .S(_07064_),
    .X(_07066_));
 sky130_fd_sc_hd__clkbuf_1 _14892_ (.A(_07066_),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _14893_ (.A0(\spi0.data_packed[54] ),
    .A1(\top0.kpq[6] ),
    .S(_07064_),
    .X(_07067_));
 sky130_fd_sc_hd__clkbuf_1 _14894_ (.A(_07067_),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _14895_ (.A0(\spi0.data_packed[55] ),
    .A1(\top0.kpq[7] ),
    .S(_07064_),
    .X(_07068_));
 sky130_fd_sc_hd__clkbuf_1 _14896_ (.A(_07068_),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _14897_ (.A0(\spi0.data_packed[56] ),
    .A1(\top0.kpq[8] ),
    .S(_07064_),
    .X(_07069_));
 sky130_fd_sc_hd__clkbuf_1 _14898_ (.A(_07069_),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _14899_ (.A0(\spi0.data_packed[57] ),
    .A1(\top0.kpq[9] ),
    .S(_07064_),
    .X(_07070_));
 sky130_fd_sc_hd__clkbuf_1 _14900_ (.A(_07070_),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _14901_ (.A0(\spi0.data_packed[58] ),
    .A1(\top0.kpq[10] ),
    .S(_07064_),
    .X(_07071_));
 sky130_fd_sc_hd__clkbuf_1 _14902_ (.A(_07071_),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _14903_ (.A0(\spi0.data_packed[59] ),
    .A1(\top0.kpq[11] ),
    .S(_07064_),
    .X(_07072_));
 sky130_fd_sc_hd__clkbuf_1 _14904_ (.A(_07072_),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _14905_ (.A0(\spi0.data_packed[60] ),
    .A1(\top0.kpq[12] ),
    .S(_07064_),
    .X(_07073_));
 sky130_fd_sc_hd__clkbuf_1 _14906_ (.A(_07073_),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _14907_ (.A0(\spi0.data_packed[61] ),
    .A1(\top0.kpq[13] ),
    .S(_07064_),
    .X(_07074_));
 sky130_fd_sc_hd__clkbuf_1 _14908_ (.A(_07074_),
    .X(_00065_));
 sky130_fd_sc_hd__buf_4 _14909_ (.A(_07041_),
    .X(_07075_));
 sky130_fd_sc_hd__mux2_1 _14910_ (.A0(\spi0.data_packed[62] ),
    .A1(\top0.kpq[14] ),
    .S(_07075_),
    .X(_07076_));
 sky130_fd_sc_hd__clkbuf_1 _14911_ (.A(_07076_),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _14912_ (.A0(\spi0.data_packed[63] ),
    .A1(\top0.kpq[15] ),
    .S(_07075_),
    .X(_07077_));
 sky130_fd_sc_hd__clkbuf_1 _14913_ (.A(_07077_),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_1 _14914_ (.A0(\spi0.data_packed[32] ),
    .A1(\top0.kid[0] ),
    .S(_07075_),
    .X(_07078_));
 sky130_fd_sc_hd__clkbuf_1 _14915_ (.A(_07078_),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_1 _14916_ (.A0(\spi0.data_packed[33] ),
    .A1(\top0.kid[1] ),
    .S(_07075_),
    .X(_07079_));
 sky130_fd_sc_hd__clkbuf_1 _14917_ (.A(_07079_),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _14918_ (.A0(\spi0.data_packed[34] ),
    .A1(\top0.kid[2] ),
    .S(_07075_),
    .X(_07080_));
 sky130_fd_sc_hd__clkbuf_1 _14919_ (.A(_07080_),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _14920_ (.A0(\spi0.data_packed[35] ),
    .A1(\top0.kid[3] ),
    .S(_07075_),
    .X(_07081_));
 sky130_fd_sc_hd__clkbuf_1 _14921_ (.A(_07081_),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _14922_ (.A0(\spi0.data_packed[36] ),
    .A1(\top0.kid[4] ),
    .S(_07075_),
    .X(_07082_));
 sky130_fd_sc_hd__clkbuf_1 _14923_ (.A(_07082_),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _14924_ (.A0(\spi0.data_packed[37] ),
    .A1(\top0.kid[5] ),
    .S(_07075_),
    .X(_07083_));
 sky130_fd_sc_hd__clkbuf_1 _14925_ (.A(_07083_),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _14926_ (.A0(\spi0.data_packed[38] ),
    .A1(\top0.kid[6] ),
    .S(_07075_),
    .X(_07084_));
 sky130_fd_sc_hd__clkbuf_1 _14927_ (.A(_07084_),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _14928_ (.A0(\spi0.data_packed[39] ),
    .A1(\top0.kid[7] ),
    .S(_07075_),
    .X(_07085_));
 sky130_fd_sc_hd__clkbuf_1 _14929_ (.A(_07085_),
    .X(_00075_));
 sky130_fd_sc_hd__buf_4 _14930_ (.A(_07041_),
    .X(_07086_));
 sky130_fd_sc_hd__mux2_1 _14931_ (.A0(\spi0.data_packed[40] ),
    .A1(\top0.kid[8] ),
    .S(_07086_),
    .X(_07087_));
 sky130_fd_sc_hd__clkbuf_1 _14932_ (.A(_07087_),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _14933_ (.A0(\spi0.data_packed[41] ),
    .A1(\top0.kid[9] ),
    .S(_07086_),
    .X(_07088_));
 sky130_fd_sc_hd__clkbuf_1 _14934_ (.A(_07088_),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _14935_ (.A0(\spi0.data_packed[42] ),
    .A1(\top0.kid[10] ),
    .S(_07086_),
    .X(_07089_));
 sky130_fd_sc_hd__clkbuf_1 _14936_ (.A(_07089_),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _14937_ (.A0(\spi0.data_packed[43] ),
    .A1(\top0.kid[11] ),
    .S(_07086_),
    .X(_07090_));
 sky130_fd_sc_hd__clkbuf_1 _14938_ (.A(_07090_),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _14939_ (.A0(\spi0.data_packed[44] ),
    .A1(\top0.kid[12] ),
    .S(_07086_),
    .X(_07091_));
 sky130_fd_sc_hd__clkbuf_1 _14940_ (.A(_07091_),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _14941_ (.A0(\spi0.data_packed[45] ),
    .A1(\top0.kid[13] ),
    .S(_07086_),
    .X(_07092_));
 sky130_fd_sc_hd__clkbuf_1 _14942_ (.A(_07092_),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _14943_ (.A0(\spi0.data_packed[46] ),
    .A1(\top0.kid[14] ),
    .S(_07086_),
    .X(_07093_));
 sky130_fd_sc_hd__clkbuf_1 _14944_ (.A(_07093_),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _14945_ (.A0(\spi0.data_packed[47] ),
    .A1(\top0.kid[15] ),
    .S(_07086_),
    .X(_07094_));
 sky130_fd_sc_hd__clkbuf_1 _14946_ (.A(_07094_),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _14947_ (.A0(\spi0.data_packed[16] ),
    .A1(\top0.kiq[0] ),
    .S(_07086_),
    .X(_07095_));
 sky130_fd_sc_hd__clkbuf_1 _14948_ (.A(_07095_),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _14949_ (.A0(\spi0.data_packed[17] ),
    .A1(\top0.kiq[1] ),
    .S(_07086_),
    .X(_07096_));
 sky130_fd_sc_hd__clkbuf_1 _14950_ (.A(_07096_),
    .X(_00085_));
 sky130_fd_sc_hd__buf_4 _14951_ (.A(_07041_),
    .X(_07097_));
 sky130_fd_sc_hd__mux2_1 _14952_ (.A0(\spi0.data_packed[18] ),
    .A1(\top0.kiq[2] ),
    .S(_07097_),
    .X(_07098_));
 sky130_fd_sc_hd__clkbuf_1 _14953_ (.A(_07098_),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_1 _14954_ (.A0(\spi0.data_packed[19] ),
    .A1(\top0.kiq[3] ),
    .S(_07097_),
    .X(_07099_));
 sky130_fd_sc_hd__clkbuf_1 _14955_ (.A(_07099_),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _14956_ (.A0(\spi0.data_packed[20] ),
    .A1(\top0.kiq[4] ),
    .S(_07097_),
    .X(_07100_));
 sky130_fd_sc_hd__clkbuf_1 _14957_ (.A(_07100_),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _14958_ (.A0(\spi0.data_packed[21] ),
    .A1(\top0.kiq[5] ),
    .S(_07097_),
    .X(_07101_));
 sky130_fd_sc_hd__clkbuf_1 _14959_ (.A(_07101_),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _14960_ (.A0(\spi0.data_packed[22] ),
    .A1(\top0.kiq[6] ),
    .S(_07097_),
    .X(_07102_));
 sky130_fd_sc_hd__clkbuf_1 _14961_ (.A(_07102_),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _14962_ (.A0(\spi0.data_packed[23] ),
    .A1(\top0.kiq[7] ),
    .S(_07097_),
    .X(_07103_));
 sky130_fd_sc_hd__clkbuf_1 _14963_ (.A(_07103_),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _14964_ (.A0(\spi0.data_packed[24] ),
    .A1(\top0.kiq[8] ),
    .S(_07097_),
    .X(_07104_));
 sky130_fd_sc_hd__clkbuf_1 _14965_ (.A(_07104_),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _14966_ (.A0(\spi0.data_packed[25] ),
    .A1(\top0.kiq[9] ),
    .S(_07097_),
    .X(_07105_));
 sky130_fd_sc_hd__clkbuf_1 _14967_ (.A(_07105_),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _14968_ (.A0(\spi0.data_packed[26] ),
    .A1(\top0.kiq[10] ),
    .S(_07097_),
    .X(_07106_));
 sky130_fd_sc_hd__clkbuf_1 _14969_ (.A(_07106_),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _14970_ (.A0(\spi0.data_packed[27] ),
    .A1(\top0.kiq[11] ),
    .S(_07097_),
    .X(_07107_));
 sky130_fd_sc_hd__clkbuf_1 _14971_ (.A(_07107_),
    .X(_00095_));
 sky130_fd_sc_hd__clkbuf_4 _14972_ (.A(_07041_),
    .X(_07108_));
 sky130_fd_sc_hd__mux2_1 _14973_ (.A0(\spi0.data_packed[28] ),
    .A1(\top0.kiq[12] ),
    .S(_07108_),
    .X(_07109_));
 sky130_fd_sc_hd__clkbuf_1 _14974_ (.A(_07109_),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _14975_ (.A0(\spi0.data_packed[29] ),
    .A1(\top0.kiq[13] ),
    .S(_07108_),
    .X(_07110_));
 sky130_fd_sc_hd__clkbuf_1 _14976_ (.A(_07110_),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _14977_ (.A0(\spi0.data_packed[30] ),
    .A1(\top0.kiq[14] ),
    .S(_07108_),
    .X(_07111_));
 sky130_fd_sc_hd__clkbuf_1 _14978_ (.A(_07111_),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _14979_ (.A0(\spi0.data_packed[31] ),
    .A1(\top0.kiq[15] ),
    .S(_07108_),
    .X(_07112_));
 sky130_fd_sc_hd__clkbuf_1 _14980_ (.A(_07112_),
    .X(_00099_));
 sky130_fd_sc_hd__nor2_1 _14981_ (.A(\top0.svm0.state[1] ),
    .B(\top0.svm0.state[0] ),
    .Y(_07113_));
 sky130_fd_sc_hd__and2_1 _14982_ (.A(\top0.start_svm ),
    .B(_07113_),
    .X(_07114_));
 sky130_fd_sc_hd__inv_2 _14983_ (.A(net171),
    .Y(_07115_));
 sky130_fd_sc_hd__mux2_1 _14984_ (.A0(_06276_),
    .A1(_07114_),
    .S(_07115_),
    .X(_07116_));
 sky130_fd_sc_hd__buf_2 _14985_ (.A(_07116_),
    .X(_07117_));
 sky130_fd_sc_hd__or2_1 _14986_ (.A(\top0.svm0.delta[0] ),
    .B(_07117_),
    .X(_07118_));
 sky130_fd_sc_hd__clkbuf_1 _14987_ (.A(_07118_),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _14988_ (.A0(\spi0.data_packed[0] ),
    .A1(\top0.periodTop[0] ),
    .S(_07108_),
    .X(_07119_));
 sky130_fd_sc_hd__clkbuf_1 _14989_ (.A(_07119_),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _14990_ (.A0(\spi0.data_packed[1] ),
    .A1(\top0.periodTop[1] ),
    .S(_07108_),
    .X(_07120_));
 sky130_fd_sc_hd__clkbuf_1 _14991_ (.A(_07120_),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _14992_ (.A0(\spi0.data_packed[2] ),
    .A1(\top0.periodTop[2] ),
    .S(_07108_),
    .X(_07121_));
 sky130_fd_sc_hd__clkbuf_1 _14993_ (.A(_07121_),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _14994_ (.A0(\spi0.data_packed[3] ),
    .A1(\top0.periodTop[3] ),
    .S(_07108_),
    .X(_07122_));
 sky130_fd_sc_hd__clkbuf_1 _14995_ (.A(_07122_),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _14996_ (.A0(\spi0.data_packed[4] ),
    .A1(\top0.periodTop[4] ),
    .S(_07108_),
    .X(_07123_));
 sky130_fd_sc_hd__clkbuf_1 _14997_ (.A(_07123_),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _14998_ (.A0(\spi0.data_packed[5] ),
    .A1(\top0.periodTop[5] ),
    .S(_07108_),
    .X(_07124_));
 sky130_fd_sc_hd__clkbuf_1 _14999_ (.A(_07124_),
    .X(_00106_));
 sky130_fd_sc_hd__clkbuf_4 _15000_ (.A(_07041_),
    .X(_07125_));
 sky130_fd_sc_hd__mux2_1 _15001_ (.A0(\spi0.data_packed[6] ),
    .A1(\top0.periodTop[6] ),
    .S(_07125_),
    .X(_07126_));
 sky130_fd_sc_hd__clkbuf_1 _15002_ (.A(_07126_),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _15003_ (.A0(\spi0.data_packed[7] ),
    .A1(\top0.periodTop[7] ),
    .S(_07125_),
    .X(_07127_));
 sky130_fd_sc_hd__clkbuf_1 _15004_ (.A(_07127_),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _15005_ (.A0(\spi0.data_packed[8] ),
    .A1(\top0.periodTop[8] ),
    .S(_07125_),
    .X(_07128_));
 sky130_fd_sc_hd__clkbuf_1 _15006_ (.A(_07128_),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _15007_ (.A0(\spi0.data_packed[9] ),
    .A1(\top0.periodTop[9] ),
    .S(_07125_),
    .X(_07129_));
 sky130_fd_sc_hd__clkbuf_1 _15008_ (.A(_07129_),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _15009_ (.A0(\spi0.data_packed[10] ),
    .A1(\top0.periodTop[10] ),
    .S(_07125_),
    .X(_07130_));
 sky130_fd_sc_hd__clkbuf_1 _15010_ (.A(_07130_),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _15011_ (.A0(\spi0.data_packed[11] ),
    .A1(\top0.periodTop[11] ),
    .S(_07125_),
    .X(_07131_));
 sky130_fd_sc_hd__clkbuf_1 _15012_ (.A(_07131_),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _15013_ (.A0(\spi0.data_packed[12] ),
    .A1(\top0.periodTop[12] ),
    .S(_07125_),
    .X(_07132_));
 sky130_fd_sc_hd__clkbuf_1 _15014_ (.A(_07132_),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _15015_ (.A0(\spi0.data_packed[13] ),
    .A1(\top0.periodTop[13] ),
    .S(_07125_),
    .X(_07133_));
 sky130_fd_sc_hd__clkbuf_1 _15016_ (.A(_07133_),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _15017_ (.A0(\spi0.data_packed[14] ),
    .A1(\top0.periodTop[14] ),
    .S(_07125_),
    .X(_07134_));
 sky130_fd_sc_hd__clkbuf_1 _15018_ (.A(_07134_),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _15019_ (.A0(\spi0.data_packed[15] ),
    .A1(net1006),
    .S(_07125_),
    .X(_07135_));
 sky130_fd_sc_hd__clkbuf_1 _15020_ (.A(_07135_),
    .X(_00116_));
 sky130_fd_sc_hd__or2_2 _15021_ (.A(net431),
    .B(net441),
    .X(_07136_));
 sky130_fd_sc_hd__or3_2 _15022_ (.A(\top0.pid_d.state[0] ),
    .B(\top0.pid_d.state[3] ),
    .C(_07136_),
    .X(_07137_));
 sky130_fd_sc_hd__clkbuf_4 _15023_ (.A(_07137_),
    .X(_07138_));
 sky130_fd_sc_hd__o21a_2 _15024_ (.A1(net435),
    .A2(_07138_),
    .B1(_05443_),
    .X(_07139_));
 sky130_fd_sc_hd__clkbuf_4 _15025_ (.A(_07139_),
    .X(_07140_));
 sky130_fd_sc_hd__nor3_2 _15026_ (.A(\top0.pid_d.state[0] ),
    .B(\top0.pid_d.state[3] ),
    .C(_07136_),
    .Y(_07141_));
 sky130_fd_sc_hd__and4b_1 _15027_ (.A_N(net437),
    .B(net432),
    .C(_05442_),
    .D(_07141_),
    .X(_07142_));
 sky130_fd_sc_hd__buf_2 _15028_ (.A(_07142_),
    .X(_07143_));
 sky130_fd_sc_hd__clkbuf_4 _15029_ (.A(_07143_),
    .X(_07144_));
 sky130_fd_sc_hd__a22o_1 _15030_ (.A1(net968),
    .A2(_07140_),
    .B1(_07144_),
    .B2(\top0.pid_d.curr_int[0] ),
    .X(_00117_));
 sky130_fd_sc_hd__a22o_1 _15031_ (.A1(\top0.pid_d.prev_int[1] ),
    .A2(_07140_),
    .B1(_07144_),
    .B2(\top0.pid_d.curr_int[1] ),
    .X(_00118_));
 sky130_fd_sc_hd__a22o_1 _15032_ (.A1(net971),
    .A2(_07140_),
    .B1(_07144_),
    .B2(\top0.pid_d.curr_int[2] ),
    .X(_00119_));
 sky130_fd_sc_hd__a22o_1 _15033_ (.A1(\top0.pid_d.prev_int[3] ),
    .A2(_07140_),
    .B1(_07144_),
    .B2(\top0.pid_d.curr_int[3] ),
    .X(_00120_));
 sky130_fd_sc_hd__a22o_1 _15034_ (.A1(net964),
    .A2(_07140_),
    .B1(_07144_),
    .B2(\top0.pid_d.curr_int[4] ),
    .X(_00121_));
 sky130_fd_sc_hd__a22o_1 _15035_ (.A1(\top0.pid_d.prev_int[5] ),
    .A2(_07140_),
    .B1(_07144_),
    .B2(\top0.pid_d.curr_int[5] ),
    .X(_00122_));
 sky130_fd_sc_hd__a22o_1 _15036_ (.A1(net938),
    .A2(_07140_),
    .B1(_07144_),
    .B2(\top0.pid_d.curr_int[6] ),
    .X(_00123_));
 sky130_fd_sc_hd__a22o_1 _15037_ (.A1(\top0.pid_d.prev_int[7] ),
    .A2(_07140_),
    .B1(_07144_),
    .B2(net911),
    .X(_00124_));
 sky130_fd_sc_hd__a22o_1 _15038_ (.A1(\top0.pid_d.prev_int[8] ),
    .A2(_07140_),
    .B1(_07144_),
    .B2(\top0.pid_d.curr_int[8] ),
    .X(_00125_));
 sky130_fd_sc_hd__a22o_1 _15039_ (.A1(net990),
    .A2(_07140_),
    .B1(_07144_),
    .B2(\top0.pid_d.curr_int[9] ),
    .X(_00126_));
 sky130_fd_sc_hd__a22o_1 _15040_ (.A1(\top0.pid_d.prev_int[10] ),
    .A2(_07139_),
    .B1(_07143_),
    .B2(net828),
    .X(_00127_));
 sky130_fd_sc_hd__a22o_1 _15041_ (.A1(\top0.pid_d.prev_int[11] ),
    .A2(_07139_),
    .B1(_07143_),
    .B2(\top0.pid_d.curr_int[11] ),
    .X(_00128_));
 sky130_fd_sc_hd__a22o_1 _15042_ (.A1(\top0.pid_d.prev_int[12] ),
    .A2(_07139_),
    .B1(_07143_),
    .B2(net978),
    .X(_00129_));
 sky130_fd_sc_hd__a22o_1 _15043_ (.A1(net917),
    .A2(_07139_),
    .B1(_07143_),
    .B2(\top0.pid_d.curr_int[13] ),
    .X(_00130_));
 sky130_fd_sc_hd__a22o_1 _15044_ (.A1(net941),
    .A2(_07139_),
    .B1(_07143_),
    .B2(\top0.pid_d.curr_int[14] ),
    .X(_00131_));
 sky130_fd_sc_hd__a22o_1 _15045_ (.A1(net815),
    .A2(_07139_),
    .B1(_07143_),
    .B2(\top0.pid_d.curr_int[15] ),
    .X(_00132_));
 sky130_fd_sc_hd__and2_1 _15046_ (.A(net520),
    .B(net485),
    .X(_07145_));
 sky130_fd_sc_hd__nand2_1 _15047_ (.A(net517),
    .B(net490),
    .Y(_07146_));
 sky130_fd_sc_hd__nand2_1 _15048_ (.A(net514),
    .B(net494),
    .Y(_07147_));
 sky130_fd_sc_hd__xor2_1 _15049_ (.A(_07146_),
    .B(_07147_),
    .X(_07148_));
 sky130_fd_sc_hd__xnor2_2 _15050_ (.A(_07145_),
    .B(_07148_),
    .Y(_07149_));
 sky130_fd_sc_hd__nand2_1 _15051_ (.A(net531),
    .B(net471),
    .Y(_07150_));
 sky130_fd_sc_hd__nand2_1 _15052_ (.A(net528),
    .B(net475),
    .Y(_07151_));
 sky130_fd_sc_hd__nand2_1 _15053_ (.A(net534),
    .B(net470),
    .Y(_07152_));
 sky130_fd_sc_hd__o21ai_1 _15054_ (.A1(_07150_),
    .A2(_07151_),
    .B1(_07152_),
    .Y(_07153_));
 sky130_fd_sc_hd__a21bo_1 _15055_ (.A1(_07150_),
    .A2(_07151_),
    .B1_N(_07153_),
    .X(_07154_));
 sky130_fd_sc_hd__nand2_1 _15056_ (.A(net531),
    .B(net470),
    .Y(_07155_));
 sky130_fd_sc_hd__nand2_1 _15057_ (.A(net528),
    .B(net471),
    .Y(_07156_));
 sky130_fd_sc_hd__nand2_1 _15058_ (.A(net526),
    .B(net475),
    .Y(_07157_));
 sky130_fd_sc_hd__xnor2_1 _15059_ (.A(_07156_),
    .B(_07157_),
    .Y(_07158_));
 sky130_fd_sc_hd__xnor2_2 _15060_ (.A(_07155_),
    .B(_07158_),
    .Y(_07159_));
 sky130_fd_sc_hd__xnor2_1 _15061_ (.A(_07154_),
    .B(_07159_),
    .Y(_07160_));
 sky130_fd_sc_hd__xnor2_1 _15062_ (.A(_07149_),
    .B(_07160_),
    .Y(_07161_));
 sky130_fd_sc_hd__nand2_2 _15063_ (.A(net522),
    .B(net484),
    .Y(_07162_));
 sky130_fd_sc_hd__nand2_2 _15064_ (.A(net517),
    .B(net493),
    .Y(_07163_));
 sky130_fd_sc_hd__nand2_2 _15065_ (.A(net520),
    .B(net489),
    .Y(_07164_));
 sky130_fd_sc_hd__xnor2_2 _15066_ (.A(_07163_),
    .B(_07164_),
    .Y(_07165_));
 sky130_fd_sc_hd__xnor2_4 _15067_ (.A(_07162_),
    .B(_07165_),
    .Y(_07166_));
 sky130_fd_sc_hd__xnor2_1 _15068_ (.A(_07150_),
    .B(_07151_),
    .Y(_07167_));
 sky130_fd_sc_hd__xnor2_2 _15069_ (.A(_07152_),
    .B(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__nand2_2 _15070_ (.A(net533),
    .B(net475),
    .Y(_07169_));
 sky130_fd_sc_hd__nand2_2 _15071_ (.A(\top0.pid_q.mult0.a[2] ),
    .B(net471),
    .Y(_07170_));
 sky130_fd_sc_hd__nand2_1 _15072_ (.A(_07169_),
    .B(_07170_),
    .Y(_07171_));
 sky130_fd_sc_hd__nor2_1 _15073_ (.A(_07169_),
    .B(_07170_),
    .Y(_07172_));
 sky130_fd_sc_hd__a31o_1 _15074_ (.A1(net539),
    .A2(net470),
    .A3(_07171_),
    .B1(_07172_),
    .X(_07173_));
 sky130_fd_sc_hd__o21bai_1 _15075_ (.A1(_07166_),
    .A2(_07168_),
    .B1_N(_07173_),
    .Y(_07174_));
 sky130_fd_sc_hd__a21bo_1 _15076_ (.A1(_07166_),
    .A2(_07168_),
    .B1_N(_07174_),
    .X(_07175_));
 sky130_fd_sc_hd__xor2_1 _15077_ (.A(_07161_),
    .B(_07175_),
    .X(_07176_));
 sky130_fd_sc_hd__nand2_1 _15078_ (.A(net537),
    .B(net462),
    .Y(_07177_));
 sky130_fd_sc_hd__nand2_1 _15079_ (.A(net535),
    .B(net465),
    .Y(_07178_));
 sky130_fd_sc_hd__nand2_1 _15080_ (.A(net540),
    .B(net460),
    .Y(_07179_));
 sky130_fd_sc_hd__o22a_1 _15081_ (.A1(net540),
    .A2(_07178_),
    .B1(_07179_),
    .B2(net464),
    .X(_07180_));
 sky130_fd_sc_hd__xnor2_1 _15082_ (.A(net535),
    .B(net460),
    .Y(_07181_));
 sky130_fd_sc_hd__inv_2 _15083_ (.A(net541),
    .Y(_07182_));
 sky130_fd_sc_hd__a2bb2o_1 _15084_ (.A1_N(net460),
    .A2_N(net464),
    .B1(_07178_),
    .B2(_07182_),
    .X(_07183_));
 sky130_fd_sc_hd__a32o_1 _15085_ (.A1(net540),
    .A2(net465),
    .A3(_07181_),
    .B1(_07177_),
    .B2(_07183_),
    .X(_07184_));
 sky130_fd_sc_hd__o21ba_1 _15086_ (.A1(_07177_),
    .A2(_07180_),
    .B1_N(_07184_),
    .X(_07185_));
 sky130_fd_sc_hd__nand2_1 _15087_ (.A(_07176_),
    .B(_07185_),
    .Y(_07186_));
 sky130_fd_sc_hd__and2_1 _15088_ (.A(net537),
    .B(net460),
    .X(_07187_));
 sky130_fd_sc_hd__nand2_1 _15089_ (.A(net535),
    .B(net462),
    .Y(_07188_));
 sky130_fd_sc_hd__nand2_1 _15090_ (.A(net531),
    .B(net464),
    .Y(_07189_));
 sky130_fd_sc_hd__xor2_1 _15091_ (.A(_07188_),
    .B(_07189_),
    .X(_07190_));
 sky130_fd_sc_hd__xnor2_2 _15092_ (.A(_07187_),
    .B(_07190_),
    .Y(_07191_));
 sky130_fd_sc_hd__o21a_1 _15093_ (.A1(_07177_),
    .A2(_07178_),
    .B1(_07179_),
    .X(_07192_));
 sky130_fd_sc_hd__a21o_1 _15094_ (.A1(_07177_),
    .A2(_07178_),
    .B1(_07192_),
    .X(_07193_));
 sky130_fd_sc_hd__nand2_1 _15095_ (.A(net540),
    .B(net457),
    .Y(_07194_));
 sky130_fd_sc_hd__xor2_1 _15096_ (.A(_07193_),
    .B(_07194_),
    .X(_07195_));
 sky130_fd_sc_hd__xnor2_1 _15097_ (.A(_07191_),
    .B(_07195_),
    .Y(_07196_));
 sky130_fd_sc_hd__nand2_1 _15098_ (.A(net528),
    .B(net470),
    .Y(_07197_));
 sky130_fd_sc_hd__nand2_1 _15099_ (.A(net525),
    .B(net471),
    .Y(_07198_));
 sky130_fd_sc_hd__nand2_1 _15100_ (.A(net522),
    .B(net475),
    .Y(_07199_));
 sky130_fd_sc_hd__xor2_1 _15101_ (.A(_07198_),
    .B(_07199_),
    .X(_07200_));
 sky130_fd_sc_hd__xnor2_2 _15102_ (.A(_07197_),
    .B(_07200_),
    .Y(_07201_));
 sky130_fd_sc_hd__o21ai_1 _15103_ (.A1(_07156_),
    .A2(_07157_),
    .B1(_07155_),
    .Y(_07202_));
 sky130_fd_sc_hd__a21bo_1 _15104_ (.A1(_07156_),
    .A2(_07157_),
    .B1_N(_07202_),
    .X(_07203_));
 sky130_fd_sc_hd__nand2_2 _15105_ (.A(net494),
    .B(net511),
    .Y(_07204_));
 sky130_fd_sc_hd__nand2_1 _15106_ (.A(net514),
    .B(net490),
    .Y(_07205_));
 sky130_fd_sc_hd__nand2_1 _15107_ (.A(net517),
    .B(net485),
    .Y(_07206_));
 sky130_fd_sc_hd__xnor2_1 _15108_ (.A(_07205_),
    .B(_07206_),
    .Y(_07207_));
 sky130_fd_sc_hd__xnor2_2 _15109_ (.A(_07204_),
    .B(_07207_),
    .Y(_07208_));
 sky130_fd_sc_hd__xor2_1 _15110_ (.A(_07203_),
    .B(_07208_),
    .X(_07209_));
 sky130_fd_sc_hd__xnor2_2 _15111_ (.A(_07201_),
    .B(_07209_),
    .Y(_07210_));
 sky130_fd_sc_hd__o21ai_1 _15112_ (.A1(_07149_),
    .A2(_07159_),
    .B1(_07154_),
    .Y(_07211_));
 sky130_fd_sc_hd__nand2_1 _15113_ (.A(_07149_),
    .B(_07159_),
    .Y(_07212_));
 sky130_fd_sc_hd__and2_4 _15114_ (.A(net462),
    .B(net464),
    .X(_07213_));
 sky130_fd_sc_hd__nand4_2 _15115_ (.A(net540),
    .B(net538),
    .C(_07181_),
    .D(_07213_),
    .Y(_07214_));
 sky130_fd_sc_hd__nand3_1 _15116_ (.A(_07211_),
    .B(_07212_),
    .C(_07214_),
    .Y(_07215_));
 sky130_fd_sc_hd__a21o_1 _15117_ (.A1(_07211_),
    .A2(_07212_),
    .B1(_07214_),
    .X(_07216_));
 sky130_fd_sc_hd__nand3_1 _15118_ (.A(_07210_),
    .B(_07215_),
    .C(_07216_),
    .Y(_07217_));
 sky130_fd_sc_hd__a21o_1 _15119_ (.A1(_07215_),
    .A2(_07216_),
    .B1(_07210_),
    .X(_07218_));
 sky130_fd_sc_hd__and3_1 _15120_ (.A(_07196_),
    .B(_07217_),
    .C(_07218_),
    .X(_07219_));
 sky130_fd_sc_hd__clkbuf_2 _15121_ (.A(_07219_),
    .X(_07220_));
 sky130_fd_sc_hd__a21oi_1 _15122_ (.A1(_07217_),
    .A2(_07218_),
    .B1(_07196_),
    .Y(_07221_));
 sky130_fd_sc_hd__nor2_2 _15123_ (.A(_07161_),
    .B(_07175_),
    .Y(_07222_));
 sky130_fd_sc_hd__and4_1 _15124_ (.A(net517),
    .B(net514),
    .C(net494),
    .D(net490),
    .X(_07223_));
 sky130_fd_sc_hd__a22o_1 _15125_ (.A1(net514),
    .A2(net494),
    .B1(net490),
    .B2(net517),
    .X(_07224_));
 sky130_fd_sc_hd__o21a_1 _15126_ (.A1(_07145_),
    .A2(_07223_),
    .B1(_07224_),
    .X(_07225_));
 sky130_fd_sc_hd__inv_2 _15127_ (.A(_07225_),
    .Y(_07226_));
 sky130_fd_sc_hd__or2_1 _15128_ (.A(net489),
    .B(net484),
    .X(_07227_));
 sky130_fd_sc_hd__and2_1 _15129_ (.A(net489),
    .B(net484),
    .X(_07228_));
 sky130_fd_sc_hd__a21o_1 _15130_ (.A1(net517),
    .A2(net493),
    .B1(_07228_),
    .X(_07229_));
 sky130_fd_sc_hd__inv_2 _15131_ (.A(net521),
    .Y(_07230_));
 sky130_fd_sc_hd__a31o_1 _15132_ (.A1(net522),
    .A2(_07227_),
    .A3(_07229_),
    .B1(_07230_),
    .X(_07231_));
 sky130_fd_sc_hd__or3_1 _15133_ (.A(net520),
    .B(_07162_),
    .C(_07163_),
    .X(_07232_));
 sky130_fd_sc_hd__inv_2 _15134_ (.A(net479),
    .Y(_07233_));
 sky130_fd_sc_hd__a21o_1 _15135_ (.A1(_07231_),
    .A2(_07232_),
    .B1(_07233_),
    .X(_07234_));
 sky130_fd_sc_hd__xnor2_2 _15136_ (.A(_07226_),
    .B(_07234_),
    .Y(_07235_));
 sky130_fd_sc_hd__xnor2_2 _15137_ (.A(_07222_),
    .B(_07235_),
    .Y(_07236_));
 sky130_fd_sc_hd__or3b_1 _15138_ (.A(_07220_),
    .B(_07221_),
    .C_N(_07236_),
    .X(_07237_));
 sky130_fd_sc_hd__or2_1 _15139_ (.A(_07220_),
    .B(_07221_),
    .X(_07238_));
 sky130_fd_sc_hd__and2b_1 _15140_ (.A_N(_07236_),
    .B(_07238_),
    .X(_07239_));
 sky130_fd_sc_hd__a21o_1 _15141_ (.A1(_07186_),
    .A2(_07237_),
    .B1(_07239_),
    .X(_07240_));
 sky130_fd_sc_hd__inv_2 _15142_ (.A(net523),
    .Y(_07241_));
 sky130_fd_sc_hd__o21a_1 _15143_ (.A1(_07163_),
    .A2(_07164_),
    .B1(_07162_),
    .X(_07242_));
 sky130_fd_sc_hd__a21oi_2 _15144_ (.A1(_07163_),
    .A2(_07164_),
    .B1(_07242_),
    .Y(_07243_));
 sky130_fd_sc_hd__inv_2 _15145_ (.A(_07243_),
    .Y(_07244_));
 sky130_fd_sc_hd__nor2_1 _15146_ (.A(_07241_),
    .B(_07244_),
    .Y(_07245_));
 sky130_fd_sc_hd__a21o_1 _15147_ (.A1(_07230_),
    .A2(_07225_),
    .B1(_07222_),
    .X(_07246_));
 sky130_fd_sc_hd__o211a_1 _15148_ (.A1(_07222_),
    .A2(_07245_),
    .B1(_07226_),
    .C1(net520),
    .X(_07247_));
 sky130_fd_sc_hd__a21o_1 _15149_ (.A1(_07245_),
    .A2(_07246_),
    .B1(_07247_),
    .X(_07248_));
 sky130_fd_sc_hd__nand2_1 _15150_ (.A(net521),
    .B(net480),
    .Y(_07249_));
 sky130_fd_sc_hd__and3_1 _15151_ (.A(_07222_),
    .B(_07225_),
    .C(_07249_),
    .X(_07250_));
 sky130_fd_sc_hd__a21oi_2 _15152_ (.A1(net480),
    .A2(_07248_),
    .B1(_07250_),
    .Y(_07251_));
 sky130_fd_sc_hd__nand2_1 _15153_ (.A(_07211_),
    .B(_07212_),
    .Y(_07252_));
 sky130_fd_sc_hd__o21ai_1 _15154_ (.A1(_07252_),
    .A2(_07210_),
    .B1(_07214_),
    .Y(_07253_));
 sky130_fd_sc_hd__nand2_1 _15155_ (.A(_07252_),
    .B(_07210_),
    .Y(_07254_));
 sky130_fd_sc_hd__nand2_2 _15156_ (.A(_07253_),
    .B(_07254_),
    .Y(_07255_));
 sky130_fd_sc_hd__nand2_1 _15157_ (.A(_07204_),
    .B(_07205_),
    .Y(_07256_));
 sky130_fd_sc_hd__nor2_1 _15158_ (.A(_07204_),
    .B(_07205_),
    .Y(_07257_));
 sky130_fd_sc_hd__a31o_1 _15159_ (.A1(net517),
    .A2(net485),
    .A3(_07256_),
    .B1(_07257_),
    .X(_07258_));
 sky130_fd_sc_hd__nor2_1 _15160_ (.A(_07230_),
    .B(_07226_),
    .Y(_07259_));
 sky130_fd_sc_hd__xnor2_1 _15161_ (.A(net517),
    .B(_07259_),
    .Y(_07260_));
 sky130_fd_sc_hd__nor2_1 _15162_ (.A(_07233_),
    .B(_07260_),
    .Y(_07261_));
 sky130_fd_sc_hd__xnor2_1 _15163_ (.A(_07258_),
    .B(_07261_),
    .Y(_07262_));
 sky130_fd_sc_hd__xnor2_1 _15164_ (.A(_07255_),
    .B(_07262_),
    .Y(_07263_));
 sky130_fd_sc_hd__nand2_1 _15165_ (.A(_07203_),
    .B(_07208_),
    .Y(_07264_));
 sky130_fd_sc_hd__nor2_1 _15166_ (.A(_07203_),
    .B(_07208_),
    .Y(_07265_));
 sky130_fd_sc_hd__a21oi_4 _15167_ (.A1(_07201_),
    .A2(_07264_),
    .B1(_07265_),
    .Y(_07266_));
 sky130_fd_sc_hd__nand2_2 _15168_ (.A(net520),
    .B(net475),
    .Y(_07267_));
 sky130_fd_sc_hd__nand2_2 _15169_ (.A(net522),
    .B(net471),
    .Y(_07268_));
 sky130_fd_sc_hd__nand2_1 _15170_ (.A(net526),
    .B(net470),
    .Y(_07269_));
 sky130_fd_sc_hd__xnor2_2 _15171_ (.A(_07268_),
    .B(_07269_),
    .Y(_07270_));
 sky130_fd_sc_hd__xnor2_4 _15172_ (.A(_07267_),
    .B(_07270_),
    .Y(_07271_));
 sky130_fd_sc_hd__o21ai_1 _15173_ (.A1(_07198_),
    .A2(_07199_),
    .B1(_07197_),
    .Y(_07272_));
 sky130_fd_sc_hd__a21bo_1 _15174_ (.A1(_07198_),
    .A2(_07199_),
    .B1_N(_07272_),
    .X(_07273_));
 sky130_fd_sc_hd__and2_2 _15175_ (.A(net489),
    .B(net511),
    .X(_07274_));
 sky130_fd_sc_hd__nand2_1 _15176_ (.A(net514),
    .B(net485),
    .Y(_07275_));
 sky130_fd_sc_hd__and2_1 _15177_ (.A(net493),
    .B(net508),
    .X(_07276_));
 sky130_fd_sc_hd__xnor2_1 _15178_ (.A(_07275_),
    .B(_07276_),
    .Y(_07277_));
 sky130_fd_sc_hd__xnor2_2 _15179_ (.A(_07274_),
    .B(_07277_),
    .Y(_07278_));
 sky130_fd_sc_hd__xnor2_2 _15180_ (.A(_07273_),
    .B(_07278_),
    .Y(_07279_));
 sky130_fd_sc_hd__xnor2_4 _15181_ (.A(_07271_),
    .B(_07279_),
    .Y(_07280_));
 sky130_fd_sc_hd__xnor2_4 _15182_ (.A(_07266_),
    .B(_07280_),
    .Y(_07281_));
 sky130_fd_sc_hd__nand2_2 _15183_ (.A(net535),
    .B(net460),
    .Y(_07282_));
 sky130_fd_sc_hd__nand2_1 _15184_ (.A(net531),
    .B(net462),
    .Y(_07283_));
 sky130_fd_sc_hd__nand2_1 _15185_ (.A(net528),
    .B(net464),
    .Y(_07284_));
 sky130_fd_sc_hd__xor2_2 _15186_ (.A(_07283_),
    .B(_07284_),
    .X(_07285_));
 sky130_fd_sc_hd__xnor2_4 _15187_ (.A(_07282_),
    .B(_07285_),
    .Y(_07286_));
 sky130_fd_sc_hd__o21ba_1 _15188_ (.A1(_07188_),
    .A2(_07189_),
    .B1_N(_07187_),
    .X(_07287_));
 sky130_fd_sc_hd__a21oi_2 _15189_ (.A1(_07188_),
    .A2(_07189_),
    .B1(_07287_),
    .Y(_07288_));
 sky130_fd_sc_hd__nand2_2 _15190_ (.A(net538),
    .B(net457),
    .Y(_07289_));
 sky130_fd_sc_hd__nand2_2 _15191_ (.A(net540),
    .B(net454),
    .Y(_07290_));
 sky130_fd_sc_hd__xor2_4 _15192_ (.A(_07289_),
    .B(_07290_),
    .X(_07291_));
 sky130_fd_sc_hd__xnor2_2 _15193_ (.A(_07288_),
    .B(_07291_),
    .Y(_07292_));
 sky130_fd_sc_hd__xnor2_4 _15194_ (.A(_07286_),
    .B(_07292_),
    .Y(_07293_));
 sky130_fd_sc_hd__or2_1 _15195_ (.A(_07193_),
    .B(_07191_),
    .X(_07294_));
 sky130_fd_sc_hd__and2_1 _15196_ (.A(_07193_),
    .B(_07191_),
    .X(_07295_));
 sky130_fd_sc_hd__a21oi_2 _15197_ (.A1(_07194_),
    .A2(_07294_),
    .B1(_07295_),
    .Y(_07296_));
 sky130_fd_sc_hd__xor2_2 _15198_ (.A(_07293_),
    .B(_07296_),
    .X(_07297_));
 sky130_fd_sc_hd__xnor2_4 _15199_ (.A(_07281_),
    .B(_07297_),
    .Y(_07298_));
 sky130_fd_sc_hd__xnor2_1 _15200_ (.A(_07220_),
    .B(_07298_),
    .Y(_07299_));
 sky130_fd_sc_hd__xnor2_1 _15201_ (.A(_07263_),
    .B(_07299_),
    .Y(_07300_));
 sky130_fd_sc_hd__xnor2_1 _15202_ (.A(_07251_),
    .B(_07300_),
    .Y(_07301_));
 sky130_fd_sc_hd__xor2_1 _15203_ (.A(_07240_),
    .B(_07301_),
    .X(_07302_));
 sky130_fd_sc_hd__xnor2_2 _15204_ (.A(_07168_),
    .B(_07173_),
    .Y(_07303_));
 sky130_fd_sc_hd__xnor2_4 _15205_ (.A(_07166_),
    .B(_07303_),
    .Y(_07304_));
 sky130_fd_sc_hd__nand2_1 _15206_ (.A(\top0.pid_q.mult0.a[2] ),
    .B(net475),
    .Y(_07305_));
 sky130_fd_sc_hd__nand2_1 _15207_ (.A(net539),
    .B(net471),
    .Y(_07306_));
 sky130_fd_sc_hd__nand2_1 _15208_ (.A(net542),
    .B(net470),
    .Y(_07307_));
 sky130_fd_sc_hd__o21a_1 _15209_ (.A1(_07305_),
    .A2(_07306_),
    .B1(_07307_),
    .X(_07308_));
 sky130_fd_sc_hd__a21o_1 _15210_ (.A1(_07305_),
    .A2(_07306_),
    .B1(_07308_),
    .X(_07309_));
 sky130_fd_sc_hd__nand2_2 _15211_ (.A(net539),
    .B(net470),
    .Y(_07310_));
 sky130_fd_sc_hd__xnor2_2 _15212_ (.A(_07169_),
    .B(_07170_),
    .Y(_07311_));
 sky130_fd_sc_hd__xnor2_4 _15213_ (.A(_07310_),
    .B(_07311_),
    .Y(_07312_));
 sky130_fd_sc_hd__nand2_2 _15214_ (.A(net520),
    .B(net493),
    .Y(_07313_));
 sky130_fd_sc_hd__nand2_1 _15215_ (.A(net525),
    .B(net487),
    .Y(_07314_));
 sky130_fd_sc_hd__nand2_1 _15216_ (.A(net522),
    .B(net491),
    .Y(_07315_));
 sky130_fd_sc_hd__xnor2_1 _15217_ (.A(_07314_),
    .B(_07315_),
    .Y(_07316_));
 sky130_fd_sc_hd__xnor2_1 _15218_ (.A(_07313_),
    .B(_07316_),
    .Y(_07317_));
 sky130_fd_sc_hd__o21a_1 _15219_ (.A1(_07309_),
    .A2(_07312_),
    .B1(_07317_),
    .X(_07318_));
 sky130_fd_sc_hd__a21oi_4 _15220_ (.A1(_07309_),
    .A2(_07312_),
    .B1(_07318_),
    .Y(_07319_));
 sky130_fd_sc_hd__inv_2 _15221_ (.A(net527),
    .Y(_07320_));
 sky130_fd_sc_hd__nor2_2 _15222_ (.A(_07313_),
    .B(_07315_),
    .Y(_07321_));
 sky130_fd_sc_hd__nand2_1 _15223_ (.A(_07313_),
    .B(_07315_),
    .Y(_07322_));
 sky130_fd_sc_hd__o21ai_1 _15224_ (.A1(net487),
    .A2(_07321_),
    .B1(_07322_),
    .Y(_07323_));
 sky130_fd_sc_hd__nor2_1 _15225_ (.A(_07320_),
    .B(_07323_),
    .Y(_07324_));
 sky130_fd_sc_hd__a21o_1 _15226_ (.A1(_07304_),
    .A2(_07319_),
    .B1(_07324_),
    .X(_07325_));
 sky130_fd_sc_hd__a22o_1 _15227_ (.A1(_07304_),
    .A2(_07319_),
    .B1(_07243_),
    .B2(_07241_),
    .X(_07326_));
 sky130_fd_sc_hd__a32o_1 _15228_ (.A1(net522),
    .A2(_07244_),
    .A3(_07325_),
    .B1(_07326_),
    .B2(_07324_),
    .X(_07327_));
 sky130_fd_sc_hd__and2_1 _15229_ (.A(_07304_),
    .B(_07319_),
    .X(_07328_));
 sky130_fd_sc_hd__o211a_1 _15230_ (.A1(_07241_),
    .A2(_07233_),
    .B1(_07328_),
    .C1(_07243_),
    .X(_07329_));
 sky130_fd_sc_hd__a21oi_2 _15231_ (.A1(net481),
    .A2(_07327_),
    .B1(_07329_),
    .Y(_07330_));
 sky130_fd_sc_hd__xor2_1 _15232_ (.A(_07186_),
    .B(_07236_),
    .X(_07331_));
 sky130_fd_sc_hd__xnor2_2 _15233_ (.A(_07238_),
    .B(_07331_),
    .Y(_07332_));
 sky130_fd_sc_hd__xnor2_1 _15234_ (.A(_07176_),
    .B(_07185_),
    .Y(_07333_));
 sky130_fd_sc_hd__nor2_1 _15235_ (.A(_07304_),
    .B(_07319_),
    .Y(_07334_));
 sky130_fd_sc_hd__nand2_2 _15236_ (.A(net537),
    .B(net464),
    .Y(_07335_));
 sky130_fd_sc_hd__nand2_1 _15237_ (.A(net541),
    .B(net462),
    .Y(_07336_));
 sky130_fd_sc_hd__xnor2_1 _15238_ (.A(_07335_),
    .B(_07336_),
    .Y(_07337_));
 sky130_fd_sc_hd__a21o_1 _15239_ (.A1(net520),
    .A2(net493),
    .B1(_07228_),
    .X(_07338_));
 sky130_fd_sc_hd__a31o_1 _15240_ (.A1(net525),
    .A2(_07227_),
    .A3(_07338_),
    .B1(_07241_),
    .X(_07339_));
 sky130_fd_sc_hd__or3_1 _15241_ (.A(net522),
    .B(_07314_),
    .C(_07313_),
    .X(_07340_));
 sky130_fd_sc_hd__a21o_1 _15242_ (.A1(_07339_),
    .A2(_07340_),
    .B1(_07233_),
    .X(_07341_));
 sky130_fd_sc_hd__xnor2_1 _15243_ (.A(_07243_),
    .B(_07341_),
    .Y(_07342_));
 sky130_fd_sc_hd__or4b_1 _15244_ (.A(_07328_),
    .B(_07334_),
    .C(_07337_),
    .D_N(_07342_),
    .X(_07343_));
 sky130_fd_sc_hd__xor2_2 _15245_ (.A(_07304_),
    .B(_07319_),
    .X(_07344_));
 sky130_fd_sc_hd__xor2_2 _15246_ (.A(_07335_),
    .B(_07336_),
    .X(_07345_));
 sky130_fd_sc_hd__and3_1 _15247_ (.A(_07304_),
    .B(_07319_),
    .C(_07342_),
    .X(_07346_));
 sky130_fd_sc_hd__a21oi_1 _15248_ (.A1(_07304_),
    .A2(_07319_),
    .B1(_07342_),
    .Y(_07347_));
 sky130_fd_sc_hd__o2bb2a_1 _15249_ (.A1_N(_07344_),
    .A2_N(_07345_),
    .B1(_07346_),
    .B2(_07347_),
    .X(_07348_));
 sky130_fd_sc_hd__a21o_1 _15250_ (.A1(_07333_),
    .A2(_07343_),
    .B1(_07348_),
    .X(_07349_));
 sky130_fd_sc_hd__nand3_1 _15251_ (.A(_07330_),
    .B(_07332_),
    .C(_07349_),
    .Y(_07350_));
 sky130_fd_sc_hd__nand2_1 _15252_ (.A(_07332_),
    .B(_07349_),
    .Y(_07351_));
 sky130_fd_sc_hd__o21ai_1 _15253_ (.A1(_07332_),
    .A2(_07349_),
    .B1(_07330_),
    .Y(_07352_));
 sky130_fd_sc_hd__xnor2_1 _15254_ (.A(_07309_),
    .B(_07317_),
    .Y(_07353_));
 sky130_fd_sc_hd__xnor2_1 _15255_ (.A(_07312_),
    .B(_07353_),
    .Y(_07354_));
 sky130_fd_sc_hd__and4_1 _15256_ (.A(net542),
    .B(net539),
    .C(net471),
    .D(net475),
    .X(_07355_));
 sky130_fd_sc_hd__nand2_1 _15257_ (.A(net527),
    .B(net491),
    .Y(_07356_));
 sky130_fd_sc_hd__nand2_1 _15258_ (.A(net524),
    .B(net495),
    .Y(_07357_));
 sky130_fd_sc_hd__xor2_1 _15259_ (.A(_07356_),
    .B(_07357_),
    .X(_07358_));
 sky130_fd_sc_hd__nand2_1 _15260_ (.A(net1026),
    .B(net487),
    .Y(_07359_));
 sky130_fd_sc_hd__xnor2_2 _15261_ (.A(_07358_),
    .B(_07359_),
    .Y(_07360_));
 sky130_fd_sc_hd__xor2_1 _15262_ (.A(_07305_),
    .B(_07306_),
    .X(_07361_));
 sky130_fd_sc_hd__xnor2_1 _15263_ (.A(_07307_),
    .B(_07361_),
    .Y(_07362_));
 sky130_fd_sc_hd__o21a_1 _15264_ (.A1(_07355_),
    .A2(_07360_),
    .B1(_07362_),
    .X(_07363_));
 sky130_fd_sc_hd__a21o_1 _15265_ (.A1(_07355_),
    .A2(_07360_),
    .B1(_07363_),
    .X(_07364_));
 sky130_fd_sc_hd__nand2b_2 _15266_ (.A_N(_07354_),
    .B(_07364_),
    .Y(_07365_));
 sky130_fd_sc_hd__inv_2 _15267_ (.A(net484),
    .Y(_07366_));
 sky130_fd_sc_hd__nor2_1 _15268_ (.A(_07366_),
    .B(net479),
    .Y(_07367_));
 sky130_fd_sc_hd__a22o_1 _15269_ (.A1(net479),
    .A2(_07323_),
    .B1(_07367_),
    .B2(_07322_),
    .X(_07368_));
 sky130_fd_sc_hd__nand2_1 _15270_ (.A(net525),
    .B(net479),
    .Y(_07369_));
 sky130_fd_sc_hd__a22oi_2 _15271_ (.A1(net525),
    .A2(_07368_),
    .B1(_07369_),
    .B2(_07321_),
    .Y(_07370_));
 sky130_fd_sc_hd__nand2_1 _15272_ (.A(_07365_),
    .B(_07370_),
    .Y(_07371_));
 sky130_fd_sc_hd__and4_1 _15273_ (.A(net527),
    .B(net524),
    .C(net495),
    .D(net491),
    .X(_07372_));
 sky130_fd_sc_hd__a22o_1 _15274_ (.A1(net524),
    .A2(net495),
    .B1(net491),
    .B2(net527),
    .X(_07373_));
 sky130_fd_sc_hd__o211a_2 _15275_ (.A1(net487),
    .A2(_07372_),
    .B1(_07373_),
    .C1(net1026),
    .X(_07374_));
 sky130_fd_sc_hd__nor2_1 _15276_ (.A(_07365_),
    .B(_07370_),
    .Y(_07375_));
 sky130_fd_sc_hd__a31oi_4 _15277_ (.A1(net479),
    .A2(_07371_),
    .A3(_07374_),
    .B1(_07375_),
    .Y(_07376_));
 sky130_fd_sc_hd__inv_2 _15278_ (.A(_07376_),
    .Y(_07377_));
 sky130_fd_sc_hd__or4_1 _15279_ (.A(_07328_),
    .B(_07334_),
    .C(_07337_),
    .D(_07342_),
    .X(_07378_));
 sky130_fd_sc_hd__a211o_1 _15280_ (.A1(_07344_),
    .A2(_07345_),
    .B1(_07346_),
    .C1(_07347_),
    .X(_07379_));
 sky130_fd_sc_hd__nand3_1 _15281_ (.A(_07333_),
    .B(_07378_),
    .C(_07379_),
    .Y(_07380_));
 sky130_fd_sc_hd__a21o_1 _15282_ (.A1(_07378_),
    .A2(_07379_),
    .B1(_07333_),
    .X(_07381_));
 sky130_fd_sc_hd__o21ai_1 _15283_ (.A1(net525),
    .A2(_07374_),
    .B1(net479),
    .Y(_07382_));
 sky130_fd_sc_hd__o211a_1 _15284_ (.A1(_07233_),
    .A2(_07374_),
    .B1(_07322_),
    .C1(net487),
    .X(_07383_));
 sky130_fd_sc_hd__a21o_1 _15285_ (.A1(_07321_),
    .A2(_07374_),
    .B1(_07383_),
    .X(_07384_));
 sky130_fd_sc_hd__nand2_1 _15286_ (.A(net525),
    .B(_07366_),
    .Y(_07385_));
 sky130_fd_sc_hd__mux2_1 _15287_ (.A0(_07385_),
    .A1(net525),
    .S(_07374_),
    .X(_07386_));
 sky130_fd_sc_hd__o32a_1 _15288_ (.A1(_07320_),
    .A2(_07322_),
    .A3(_07374_),
    .B1(_07386_),
    .B2(_07321_),
    .X(_07387_));
 sky130_fd_sc_hd__nor2_1 _15289_ (.A(_07233_),
    .B(_07387_),
    .Y(_07388_));
 sky130_fd_sc_hd__a221o_1 _15290_ (.A1(_07321_),
    .A2(_07382_),
    .B1(_07384_),
    .B2(net525),
    .C1(_07388_),
    .X(_07389_));
 sky130_fd_sc_hd__xor2_2 _15291_ (.A(_07365_),
    .B(_07389_),
    .X(_07390_));
 sky130_fd_sc_hd__xnor2_2 _15292_ (.A(_07344_),
    .B(_07345_),
    .Y(_07391_));
 sky130_fd_sc_hd__nand2_1 _15293_ (.A(_07390_),
    .B(_07391_),
    .Y(_07392_));
 sky130_fd_sc_hd__nand2_1 _15294_ (.A(net542),
    .B(net464),
    .Y(_07393_));
 sky130_fd_sc_hd__xor2_1 _15295_ (.A(_07354_),
    .B(_07364_),
    .X(_07394_));
 sky130_fd_sc_hd__nor2_1 _15296_ (.A(_07393_),
    .B(_07394_),
    .Y(_07395_));
 sky130_fd_sc_hd__o21bai_1 _15297_ (.A1(_07390_),
    .A2(_07391_),
    .B1_N(_07395_),
    .Y(_07396_));
 sky130_fd_sc_hd__a22o_1 _15298_ (.A1(_07380_),
    .A2(_07381_),
    .B1(_07392_),
    .B2(_07396_),
    .X(_07397_));
 sky130_fd_sc_hd__and4_1 _15299_ (.A(_07380_),
    .B(_07381_),
    .C(_07392_),
    .D(_07396_),
    .X(_07398_));
 sky130_fd_sc_hd__a21o_1 _15300_ (.A1(_07377_),
    .A2(_07397_),
    .B1(_07398_),
    .X(_07399_));
 sky130_fd_sc_hd__a21o_1 _15301_ (.A1(_07351_),
    .A2(_07352_),
    .B1(_07399_),
    .X(_07400_));
 sky130_fd_sc_hd__a22o_1 _15302_ (.A1(net527),
    .A2(net495),
    .B1(net491),
    .B2(net1026),
    .X(_07401_));
 sky130_fd_sc_hd__and4_1 _15303_ (.A(net1026),
    .B(net527),
    .C(net495),
    .D(net491),
    .X(_07402_));
 sky130_fd_sc_hd__a21o_1 _15304_ (.A1(net487),
    .A2(_07401_),
    .B1(_07402_),
    .X(_07403_));
 sky130_fd_sc_hd__and2_1 _15305_ (.A(net533),
    .B(_07403_),
    .X(_07404_));
 sky130_fd_sc_hd__nand2_1 _15306_ (.A(net479),
    .B(_07404_),
    .Y(_07405_));
 sky130_fd_sc_hd__nor2_1 _15307_ (.A(net1026),
    .B(_07372_),
    .Y(_07406_));
 sky130_fd_sc_hd__nand2_1 _15308_ (.A(net539),
    .B(net478),
    .Y(_07407_));
 sky130_fd_sc_hd__and3_1 _15309_ (.A(net542),
    .B(net471),
    .C(_07407_),
    .X(_07408_));
 sky130_fd_sc_hd__a21oi_1 _15310_ (.A1(net542),
    .A2(net471),
    .B1(_07407_),
    .Y(_07409_));
 sky130_fd_sc_hd__nand2_1 _15311_ (.A(net1026),
    .B(net491),
    .Y(_07410_));
 sky130_fd_sc_hd__nand2_1 _15312_ (.A(net527),
    .B(net495),
    .Y(_07411_));
 sky130_fd_sc_hd__and2_1 _15313_ (.A(net533),
    .B(net487),
    .X(_07412_));
 sky130_fd_sc_hd__xor2_1 _15314_ (.A(_07411_),
    .B(_07412_),
    .X(_07413_));
 sky130_fd_sc_hd__xnor2_2 _15315_ (.A(_07410_),
    .B(_07413_),
    .Y(_07414_));
 sky130_fd_sc_hd__o21ba_1 _15316_ (.A1(_07408_),
    .A2(_07409_),
    .B1_N(_07414_),
    .X(_07415_));
 sky130_fd_sc_hd__xnor2_1 _15317_ (.A(_07362_),
    .B(_07360_),
    .Y(_07416_));
 sky130_fd_sc_hd__xnor2_1 _15318_ (.A(_07355_),
    .B(_07416_),
    .Y(_07417_));
 sky130_fd_sc_hd__nand2_1 _15319_ (.A(_07415_),
    .B(_07417_),
    .Y(_07418_));
 sky130_fd_sc_hd__a21o_1 _15320_ (.A1(net1026),
    .A2(net487),
    .B1(_07372_),
    .X(_07419_));
 sky130_fd_sc_hd__nand2_1 _15321_ (.A(_07373_),
    .B(_07419_),
    .Y(_07420_));
 sky130_fd_sc_hd__xor2_1 _15322_ (.A(net1026),
    .B(_07404_),
    .X(_07421_));
 sky130_fd_sc_hd__nand2_1 _15323_ (.A(net479),
    .B(_07421_),
    .Y(_07422_));
 sky130_fd_sc_hd__xnor2_1 _15324_ (.A(_07420_),
    .B(_07422_),
    .Y(_07423_));
 sky130_fd_sc_hd__and2_1 _15325_ (.A(_07418_),
    .B(_07423_),
    .X(_07424_));
 sky130_fd_sc_hd__xor2_1 _15326_ (.A(_07393_),
    .B(_07394_),
    .X(_07425_));
 sky130_fd_sc_hd__o21ba_1 _15327_ (.A1(_07418_),
    .A2(_07423_),
    .B1_N(_07425_),
    .X(_07426_));
 sky130_fd_sc_hd__o32a_1 _15328_ (.A1(_07374_),
    .A2(_07405_),
    .A3(_07406_),
    .B1(_07424_),
    .B2(_07426_),
    .X(_07427_));
 sky130_fd_sc_hd__xor2_1 _15329_ (.A(_07391_),
    .B(_07395_),
    .X(_07428_));
 sky130_fd_sc_hd__xnor2_1 _15330_ (.A(_07390_),
    .B(_07428_),
    .Y(_07429_));
 sky130_fd_sc_hd__nand2_1 _15331_ (.A(_07427_),
    .B(_07429_),
    .Y(_07430_));
 sky130_fd_sc_hd__xor2_1 _15332_ (.A(_07418_),
    .B(_07423_),
    .X(_07431_));
 sky130_fd_sc_hd__xnor2_1 _15333_ (.A(_07425_),
    .B(_07431_),
    .Y(_07432_));
 sky130_fd_sc_hd__xnor2_1 _15334_ (.A(net539),
    .B(net472),
    .Y(_07433_));
 sky130_fd_sc_hd__and2_1 _15335_ (.A(_07414_),
    .B(_07433_),
    .X(_07434_));
 sky130_fd_sc_hd__nor2_1 _15336_ (.A(_07414_),
    .B(_07433_),
    .Y(_07435_));
 sky130_fd_sc_hd__nand2_4 _15337_ (.A(net528),
    .B(net495),
    .Y(_07436_));
 sky130_fd_sc_hd__nand2_2 _15338_ (.A(net531),
    .B(net491),
    .Y(_07437_));
 sky130_fd_sc_hd__nand2_1 _15339_ (.A(net534),
    .B(net487),
    .Y(_07438_));
 sky130_fd_sc_hd__xnor2_2 _15340_ (.A(_07437_),
    .B(_07438_),
    .Y(_07439_));
 sky130_fd_sc_hd__xnor2_4 _15341_ (.A(_07436_),
    .B(_07439_),
    .Y(_07440_));
 sky130_fd_sc_hd__nand2_1 _15342_ (.A(net542),
    .B(net475),
    .Y(_07441_));
 sky130_fd_sc_hd__or4_2 _15343_ (.A(_07434_),
    .B(_07435_),
    .C(_07440_),
    .D(_07441_),
    .X(_07442_));
 sky130_fd_sc_hd__o21a_1 _15344_ (.A1(_07402_),
    .A2(_07412_),
    .B1(_07401_),
    .X(_07443_));
 sky130_fd_sc_hd__nor2_1 _15345_ (.A(_07436_),
    .B(_07437_),
    .Y(_07444_));
 sky130_fd_sc_hd__a21oi_1 _15346_ (.A1(_07436_),
    .A2(_07437_),
    .B1(_07366_),
    .Y(_07445_));
 sky130_fd_sc_hd__o21ai_2 _15347_ (.A1(_07444_),
    .A2(_07445_),
    .B1(net534),
    .Y(_07446_));
 sky130_fd_sc_hd__nor2_1 _15348_ (.A(net533),
    .B(_07402_),
    .Y(_07447_));
 sky130_fd_sc_hd__a31o_1 _15349_ (.A1(net533),
    .A2(net482),
    .A3(_07403_),
    .B1(_07447_),
    .X(_07448_));
 sky130_fd_sc_hd__a2bb2o_1 _15350_ (.A1_N(net482),
    .A2_N(_07443_),
    .B1(_07446_),
    .B2(_07448_),
    .X(_07449_));
 sky130_fd_sc_hd__xnor2_1 _15351_ (.A(_07415_),
    .B(_07417_),
    .Y(_07450_));
 sky130_fd_sc_hd__or4_1 _15352_ (.A(_07233_),
    .B(_07404_),
    .C(_07446_),
    .D(_07447_),
    .X(_07451_));
 sky130_fd_sc_hd__a21o_1 _15353_ (.A1(_07442_),
    .A2(_07451_),
    .B1(_07449_),
    .X(_07452_));
 sky130_fd_sc_hd__a22o_1 _15354_ (.A1(_07442_),
    .A2(_07449_),
    .B1(_07450_),
    .B2(_07452_),
    .X(_07453_));
 sky130_fd_sc_hd__nand2_1 _15355_ (.A(_07432_),
    .B(_07453_),
    .Y(_07454_));
 sky130_fd_sc_hd__and2_1 _15356_ (.A(net531),
    .B(net493),
    .X(_07455_));
 sky130_fd_sc_hd__clkbuf_2 _15357_ (.A(_07455_),
    .X(_07456_));
 sky130_fd_sc_hd__nand2_1 _15358_ (.A(net534),
    .B(net491),
    .Y(_07457_));
 sky130_fd_sc_hd__a21bo_1 _15359_ (.A1(net486),
    .A2(_07456_),
    .B1_N(_07457_),
    .X(_07458_));
 sky130_fd_sc_hd__o211a_1 _15360_ (.A1(net486),
    .A2(_07456_),
    .B1(_07458_),
    .C1(net537),
    .X(_07459_));
 sky130_fd_sc_hd__o2111a_1 _15361_ (.A1(net534),
    .A2(_07444_),
    .B1(_07446_),
    .C1(_07459_),
    .D1(net479),
    .X(_07460_));
 sky130_fd_sc_hd__xnor2_1 _15362_ (.A(net533),
    .B(_07446_),
    .Y(_07461_));
 sky130_fd_sc_hd__nand2_1 _15363_ (.A(net482),
    .B(_07461_),
    .Y(_07462_));
 sky130_fd_sc_hd__xnor2_1 _15364_ (.A(_07443_),
    .B(_07462_),
    .Y(_07463_));
 sky130_fd_sc_hd__xnor2_1 _15365_ (.A(_07442_),
    .B(_07463_),
    .Y(_07464_));
 sky130_fd_sc_hd__xnor2_1 _15366_ (.A(_07450_),
    .B(_07464_),
    .Y(_07465_));
 sky130_fd_sc_hd__o211ai_1 _15367_ (.A1(_07228_),
    .A2(_07456_),
    .B1(net537),
    .C1(_07227_),
    .Y(_07466_));
 sky130_fd_sc_hd__and4b_1 _15368_ (.A_N(net534),
    .B(net484),
    .C(_07456_),
    .D(net537),
    .X(_07467_));
 sky130_fd_sc_hd__a21o_1 _15369_ (.A1(net534),
    .A2(_07466_),
    .B1(_07467_),
    .X(_07468_));
 sky130_fd_sc_hd__nand2_1 _15370_ (.A(net479),
    .B(_07468_),
    .Y(_07469_));
 sky130_fd_sc_hd__o21a_1 _15371_ (.A1(_07436_),
    .A2(_07437_),
    .B1(_07438_),
    .X(_07470_));
 sky130_fd_sc_hd__a21oi_1 _15372_ (.A1(_07436_),
    .A2(_07437_),
    .B1(_07470_),
    .Y(_07471_));
 sky130_fd_sc_hd__xnor2_1 _15373_ (.A(_07469_),
    .B(_07471_),
    .Y(_07472_));
 sky130_fd_sc_hd__a22o_1 _15374_ (.A1(net534),
    .A2(net493),
    .B1(net489),
    .B2(net537),
    .X(_07473_));
 sky130_fd_sc_hd__and4_1 _15375_ (.A(net537),
    .B(net534),
    .C(net493),
    .D(net489),
    .X(_07474_));
 sky130_fd_sc_hd__a31o_1 _15376_ (.A1(net541),
    .A2(net484),
    .A3(_07473_),
    .B1(_07474_),
    .X(_07475_));
 sky130_fd_sc_hd__or3b_1 _15377_ (.A(_07182_),
    .B(_07233_),
    .C_N(_07475_),
    .X(_07476_));
 sky130_fd_sc_hd__and3_1 _15378_ (.A(net535),
    .B(net489),
    .C(_07456_),
    .X(_07477_));
 sky130_fd_sc_hd__or2_1 _15379_ (.A(net537),
    .B(_07477_),
    .X(_07478_));
 sky130_fd_sc_hd__nor3b_1 _15380_ (.A(_07476_),
    .B(_07459_),
    .C_N(_07478_),
    .Y(_07479_));
 sky130_fd_sc_hd__nand2_1 _15381_ (.A(net538),
    .B(net486),
    .Y(_07480_));
 sky130_fd_sc_hd__xor2_1 _15382_ (.A(_07457_),
    .B(_07480_),
    .X(_07481_));
 sky130_fd_sc_hd__xnor2_1 _15383_ (.A(_07456_),
    .B(_07481_),
    .Y(_07482_));
 sky130_fd_sc_hd__or2_1 _15384_ (.A(net534),
    .B(net487),
    .X(_07483_));
 sky130_fd_sc_hd__inv_2 _15385_ (.A(net539),
    .Y(_07484_));
 sky130_fd_sc_hd__nand2_1 _15386_ (.A(net495),
    .B(net491),
    .Y(_07485_));
 sky130_fd_sc_hd__a2111o_1 _15387_ (.A1(_07438_),
    .A2(_07483_),
    .B1(_07182_),
    .C1(_07484_),
    .D1(_07485_),
    .X(_07486_));
 sky130_fd_sc_hd__a21oi_1 _15388_ (.A1(net541),
    .A2(net482),
    .B1(_07475_),
    .Y(_07487_));
 sky130_fd_sc_hd__a21oi_1 _15389_ (.A1(_07482_),
    .A2(_07486_),
    .B1(_07487_),
    .Y(_07488_));
 sky130_fd_sc_hd__a2bb2o_1 _15390_ (.A1_N(_07482_),
    .A2_N(_07486_),
    .B1(_07476_),
    .B2(_07488_),
    .X(_07489_));
 sky130_fd_sc_hd__xor2_2 _15391_ (.A(_07440_),
    .B(_07441_),
    .X(_07490_));
 sky130_fd_sc_hd__nor2_1 _15392_ (.A(net541),
    .B(_07407_),
    .Y(_07491_));
 sky130_fd_sc_hd__and3b_1 _15393_ (.A_N(net475),
    .B(net472),
    .C(net542),
    .X(_07492_));
 sky130_fd_sc_hd__or2b_2 _15394_ (.A(net472),
    .B_N(net478),
    .X(_07493_));
 sky130_fd_sc_hd__nor3_1 _15395_ (.A(_07182_),
    .B(net539),
    .C(_07493_),
    .Y(_07494_));
 sky130_fd_sc_hd__nor2_1 _15396_ (.A(net472),
    .B(_07407_),
    .Y(_07495_));
 sky130_fd_sc_hd__mux2_1 _15397_ (.A0(_07494_),
    .A1(_07495_),
    .S(_07440_),
    .X(_07496_));
 sky130_fd_sc_hd__and3_1 _15398_ (.A(net541),
    .B(\top0.pid_q.mult0.a[1] ),
    .C(net472),
    .X(_07497_));
 sky130_fd_sc_hd__and3_1 _15399_ (.A(net541),
    .B(_07484_),
    .C(net472),
    .X(_07498_));
 sky130_fd_sc_hd__mux2_1 _15400_ (.A0(_07497_),
    .A1(_07498_),
    .S(_07440_),
    .X(_07499_));
 sky130_fd_sc_hd__or4_1 _15401_ (.A(_07491_),
    .B(_07492_),
    .C(_07496_),
    .D(_07499_),
    .X(_07500_));
 sky130_fd_sc_hd__xnor2_1 _15402_ (.A(_07414_),
    .B(_07500_),
    .Y(_07501_));
 sky130_fd_sc_hd__o21a_1 _15403_ (.A1(_07489_),
    .A2(_07490_),
    .B1(_07501_),
    .X(_07502_));
 sky130_fd_sc_hd__or2b_1 _15404_ (.A(_07456_),
    .B_N(_07457_),
    .X(_07503_));
 sky130_fd_sc_hd__a31o_1 _15405_ (.A1(net537),
    .A2(net486),
    .A3(_07503_),
    .B1(net481),
    .X(_07504_));
 sky130_fd_sc_hd__a21o_1 _15406_ (.A1(net484),
    .A2(_07473_),
    .B1(_07474_),
    .X(_07505_));
 sky130_fd_sc_hd__nand2_1 _15407_ (.A(net481),
    .B(_07459_),
    .Y(_07506_));
 sky130_fd_sc_hd__a22o_1 _15408_ (.A1(net541),
    .A2(_07505_),
    .B1(_07506_),
    .B2(_07478_),
    .X(_07507_));
 sky130_fd_sc_hd__o21a_1 _15409_ (.A1(_07477_),
    .A2(_07504_),
    .B1(_07507_),
    .X(_07508_));
 sky130_fd_sc_hd__a22o_1 _15410_ (.A1(_07501_),
    .A2(_07508_),
    .B1(_07490_),
    .B2(_07489_),
    .X(_07509_));
 sky130_fd_sc_hd__o21a_1 _15411_ (.A1(_07479_),
    .A2(_07502_),
    .B1(_07509_),
    .X(_07510_));
 sky130_fd_sc_hd__or3_1 _15412_ (.A(_07489_),
    .B(_07479_),
    .C(_07490_),
    .X(_07511_));
 sky130_fd_sc_hd__a21o_1 _15413_ (.A1(_07489_),
    .A2(_07490_),
    .B1(_07508_),
    .X(_07512_));
 sky130_fd_sc_hd__a21o_1 _15414_ (.A1(_07511_),
    .A2(_07512_),
    .B1(_07501_),
    .X(_07513_));
 sky130_fd_sc_hd__o221a_1 _15415_ (.A1(_07472_),
    .A2(_07510_),
    .B1(_07460_),
    .B2(_07465_),
    .C1(_07513_),
    .X(_07514_));
 sky130_fd_sc_hd__nor2_1 _15416_ (.A(_07432_),
    .B(_07453_),
    .Y(_07515_));
 sky130_fd_sc_hd__a211o_1 _15417_ (.A1(_07460_),
    .A2(_07465_),
    .B1(_07514_),
    .C1(_07515_),
    .X(_07516_));
 sky130_fd_sc_hd__nor2_1 _15418_ (.A(_07427_),
    .B(_07429_),
    .Y(_07517_));
 sky130_fd_sc_hd__a31o_1 _15419_ (.A1(_07430_),
    .A2(_07454_),
    .A3(_07516_),
    .B1(_07517_),
    .X(_07518_));
 sky130_fd_sc_hd__xor2_1 _15420_ (.A(_07330_),
    .B(_07349_),
    .X(_07519_));
 sky130_fd_sc_hd__xnor2_1 _15421_ (.A(_07332_),
    .B(_07519_),
    .Y(_07520_));
 sky130_fd_sc_hd__nand3_1 _15422_ (.A(_07380_),
    .B(_07381_),
    .C(_07376_),
    .Y(_07521_));
 sky130_fd_sc_hd__a21o_1 _15423_ (.A1(_07380_),
    .A2(_07381_),
    .B1(_07376_),
    .X(_07522_));
 sky130_fd_sc_hd__nand2_1 _15424_ (.A(_07392_),
    .B(_07396_),
    .Y(_07523_));
 sky130_fd_sc_hd__a21o_1 _15425_ (.A1(_07521_),
    .A2(_07522_),
    .B1(_07523_),
    .X(_07524_));
 sky130_fd_sc_hd__nand3_1 _15426_ (.A(_07523_),
    .B(_07521_),
    .C(_07522_),
    .Y(_07525_));
 sky130_fd_sc_hd__o211a_1 _15427_ (.A1(_07520_),
    .A2(_07399_),
    .B1(_07524_),
    .C1(_07525_),
    .X(_07526_));
 sky130_fd_sc_hd__a32o_1 _15428_ (.A1(_07302_),
    .A2(_07350_),
    .A3(_07400_),
    .B1(_07518_),
    .B2(_07526_),
    .X(_07527_));
 sky130_fd_sc_hd__a21o_1 _15429_ (.A1(_07351_),
    .A2(_07352_),
    .B1(_07302_),
    .X(_07528_));
 sky130_fd_sc_hd__and2_1 _15430_ (.A(_07251_),
    .B(_07300_),
    .X(_07529_));
 sky130_fd_sc_hd__or2_1 _15431_ (.A(_07251_),
    .B(_07300_),
    .X(_07530_));
 sky130_fd_sc_hd__o21ai_2 _15432_ (.A1(_07240_),
    .A2(_07529_),
    .B1(_07530_),
    .Y(_07531_));
 sky130_fd_sc_hd__a21o_1 _15433_ (.A1(_07527_),
    .A2(_07528_),
    .B1(_07531_),
    .X(_07532_));
 sky130_fd_sc_hd__nand2_1 _15434_ (.A(_07266_),
    .B(_07280_),
    .Y(_07533_));
 sky130_fd_sc_hd__o21ai_2 _15435_ (.A1(_07266_),
    .A2(_07280_),
    .B1(_07294_),
    .Y(_07534_));
 sky130_fd_sc_hd__and3_1 _15436_ (.A(net494),
    .B(net489),
    .C(net508),
    .X(_07535_));
 sky130_fd_sc_hd__nand2_1 _15437_ (.A(net514),
    .B(net480),
    .Y(_07536_));
 sky130_fd_sc_hd__mux2_1 _15438_ (.A0(net480),
    .A1(_07274_),
    .S(_07366_),
    .X(_07537_));
 sky130_fd_sc_hd__nand2_1 _15439_ (.A(_07276_),
    .B(_07537_),
    .Y(_07538_));
 sky130_fd_sc_hd__o21a_1 _15440_ (.A1(_07274_),
    .A2(_07276_),
    .B1(net484),
    .X(_07539_));
 sky130_fd_sc_hd__and3_1 _15441_ (.A(net489),
    .B(net484),
    .C(net511),
    .X(_07540_));
 sky130_fd_sc_hd__nand2_1 _15442_ (.A(net480),
    .B(_07540_),
    .Y(_07541_));
 sky130_fd_sc_hd__o211a_1 _15443_ (.A1(net480),
    .A2(_07539_),
    .B1(_07541_),
    .C1(net514),
    .X(_07542_));
 sky130_fd_sc_hd__a32o_1 _15444_ (.A1(net511),
    .A2(_07535_),
    .A3(_07536_),
    .B1(_07538_),
    .B2(_07542_),
    .X(_07543_));
 sky130_fd_sc_hd__and3_1 _15445_ (.A(net518),
    .B(net480),
    .C(_07258_),
    .X(_07544_));
 sky130_fd_sc_hd__xor2_1 _15446_ (.A(_07543_),
    .B(_07544_),
    .X(_07545_));
 sky130_fd_sc_hd__nand3_2 _15447_ (.A(_07533_),
    .B(_07534_),
    .C(_07545_),
    .Y(_07546_));
 sky130_fd_sc_hd__a21o_1 _15448_ (.A1(_07533_),
    .A2(_07534_),
    .B1(_07545_),
    .X(_07547_));
 sky130_fd_sc_hd__a21o_1 _15449_ (.A1(_07273_),
    .A2(_07271_),
    .B1(_07278_),
    .X(_07548_));
 sky130_fd_sc_hd__o21a_1 _15450_ (.A1(_07273_),
    .A2(_07271_),
    .B1(_07548_),
    .X(_07549_));
 sky130_fd_sc_hd__nand2_1 _15451_ (.A(net518),
    .B(net475),
    .Y(_07550_));
 sky130_fd_sc_hd__nand2_1 _15452_ (.A(net520),
    .B(net471),
    .Y(_07551_));
 sky130_fd_sc_hd__nand2_1 _15453_ (.A(net522),
    .B(net470),
    .Y(_07552_));
 sky130_fd_sc_hd__xnor2_1 _15454_ (.A(_07551_),
    .B(_07552_),
    .Y(_07553_));
 sky130_fd_sc_hd__xnor2_2 _15455_ (.A(_07550_),
    .B(_07553_),
    .Y(_07554_));
 sky130_fd_sc_hd__o21ai_1 _15456_ (.A1(_07267_),
    .A2(_07268_),
    .B1(_07269_),
    .Y(_07555_));
 sky130_fd_sc_hd__a21bo_1 _15457_ (.A1(_07267_),
    .A2(_07268_),
    .B1_N(_07555_),
    .X(_07556_));
 sky130_fd_sc_hd__nand2_2 _15458_ (.A(net485),
    .B(net511),
    .Y(_07557_));
 sky130_fd_sc_hd__nand2_1 _15459_ (.A(net489),
    .B(net508),
    .Y(_07558_));
 sky130_fd_sc_hd__nand2_1 _15460_ (.A(net493),
    .B(net506),
    .Y(_07559_));
 sky130_fd_sc_hd__xnor2_1 _15461_ (.A(_07558_),
    .B(_07559_),
    .Y(_07560_));
 sky130_fd_sc_hd__xnor2_2 _15462_ (.A(_07557_),
    .B(_07560_),
    .Y(_07561_));
 sky130_fd_sc_hd__xnor2_1 _15463_ (.A(_07556_),
    .B(_07561_),
    .Y(_07562_));
 sky130_fd_sc_hd__xnor2_2 _15464_ (.A(_07554_),
    .B(_07562_),
    .Y(_07563_));
 sky130_fd_sc_hd__xnor2_2 _15465_ (.A(_07549_),
    .B(_07563_),
    .Y(_07564_));
 sky130_fd_sc_hd__nand2_1 _15466_ (.A(net526),
    .B(net464),
    .Y(_07565_));
 sky130_fd_sc_hd__nand2_1 _15467_ (.A(net528),
    .B(net462),
    .Y(_07566_));
 sky130_fd_sc_hd__nand2_1 _15468_ (.A(net531),
    .B(net460),
    .Y(_07567_));
 sky130_fd_sc_hd__xnor2_1 _15469_ (.A(_07566_),
    .B(_07567_),
    .Y(_07568_));
 sky130_fd_sc_hd__xnor2_1 _15470_ (.A(_07565_),
    .B(_07568_),
    .Y(_07569_));
 sky130_fd_sc_hd__nand4_1 _15471_ (.A(net531),
    .B(net528),
    .C(net462),
    .D(net464),
    .Y(_07570_));
 sky130_fd_sc_hd__a22oi_1 _15472_ (.A1(net531),
    .A2(net462),
    .B1(net464),
    .B2(net528),
    .Y(_07571_));
 sky130_fd_sc_hd__a21oi_2 _15473_ (.A1(_07282_),
    .A2(_07570_),
    .B1(_07571_),
    .Y(_07572_));
 sky130_fd_sc_hd__and4_1 _15474_ (.A(net540),
    .B(net538),
    .C(net454),
    .D(net457),
    .X(_07573_));
 sky130_fd_sc_hd__xnor2_1 _15475_ (.A(_07572_),
    .B(_07573_),
    .Y(_07574_));
 sky130_fd_sc_hd__xnor2_1 _15476_ (.A(_07569_),
    .B(_07574_),
    .Y(_07575_));
 sky130_fd_sc_hd__nand2_1 _15477_ (.A(net535),
    .B(net457),
    .Y(_07576_));
 sky130_fd_sc_hd__nand2_1 _15478_ (.A(net538),
    .B(net454),
    .Y(_07577_));
 sky130_fd_sc_hd__nand2_1 _15479_ (.A(net540),
    .B(net451),
    .Y(_07578_));
 sky130_fd_sc_hd__xnor2_1 _15480_ (.A(_07577_),
    .B(_07578_),
    .Y(_07579_));
 sky130_fd_sc_hd__xnor2_1 _15481_ (.A(_07576_),
    .B(_07579_),
    .Y(_07580_));
 sky130_fd_sc_hd__xnor2_1 _15482_ (.A(_07575_),
    .B(_07580_),
    .Y(_07581_));
 sky130_fd_sc_hd__o21a_1 _15483_ (.A1(_07286_),
    .A2(_07291_),
    .B1(_07288_),
    .X(_07582_));
 sky130_fd_sc_hd__a21oi_1 _15484_ (.A1(_07286_),
    .A2(_07291_),
    .B1(_07582_),
    .Y(_07583_));
 sky130_fd_sc_hd__xnor2_1 _15485_ (.A(_07581_),
    .B(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__xnor2_2 _15486_ (.A(_07564_),
    .B(_07584_),
    .Y(_07585_));
 sky130_fd_sc_hd__a21oi_1 _15487_ (.A1(_07546_),
    .A2(_07547_),
    .B1(_07585_),
    .Y(_07586_));
 sky130_fd_sc_hd__and3_1 _15488_ (.A(_07585_),
    .B(_07546_),
    .C(_07547_),
    .X(_07587_));
 sky130_fd_sc_hd__nor2_1 _15489_ (.A(_07194_),
    .B(_07295_),
    .Y(_07588_));
 sky130_fd_sc_hd__nor2_1 _15490_ (.A(_07293_),
    .B(_07588_),
    .Y(_07589_));
 sky130_fd_sc_hd__nor2_1 _15491_ (.A(_07193_),
    .B(_07191_),
    .Y(_07590_));
 sky130_fd_sc_hd__nand2_1 _15492_ (.A(_07293_),
    .B(_07296_),
    .Y(_07591_));
 sky130_fd_sc_hd__mux2_1 _15493_ (.A0(_07590_),
    .A1(_07591_),
    .S(_07281_),
    .X(_07592_));
 sky130_fd_sc_hd__nor2_1 _15494_ (.A(_07589_),
    .B(_07592_),
    .Y(_07593_));
 sky130_fd_sc_hd__o21bai_1 _15495_ (.A1(_07586_),
    .A2(_07587_),
    .B1_N(_07593_),
    .Y(_07594_));
 sky130_fd_sc_hd__or3b_1 _15496_ (.A(_07586_),
    .B(_07587_),
    .C_N(_07593_),
    .X(_07595_));
 sky130_fd_sc_hd__nand2_1 _15497_ (.A(_07594_),
    .B(_07595_),
    .Y(_07596_));
 sky130_fd_sc_hd__nor2_1 _15498_ (.A(net517),
    .B(_07257_),
    .Y(_07597_));
 sky130_fd_sc_hd__nor2_1 _15499_ (.A(_07544_),
    .B(_07597_),
    .Y(_07598_));
 sky130_fd_sc_hd__o22a_2 _15500_ (.A1(net480),
    .A2(_07258_),
    .B1(_07259_),
    .B2(_07598_),
    .X(_07599_));
 sky130_fd_sc_hd__nand2_1 _15501_ (.A(_07298_),
    .B(_07599_),
    .Y(_07600_));
 sky130_fd_sc_hd__inv_2 _15502_ (.A(_07599_),
    .Y(_07601_));
 sky130_fd_sc_hd__o21ba_1 _15503_ (.A1(_07255_),
    .A2(_07601_),
    .B1_N(_07298_),
    .X(_07602_));
 sky130_fd_sc_hd__and2_1 _15504_ (.A(net517),
    .B(_07258_),
    .X(_07603_));
 sky130_fd_sc_hd__or4_2 _15505_ (.A(_07226_),
    .B(_07249_),
    .C(_07597_),
    .D(_07603_),
    .X(_07604_));
 sky130_fd_sc_hd__o22ai_1 _15506_ (.A1(_07255_),
    .A2(_07600_),
    .B1(_07602_),
    .B2(_07604_),
    .Y(_07605_));
 sky130_fd_sc_hd__a21bo_1 _15507_ (.A1(_07253_),
    .A2(_07254_),
    .B1_N(_07604_),
    .X(_07606_));
 sky130_fd_sc_hd__a21o_1 _15508_ (.A1(_07298_),
    .A2(_07599_),
    .B1(_07606_),
    .X(_07607_));
 sky130_fd_sc_hd__or2_1 _15509_ (.A(_07298_),
    .B(_07599_),
    .X(_07608_));
 sky130_fd_sc_hd__a21oi_1 _15510_ (.A1(_07607_),
    .A2(_07608_),
    .B1(_07220_),
    .Y(_07609_));
 sky130_fd_sc_hd__and2_1 _15511_ (.A(_07255_),
    .B(_07601_),
    .X(_07610_));
 sky130_fd_sc_hd__nor2_1 _15512_ (.A(_07255_),
    .B(_07604_),
    .Y(_07611_));
 sky130_fd_sc_hd__mux2_1 _15513_ (.A0(_07610_),
    .A1(_07611_),
    .S(_07298_),
    .X(_07612_));
 sky130_fd_sc_hd__a211o_1 _15514_ (.A1(_07220_),
    .A2(_07605_),
    .B1(_07609_),
    .C1(_07612_),
    .X(_07613_));
 sky130_fd_sc_hd__xnor2_1 _15515_ (.A(_07596_),
    .B(_07613_),
    .Y(_07614_));
 sky130_fd_sc_hd__a31o_1 _15516_ (.A1(_07527_),
    .A2(_07528_),
    .A3(_07531_),
    .B1(_07614_),
    .X(_07615_));
 sky130_fd_sc_hd__nand2_1 _15517_ (.A(_07532_),
    .B(_07615_),
    .Y(_07616_));
 sky130_fd_sc_hd__nand2_2 _15518_ (.A(net486),
    .B(net508),
    .Y(_07617_));
 sky130_fd_sc_hd__nand2_1 _15519_ (.A(net492),
    .B(net506),
    .Y(_07618_));
 sky130_fd_sc_hd__nand2_1 _15520_ (.A(net495),
    .B(net505),
    .Y(_07619_));
 sky130_fd_sc_hd__xnor2_1 _15521_ (.A(_07618_),
    .B(_07619_),
    .Y(_07620_));
 sky130_fd_sc_hd__xnor2_2 _15522_ (.A(_07617_),
    .B(_07620_),
    .Y(_07621_));
 sky130_fd_sc_hd__o21ai_1 _15523_ (.A1(_07550_),
    .A2(_07551_),
    .B1(_07552_),
    .Y(_07622_));
 sky130_fd_sc_hd__a21bo_1 _15524_ (.A1(_07550_),
    .A2(_07551_),
    .B1_N(_07622_),
    .X(_07623_));
 sky130_fd_sc_hd__nand2_2 _15525_ (.A(net478),
    .B(net514),
    .Y(_07624_));
 sky130_fd_sc_hd__nand2_1 _15526_ (.A(net472),
    .B(net518),
    .Y(_07625_));
 sky130_fd_sc_hd__nand2_1 _15527_ (.A(net470),
    .B(net520),
    .Y(_07626_));
 sky130_fd_sc_hd__xnor2_1 _15528_ (.A(_07625_),
    .B(_07626_),
    .Y(_07627_));
 sky130_fd_sc_hd__xnor2_2 _15529_ (.A(_07624_),
    .B(_07627_),
    .Y(_07628_));
 sky130_fd_sc_hd__xnor2_1 _15530_ (.A(_07623_),
    .B(_07628_),
    .Y(_07629_));
 sky130_fd_sc_hd__xnor2_2 _15531_ (.A(_07621_),
    .B(_07629_),
    .Y(_07630_));
 sky130_fd_sc_hd__a21bo_1 _15532_ (.A1(_07572_),
    .A2(_07573_),
    .B1_N(_07569_),
    .X(_07631_));
 sky130_fd_sc_hd__o21ai_1 _15533_ (.A1(_07572_),
    .A2(_07573_),
    .B1(_07631_),
    .Y(_07632_));
 sky130_fd_sc_hd__o21a_1 _15534_ (.A1(_07556_),
    .A2(_07561_),
    .B1(_07554_),
    .X(_07633_));
 sky130_fd_sc_hd__a21o_1 _15535_ (.A1(_07556_),
    .A2(_07561_),
    .B1(_07633_),
    .X(_07634_));
 sky130_fd_sc_hd__xnor2_1 _15536_ (.A(_07632_),
    .B(_07634_),
    .Y(_07635_));
 sky130_fd_sc_hd__xnor2_2 _15537_ (.A(_07630_),
    .B(_07635_),
    .Y(_07636_));
 sky130_fd_sc_hd__nor2_1 _15538_ (.A(_07575_),
    .B(_07580_),
    .Y(_07637_));
 sky130_fd_sc_hd__nand2_2 _15539_ (.A(net465),
    .B(net522),
    .Y(_07638_));
 sky130_fd_sc_hd__nand2_1 _15540_ (.A(net462),
    .B(net526),
    .Y(_07639_));
 sky130_fd_sc_hd__nand2_1 _15541_ (.A(net460),
    .B(net528),
    .Y(_07640_));
 sky130_fd_sc_hd__xnor2_1 _15542_ (.A(_07639_),
    .B(_07640_),
    .Y(_07641_));
 sky130_fd_sc_hd__xnor2_2 _15543_ (.A(_07638_),
    .B(_07641_),
    .Y(_07642_));
 sky130_fd_sc_hd__o21a_1 _15544_ (.A1(_07576_),
    .A2(_07577_),
    .B1(_07578_),
    .X(_07643_));
 sky130_fd_sc_hd__a21o_1 _15545_ (.A1(_07576_),
    .A2(_07577_),
    .B1(_07643_),
    .X(_07644_));
 sky130_fd_sc_hd__o21a_1 _15546_ (.A1(_07565_),
    .A2(_07566_),
    .B1(_07567_),
    .X(_07645_));
 sky130_fd_sc_hd__a21o_1 _15547_ (.A1(_07565_),
    .A2(_07566_),
    .B1(_07645_),
    .X(_07646_));
 sky130_fd_sc_hd__xnor2_1 _15548_ (.A(_07644_),
    .B(_07646_),
    .Y(_07647_));
 sky130_fd_sc_hd__xnor2_1 _15549_ (.A(_07642_),
    .B(_07647_),
    .Y(_07648_));
 sky130_fd_sc_hd__nand2_1 _15550_ (.A(net448),
    .B(net540),
    .Y(_07649_));
 sky130_fd_sc_hd__nand2_1 _15551_ (.A(net457),
    .B(net531),
    .Y(_07650_));
 sky130_fd_sc_hd__nand2_1 _15552_ (.A(net454),
    .B(net536),
    .Y(_07651_));
 sky130_fd_sc_hd__nand2_1 _15553_ (.A(net451),
    .B(net538),
    .Y(_07652_));
 sky130_fd_sc_hd__xnor2_1 _15554_ (.A(_07651_),
    .B(_07652_),
    .Y(_07653_));
 sky130_fd_sc_hd__xnor2_1 _15555_ (.A(_07650_),
    .B(_07653_),
    .Y(_07654_));
 sky130_fd_sc_hd__xnor2_1 _15556_ (.A(_07649_),
    .B(_07654_),
    .Y(_07655_));
 sky130_fd_sc_hd__nor2_1 _15557_ (.A(_07648_),
    .B(_07655_),
    .Y(_07656_));
 sky130_fd_sc_hd__and2_1 _15558_ (.A(_07648_),
    .B(_07655_),
    .X(_07657_));
 sky130_fd_sc_hd__or2_1 _15559_ (.A(_07656_),
    .B(_07657_),
    .X(_07658_));
 sky130_fd_sc_hd__xor2_1 _15560_ (.A(_07637_),
    .B(_07658_),
    .X(_07659_));
 sky130_fd_sc_hd__xnor2_2 _15561_ (.A(_07636_),
    .B(_07659_),
    .Y(_07660_));
 sky130_fd_sc_hd__nand2_1 _15562_ (.A(_07288_),
    .B(_07286_),
    .Y(_07661_));
 sky130_fd_sc_hd__a21o_1 _15563_ (.A1(_07563_),
    .A2(_07661_),
    .B1(_07549_),
    .X(_07662_));
 sky130_fd_sc_hd__o21a_2 _15564_ (.A1(_07563_),
    .A2(_07661_),
    .B1(_07662_),
    .X(_07663_));
 sky130_fd_sc_hd__o21a_1 _15565_ (.A1(_07557_),
    .A2(_07558_),
    .B1(_07559_),
    .X(_07664_));
 sky130_fd_sc_hd__a21oi_1 _15566_ (.A1(_07557_),
    .A2(_07558_),
    .B1(_07664_),
    .Y(_07665_));
 sky130_fd_sc_hd__o21a_1 _15567_ (.A1(net484),
    .A2(_07274_),
    .B1(_07276_),
    .X(_07666_));
 sky130_fd_sc_hd__o21ai_2 _15568_ (.A1(_07540_),
    .A2(_07666_),
    .B1(net514),
    .Y(_07667_));
 sky130_fd_sc_hd__xnor2_1 _15569_ (.A(net511),
    .B(_07667_),
    .Y(_07668_));
 sky130_fd_sc_hd__nand2_1 _15570_ (.A(net480),
    .B(_07668_),
    .Y(_07669_));
 sky130_fd_sc_hd__xnor2_1 _15571_ (.A(_07665_),
    .B(_07669_),
    .Y(_07670_));
 sky130_fd_sc_hd__xnor2_2 _15572_ (.A(_07663_),
    .B(_07670_),
    .Y(_07671_));
 sky130_fd_sc_hd__o21ai_1 _15573_ (.A1(_07288_),
    .A2(_07286_),
    .B1(_07291_),
    .Y(_07672_));
 sky130_fd_sc_hd__o21ai_1 _15574_ (.A1(_07564_),
    .A2(_07672_),
    .B1(_07581_),
    .Y(_07673_));
 sky130_fd_sc_hd__nand2_1 _15575_ (.A(_07564_),
    .B(_07583_),
    .Y(_07674_));
 sky130_fd_sc_hd__o211a_1 _15576_ (.A1(_07564_),
    .A2(_07661_),
    .B1(_07673_),
    .C1(_07674_),
    .X(_07675_));
 sky130_fd_sc_hd__xnor2_1 _15577_ (.A(_07671_),
    .B(_07675_),
    .Y(_07676_));
 sky130_fd_sc_hd__xnor2_1 _15578_ (.A(_07660_),
    .B(_07676_),
    .Y(_07677_));
 sky130_fd_sc_hd__inv_2 _15579_ (.A(_07296_),
    .Y(_07678_));
 sky130_fd_sc_hd__mux2_1 _15580_ (.A0(_07590_),
    .A1(_07678_),
    .S(_07281_),
    .X(_07679_));
 sky130_fd_sc_hd__inv_2 _15581_ (.A(_07281_),
    .Y(_07680_));
 sky130_fd_sc_hd__a21oi_1 _15582_ (.A1(_07680_),
    .A2(_07588_),
    .B1(_07293_),
    .Y(_07681_));
 sky130_fd_sc_hd__nand2_1 _15583_ (.A(_07546_),
    .B(_07547_),
    .Y(_07682_));
 sky130_fd_sc_hd__a2bb2oi_1 _15584_ (.A1_N(_07589_),
    .A2_N(_07592_),
    .B1(_07546_),
    .B2(_07547_),
    .Y(_07683_));
 sky130_fd_sc_hd__o32a_1 _15585_ (.A1(_07679_),
    .A2(_07681_),
    .A3(_07682_),
    .B1(_07683_),
    .B2(_07585_),
    .X(_07684_));
 sky130_fd_sc_hd__o211a_1 _15586_ (.A1(_07543_),
    .A2(_07544_),
    .B1(_07533_),
    .C1(_07534_),
    .X(_07685_));
 sky130_fd_sc_hd__a21o_1 _15587_ (.A1(_07543_),
    .A2(_07544_),
    .B1(_07685_),
    .X(_07686_));
 sky130_fd_sc_hd__xor2_1 _15588_ (.A(_07684_),
    .B(_07686_),
    .X(_07687_));
 sky130_fd_sc_hd__xor2_1 _15589_ (.A(_07677_),
    .B(_07687_),
    .X(_07688_));
 sky130_fd_sc_hd__o211a_1 _15590_ (.A1(_07255_),
    .A2(_07604_),
    .B1(_07595_),
    .C1(_07594_),
    .X(_07689_));
 sky130_fd_sc_hd__a2bb2o_1 _15591_ (.A1_N(_07610_),
    .A2_N(_07689_),
    .B1(_07220_),
    .B2(_07298_),
    .X(_07690_));
 sky130_fd_sc_hd__or2_1 _15592_ (.A(_07220_),
    .B(_07298_),
    .X(_07691_));
 sky130_fd_sc_hd__a22o_1 _15593_ (.A1(_07599_),
    .A2(_07606_),
    .B1(_07691_),
    .B2(_07596_),
    .X(_07692_));
 sky130_fd_sc_hd__or2_1 _15594_ (.A(_07596_),
    .B(_07691_),
    .X(_07693_));
 sky130_fd_sc_hd__and4_2 _15595_ (.A(_07688_),
    .B(_07690_),
    .C(_07692_),
    .D(_07693_),
    .X(_07694_));
 sky130_fd_sc_hd__a31oi_2 _15596_ (.A1(_07690_),
    .A2(_07692_),
    .A3(_07693_),
    .B1(_07688_),
    .Y(_07695_));
 sky130_fd_sc_hd__or2_1 _15597_ (.A(_07694_),
    .B(_07695_),
    .X(_07696_));
 sky130_fd_sc_hd__xnor2_2 _15598_ (.A(_07616_),
    .B(_07696_),
    .Y(_07697_));
 sky130_fd_sc_hd__or2_2 _15599_ (.A(net553),
    .B(net543),
    .X(_07698_));
 sky130_fd_sc_hd__nor3_1 _15600_ (.A(\top0.pid_q.state[0] ),
    .B(net546),
    .C(_07698_),
    .Y(_07699_));
 sky130_fd_sc_hd__clkbuf_4 _15601_ (.A(_07699_),
    .X(_07700_));
 sky130_fd_sc_hd__nand2_1 _15602_ (.A(net548),
    .B(_07700_),
    .Y(_07701_));
 sky130_fd_sc_hd__nor2_1 _15603_ (.A(_07697_),
    .B(_07701_),
    .Y(_07702_));
 sky130_fd_sc_hd__or3_1 _15604_ (.A(\top0.pid_q.state[0] ),
    .B(net546),
    .C(_07698_),
    .X(_07703_));
 sky130_fd_sc_hd__buf_2 _15605_ (.A(_07703_),
    .X(_07704_));
 sky130_fd_sc_hd__clkbuf_4 _15606_ (.A(_07704_),
    .X(_07705_));
 sky130_fd_sc_hd__inv_2 _15607_ (.A(\top0.pid_q.curr_int[0] ),
    .Y(_07706_));
 sky130_fd_sc_hd__nor2_1 _15608_ (.A(_07706_),
    .B(_07704_),
    .Y(_07707_));
 sky130_fd_sc_hd__mux2_1 _15609_ (.A0(_07707_),
    .A1(_07706_),
    .S(\top0.pid_q.out[0] ),
    .X(_07708_));
 sky130_fd_sc_hd__a22o_1 _15610_ (.A1(\top0.pid_q.out[0] ),
    .A2(_07705_),
    .B1(_07708_),
    .B2(net544),
    .X(_07709_));
 sky130_fd_sc_hd__buf_4 _15611_ (.A(net1019),
    .X(_07710_));
 sky130_fd_sc_hd__o21a_1 _15612_ (.A1(_07702_),
    .A2(_07709_),
    .B1(_07710_),
    .X(_00133_));
 sky130_fd_sc_hd__inv_2 _15613_ (.A(_07694_),
    .Y(_07711_));
 sky130_fd_sc_hd__a21o_1 _15614_ (.A1(_07616_),
    .A2(_07711_),
    .B1(_07695_),
    .X(_07712_));
 sky130_fd_sc_hd__nor2_1 _15615_ (.A(_07585_),
    .B(_07683_),
    .Y(_07713_));
 sky130_fd_sc_hd__a31o_1 _15616_ (.A1(_07593_),
    .A2(_07546_),
    .A3(_07547_),
    .B1(_07713_),
    .X(_07714_));
 sky130_fd_sc_hd__o21ba_1 _15617_ (.A1(_07714_),
    .A2(_07686_),
    .B1_N(_07677_),
    .X(_07715_));
 sky130_fd_sc_hd__a21oi_1 _15618_ (.A1(_07714_),
    .A2(_07686_),
    .B1(_07715_),
    .Y(_07716_));
 sky130_fd_sc_hd__o21ba_1 _15619_ (.A1(_07636_),
    .A2(_07658_),
    .B1_N(_07637_),
    .X(_07717_));
 sky130_fd_sc_hd__a21o_1 _15620_ (.A1(_07636_),
    .A2(_07658_),
    .B1(_07717_),
    .X(_07718_));
 sky130_fd_sc_hd__nand2_2 _15621_ (.A(net477),
    .B(net512),
    .Y(_07719_));
 sky130_fd_sc_hd__nand2_1 _15622_ (.A(net474),
    .B(net514),
    .Y(_07720_));
 sky130_fd_sc_hd__nand2_1 _15623_ (.A(net469),
    .B(net518),
    .Y(_07721_));
 sky130_fd_sc_hd__xnor2_1 _15624_ (.A(_07720_),
    .B(_07721_),
    .Y(_07722_));
 sky130_fd_sc_hd__xnor2_2 _15625_ (.A(_07719_),
    .B(_07722_),
    .Y(_07723_));
 sky130_fd_sc_hd__o21ai_1 _15626_ (.A1(_07624_),
    .A2(_07625_),
    .B1(_07626_),
    .Y(_07724_));
 sky130_fd_sc_hd__a21bo_1 _15627_ (.A1(_07624_),
    .A2(_07625_),
    .B1_N(_07724_),
    .X(_07725_));
 sky130_fd_sc_hd__and2_1 _15628_ (.A(net496),
    .B(net502),
    .X(_07726_));
 sky130_fd_sc_hd__nand2_1 _15629_ (.A(net506),
    .B(net488),
    .Y(_07727_));
 sky130_fd_sc_hd__nand2_1 _15630_ (.A(net505),
    .B(net492),
    .Y(_07728_));
 sky130_fd_sc_hd__xor2_1 _15631_ (.A(_07727_),
    .B(_07728_),
    .X(_07729_));
 sky130_fd_sc_hd__xnor2_2 _15632_ (.A(_07726_),
    .B(_07729_),
    .Y(_07730_));
 sky130_fd_sc_hd__xnor2_1 _15633_ (.A(_07725_),
    .B(_07730_),
    .Y(_07731_));
 sky130_fd_sc_hd__xnor2_2 _15634_ (.A(_07723_),
    .B(_07731_),
    .Y(_07732_));
 sky130_fd_sc_hd__o21a_1 _15635_ (.A1(_07642_),
    .A2(_07646_),
    .B1(_07644_),
    .X(_07733_));
 sky130_fd_sc_hd__a21o_1 _15636_ (.A1(_07642_),
    .A2(_07646_),
    .B1(_07733_),
    .X(_07734_));
 sky130_fd_sc_hd__o21a_1 _15637_ (.A1(_07623_),
    .A2(_07628_),
    .B1(_07621_),
    .X(_07735_));
 sky130_fd_sc_hd__a21o_1 _15638_ (.A1(_07623_),
    .A2(_07628_),
    .B1(_07735_),
    .X(_07736_));
 sky130_fd_sc_hd__xnor2_1 _15639_ (.A(_07734_),
    .B(_07736_),
    .Y(_07737_));
 sky130_fd_sc_hd__xnor2_2 _15640_ (.A(_07732_),
    .B(_07737_),
    .Y(_07738_));
 sky130_fd_sc_hd__nand2_2 _15641_ (.A(net465),
    .B(net520),
    .Y(_07739_));
 sky130_fd_sc_hd__nand2_1 _15642_ (.A(net462),
    .B(net522),
    .Y(_07740_));
 sky130_fd_sc_hd__nand2_1 _15643_ (.A(net460),
    .B(net525),
    .Y(_07741_));
 sky130_fd_sc_hd__xnor2_1 _15644_ (.A(_07740_),
    .B(_07741_),
    .Y(_07742_));
 sky130_fd_sc_hd__xnor2_2 _15645_ (.A(_07739_),
    .B(_07742_),
    .Y(_07743_));
 sky130_fd_sc_hd__o21a_1 _15646_ (.A1(_07650_),
    .A2(_07651_),
    .B1(_07652_),
    .X(_07744_));
 sky130_fd_sc_hd__a21oi_2 _15647_ (.A1(_07650_),
    .A2(_07651_),
    .B1(_07744_),
    .Y(_07745_));
 sky130_fd_sc_hd__o21a_1 _15648_ (.A1(_07638_),
    .A2(_07639_),
    .B1(_07640_),
    .X(_07746_));
 sky130_fd_sc_hd__a21oi_2 _15649_ (.A1(_07638_),
    .A2(_07639_),
    .B1(_07746_),
    .Y(_07747_));
 sky130_fd_sc_hd__xor2_1 _15650_ (.A(_07745_),
    .B(_07747_),
    .X(_07748_));
 sky130_fd_sc_hd__xnor2_2 _15651_ (.A(_07743_),
    .B(_07748_),
    .Y(_07749_));
 sky130_fd_sc_hd__nor2_1 _15652_ (.A(_07649_),
    .B(_07654_),
    .Y(_07750_));
 sky130_fd_sc_hd__nand2_1 _15653_ (.A(net540),
    .B(net446),
    .Y(_07751_));
 sky130_fd_sc_hd__nand2_1 _15654_ (.A(net448),
    .B(net538),
    .Y(_07752_));
 sky130_fd_sc_hd__xor2_1 _15655_ (.A(_07751_),
    .B(_07752_),
    .X(_07753_));
 sky130_fd_sc_hd__nand2_1 _15656_ (.A(net457),
    .B(net529),
    .Y(_07754_));
 sky130_fd_sc_hd__nand2_1 _15657_ (.A(net454),
    .B(net532),
    .Y(_07755_));
 sky130_fd_sc_hd__nand2_1 _15658_ (.A(net451),
    .B(net536),
    .Y(_07756_));
 sky130_fd_sc_hd__xor2_1 _15659_ (.A(_07755_),
    .B(_07756_),
    .X(_07757_));
 sky130_fd_sc_hd__xnor2_1 _15660_ (.A(_07754_),
    .B(_07757_),
    .Y(_07758_));
 sky130_fd_sc_hd__xor2_1 _15661_ (.A(_07753_),
    .B(_07758_),
    .X(_07759_));
 sky130_fd_sc_hd__xor2_1 _15662_ (.A(_07750_),
    .B(_07759_),
    .X(_07760_));
 sky130_fd_sc_hd__xnor2_2 _15663_ (.A(_07749_),
    .B(_07760_),
    .Y(_07761_));
 sky130_fd_sc_hd__xor2_1 _15664_ (.A(_07656_),
    .B(_07761_),
    .X(_07762_));
 sky130_fd_sc_hd__xnor2_1 _15665_ (.A(_07738_),
    .B(_07762_),
    .Y(_07763_));
 sky130_fd_sc_hd__a21o_1 _15666_ (.A1(_07630_),
    .A2(_07634_),
    .B1(_07632_),
    .X(_07764_));
 sky130_fd_sc_hd__o21a_1 _15667_ (.A1(_07630_),
    .A2(_07634_),
    .B1(_07764_),
    .X(_07765_));
 sky130_fd_sc_hd__o21a_1 _15668_ (.A1(_07617_),
    .A2(_07618_),
    .B1(_07619_),
    .X(_07766_));
 sky130_fd_sc_hd__a21o_1 _15669_ (.A1(_07617_),
    .A2(_07618_),
    .B1(_07766_),
    .X(_07767_));
 sky130_fd_sc_hd__a21oi_1 _15670_ (.A1(_07366_),
    .A2(_07558_),
    .B1(_07559_),
    .Y(_07768_));
 sky130_fd_sc_hd__a31o_1 _15671_ (.A1(net490),
    .A2(net486),
    .A3(net508),
    .B1(_07768_),
    .X(_07769_));
 sky130_fd_sc_hd__nand2_1 _15672_ (.A(net511),
    .B(_07769_),
    .Y(_07770_));
 sky130_fd_sc_hd__xnor2_1 _15673_ (.A(net508),
    .B(_07770_),
    .Y(_07771_));
 sky130_fd_sc_hd__nand2_1 _15674_ (.A(net481),
    .B(_07771_),
    .Y(_07772_));
 sky130_fd_sc_hd__xnor2_1 _15675_ (.A(_07767_),
    .B(_07772_),
    .Y(_07773_));
 sky130_fd_sc_hd__xnor2_1 _15676_ (.A(_07765_),
    .B(_07773_),
    .Y(_07774_));
 sky130_fd_sc_hd__nor2_1 _15677_ (.A(_07763_),
    .B(_07774_),
    .Y(_07775_));
 sky130_fd_sc_hd__and2_1 _15678_ (.A(_07763_),
    .B(_07774_),
    .X(_07776_));
 sky130_fd_sc_hd__nor2_1 _15679_ (.A(_07775_),
    .B(_07776_),
    .Y(_07777_));
 sky130_fd_sc_hd__xnor2_1 _15680_ (.A(_07718_),
    .B(_07777_),
    .Y(_07778_));
 sky130_fd_sc_hd__inv_2 _15681_ (.A(_07665_),
    .Y(_07779_));
 sky130_fd_sc_hd__nand2_1 _15682_ (.A(_07663_),
    .B(_07667_),
    .Y(_07780_));
 sky130_fd_sc_hd__inv_2 _15683_ (.A(net506),
    .Y(_07781_));
 sky130_fd_sc_hd__or3b_1 _15684_ (.A(_07781_),
    .B(net511),
    .C_N(_07535_),
    .X(_07782_));
 sky130_fd_sc_hd__a21oi_1 _15685_ (.A1(_07663_),
    .A2(_07782_),
    .B1(_07667_),
    .Y(_07783_));
 sky130_fd_sc_hd__a31o_1 _15686_ (.A1(net511),
    .A2(_07779_),
    .A3(_07780_),
    .B1(_07783_),
    .X(_07784_));
 sky130_fd_sc_hd__a211o_1 _15687_ (.A1(net511),
    .A2(net480),
    .B1(_07663_),
    .C1(_07779_),
    .X(_07785_));
 sky130_fd_sc_hd__a21bo_1 _15688_ (.A1(net481),
    .A2(_07784_),
    .B1_N(_07785_),
    .X(_07786_));
 sky130_fd_sc_hd__nand2_1 _15689_ (.A(_07671_),
    .B(_07675_),
    .Y(_07787_));
 sky130_fd_sc_hd__nor2_1 _15690_ (.A(_07671_),
    .B(_07675_),
    .Y(_07788_));
 sky130_fd_sc_hd__a21oi_2 _15691_ (.A1(_07660_),
    .A2(_07787_),
    .B1(_07788_),
    .Y(_07789_));
 sky130_fd_sc_hd__xor2_1 _15692_ (.A(_07786_),
    .B(_07789_),
    .X(_07790_));
 sky130_fd_sc_hd__xnor2_1 _15693_ (.A(_07778_),
    .B(_07790_),
    .Y(_07791_));
 sky130_fd_sc_hd__nor2_1 _15694_ (.A(_07716_),
    .B(_07791_),
    .Y(_07792_));
 sky130_fd_sc_hd__nand2_1 _15695_ (.A(_07716_),
    .B(_07791_),
    .Y(_07793_));
 sky130_fd_sc_hd__and2b_1 _15696_ (.A_N(_07792_),
    .B(_07793_),
    .X(_07794_));
 sky130_fd_sc_hd__xnor2_2 _15697_ (.A(_07712_),
    .B(_07794_),
    .Y(_07795_));
 sky130_fd_sc_hd__nand2_1 _15698_ (.A(\top0.pid_q.out[0] ),
    .B(\top0.pid_q.curr_int[0] ),
    .Y(_07796_));
 sky130_fd_sc_hd__xor2_1 _15699_ (.A(\top0.pid_q.out[1] ),
    .B(\top0.pid_q.curr_int[1] ),
    .X(_07797_));
 sky130_fd_sc_hd__xnor2_1 _15700_ (.A(_07796_),
    .B(_07797_),
    .Y(_07798_));
 sky130_fd_sc_hd__a221o_1 _15701_ (.A1(net549),
    .A2(_07795_),
    .B1(_07798_),
    .B2(net544),
    .C1(_07705_),
    .X(_07799_));
 sky130_fd_sc_hd__o211a_1 _15702_ (.A1(\top0.pid_q.out[1] ),
    .A2(_07700_),
    .B1(_07799_),
    .C1(_07710_),
    .X(_00134_));
 sky130_fd_sc_hd__clkbuf_4 _15703_ (.A(_05443_),
    .X(_07800_));
 sky130_fd_sc_hd__nor2_1 _15704_ (.A(\top0.pid_q.out[2] ),
    .B(_07703_),
    .Y(_07801_));
 sky130_fd_sc_hd__a22o_1 _15705_ (.A1(\top0.pid_q.out[0] ),
    .A2(\top0.pid_q.curr_int[0] ),
    .B1(\top0.pid_q.curr_int[1] ),
    .B2(\top0.pid_q.out[1] ),
    .X(_07802_));
 sky130_fd_sc_hd__or2_1 _15706_ (.A(\top0.pid_q.out[1] ),
    .B(\top0.pid_q.curr_int[1] ),
    .X(_07803_));
 sky130_fd_sc_hd__nand2_1 _15707_ (.A(_07802_),
    .B(_07803_),
    .Y(_07804_));
 sky130_fd_sc_hd__xnor2_1 _15708_ (.A(\top0.pid_q.curr_int[2] ),
    .B(_07804_),
    .Y(_07805_));
 sky130_fd_sc_hd__mux2_1 _15709_ (.A0(\top0.pid_q.out[2] ),
    .A1(_07801_),
    .S(_07805_),
    .X(_07806_));
 sky130_fd_sc_hd__a221o_1 _15710_ (.A1(_07527_),
    .A2(_07528_),
    .B1(_07531_),
    .B2(_07614_),
    .C1(_07694_),
    .X(_07807_));
 sky130_fd_sc_hd__nor2_1 _15711_ (.A(_07531_),
    .B(_07614_),
    .Y(_07808_));
 sky130_fd_sc_hd__o21bai_1 _15712_ (.A1(_07695_),
    .A2(_07808_),
    .B1_N(_07694_),
    .Y(_07809_));
 sky130_fd_sc_hd__a31o_2 _15713_ (.A1(_07793_),
    .A2(_07807_),
    .A3(_07809_),
    .B1(_07792_),
    .X(_07810_));
 sky130_fd_sc_hd__o21a_1 _15714_ (.A1(_07786_),
    .A2(_07789_),
    .B1(_07778_),
    .X(_07811_));
 sky130_fd_sc_hd__a21oi_1 _15715_ (.A1(_07786_),
    .A2(_07789_),
    .B1(_07811_),
    .Y(_07812_));
 sky130_fd_sc_hd__nand2_2 _15716_ (.A(net474),
    .B(net512),
    .Y(_07813_));
 sky130_fd_sc_hd__nand2_1 _15717_ (.A(net469),
    .B(net515),
    .Y(_07814_));
 sky130_fd_sc_hd__nand2_1 _15718_ (.A(net477),
    .B(net509),
    .Y(_07815_));
 sky130_fd_sc_hd__xnor2_1 _15719_ (.A(_07814_),
    .B(_07815_),
    .Y(_07816_));
 sky130_fd_sc_hd__xnor2_2 _15720_ (.A(_07813_),
    .B(_07816_),
    .Y(_07817_));
 sky130_fd_sc_hd__o21ai_1 _15721_ (.A1(_07719_),
    .A2(_07720_),
    .B1(_07721_),
    .Y(_07818_));
 sky130_fd_sc_hd__a21bo_1 _15722_ (.A1(_07719_),
    .A2(_07720_),
    .B1_N(_07818_),
    .X(_07819_));
 sky130_fd_sc_hd__nand2_1 _15723_ (.A(net496),
    .B(net499),
    .Y(_07820_));
 sky130_fd_sc_hd__nand2_1 _15724_ (.A(net505),
    .B(net488),
    .Y(_07821_));
 sky130_fd_sc_hd__nand2_1 _15725_ (.A(net492),
    .B(net502),
    .Y(_07822_));
 sky130_fd_sc_hd__xnor2_1 _15726_ (.A(_07821_),
    .B(_07822_),
    .Y(_07823_));
 sky130_fd_sc_hd__xnor2_2 _15727_ (.A(_07820_),
    .B(_07823_),
    .Y(_07824_));
 sky130_fd_sc_hd__xnor2_1 _15728_ (.A(_07819_),
    .B(_07824_),
    .Y(_07825_));
 sky130_fd_sc_hd__xnor2_2 _15729_ (.A(_07817_),
    .B(_07825_),
    .Y(_07826_));
 sky130_fd_sc_hd__a21bo_1 _15730_ (.A1(_07745_),
    .A2(_07747_),
    .B1_N(_07743_),
    .X(_07827_));
 sky130_fd_sc_hd__o21ai_2 _15731_ (.A1(_07745_),
    .A2(_07747_),
    .B1(_07827_),
    .Y(_07828_));
 sky130_fd_sc_hd__o21a_1 _15732_ (.A1(_07725_),
    .A2(_07730_),
    .B1(_07723_),
    .X(_07829_));
 sky130_fd_sc_hd__a21o_1 _15733_ (.A1(_07725_),
    .A2(_07730_),
    .B1(_07829_),
    .X(_07830_));
 sky130_fd_sc_hd__xnor2_1 _15734_ (.A(_07828_),
    .B(_07830_),
    .Y(_07831_));
 sky130_fd_sc_hd__xnor2_2 _15735_ (.A(_07826_),
    .B(_07831_),
    .Y(_07832_));
 sky130_fd_sc_hd__nand2_1 _15736_ (.A(net457),
    .B(net526),
    .Y(_07833_));
 sky130_fd_sc_hd__nand2_1 _15737_ (.A(net451),
    .B(net532),
    .Y(_07834_));
 sky130_fd_sc_hd__nand2_1 _15738_ (.A(net454),
    .B(net528),
    .Y(_07835_));
 sky130_fd_sc_hd__xnor2_1 _15739_ (.A(_07834_),
    .B(_07835_),
    .Y(_07836_));
 sky130_fd_sc_hd__xnor2_1 _15740_ (.A(_07833_),
    .B(_07836_),
    .Y(_07837_));
 sky130_fd_sc_hd__nand2_2 _15741_ (.A(net538),
    .B(net446),
    .Y(_07838_));
 sky130_fd_sc_hd__and2_1 _15742_ (.A(net448),
    .B(net536),
    .X(_07839_));
 sky130_fd_sc_hd__o21ba_1 _15743_ (.A1(net448),
    .A2(_07838_),
    .B1_N(_07839_),
    .X(_07840_));
 sky130_fd_sc_hd__xor2_1 _15744_ (.A(net443),
    .B(_07838_),
    .X(_07841_));
 sky130_fd_sc_hd__nand2_1 _15745_ (.A(_07182_),
    .B(net443),
    .Y(_07842_));
 sky130_fd_sc_hd__mux2_1 _15746_ (.A0(net443),
    .A1(_07842_),
    .S(_07838_),
    .X(_07843_));
 sky130_fd_sc_hd__o32a_1 _15747_ (.A1(net541),
    .A2(net536),
    .A3(_07841_),
    .B1(_07843_),
    .B2(net448),
    .X(_07844_));
 sky130_fd_sc_hd__nand2_1 _15748_ (.A(_07839_),
    .B(_07841_),
    .Y(_07845_));
 sky130_fd_sc_hd__o211a_1 _15749_ (.A1(_07182_),
    .A2(_07840_),
    .B1(_07844_),
    .C1(_07845_),
    .X(_07846_));
 sky130_fd_sc_hd__xnor2_1 _15750_ (.A(_07837_),
    .B(_07846_),
    .Y(_07847_));
 sky130_fd_sc_hd__nand2_1 _15751_ (.A(_07753_),
    .B(_07758_),
    .Y(_07848_));
 sky130_fd_sc_hd__nand2_1 _15752_ (.A(net465),
    .B(net518),
    .Y(_07849_));
 sky130_fd_sc_hd__nand2_1 _15753_ (.A(net460),
    .B(net523),
    .Y(_07850_));
 sky130_fd_sc_hd__nand2_1 _15754_ (.A(net461),
    .B(net521),
    .Y(_07851_));
 sky130_fd_sc_hd__xnor2_1 _15755_ (.A(_07850_),
    .B(_07851_),
    .Y(_07852_));
 sky130_fd_sc_hd__xnor2_1 _15756_ (.A(_07849_),
    .B(_07852_),
    .Y(_07853_));
 sky130_fd_sc_hd__o21a_1 _15757_ (.A1(_07754_),
    .A2(_07755_),
    .B1(_07756_),
    .X(_07854_));
 sky130_fd_sc_hd__a21oi_2 _15758_ (.A1(_07754_),
    .A2(_07755_),
    .B1(_07854_),
    .Y(_07855_));
 sky130_fd_sc_hd__o21a_1 _15759_ (.A1(_07739_),
    .A2(_07740_),
    .B1(_07741_),
    .X(_07856_));
 sky130_fd_sc_hd__a21oi_2 _15760_ (.A1(_07739_),
    .A2(_07740_),
    .B1(_07856_),
    .Y(_07857_));
 sky130_fd_sc_hd__xnor2_1 _15761_ (.A(_07855_),
    .B(_07857_),
    .Y(_07858_));
 sky130_fd_sc_hd__xnor2_1 _15762_ (.A(_07853_),
    .B(_07858_),
    .Y(_07859_));
 sky130_fd_sc_hd__xor2_1 _15763_ (.A(_07848_),
    .B(_07859_),
    .X(_07860_));
 sky130_fd_sc_hd__xnor2_1 _15764_ (.A(_07847_),
    .B(_07860_),
    .Y(_07861_));
 sky130_fd_sc_hd__a21o_1 _15765_ (.A1(_07749_),
    .A2(_07750_),
    .B1(_07759_),
    .X(_07862_));
 sky130_fd_sc_hd__o21a_1 _15766_ (.A1(_07749_),
    .A2(_07750_),
    .B1(_07862_),
    .X(_07863_));
 sky130_fd_sc_hd__nor2_1 _15767_ (.A(_07861_),
    .B(_07863_),
    .Y(_07864_));
 sky130_fd_sc_hd__and2_1 _15768_ (.A(_07861_),
    .B(_07863_),
    .X(_07865_));
 sky130_fd_sc_hd__nor2_1 _15769_ (.A(_07864_),
    .B(_07865_),
    .Y(_07866_));
 sky130_fd_sc_hd__xor2_2 _15770_ (.A(_07832_),
    .B(_07866_),
    .X(_07867_));
 sky130_fd_sc_hd__o21ba_1 _15771_ (.A1(_07738_),
    .A2(_07761_),
    .B1_N(_07656_),
    .X(_07868_));
 sky130_fd_sc_hd__a21o_1 _15772_ (.A1(_07738_),
    .A2(_07761_),
    .B1(_07868_),
    .X(_07869_));
 sky130_fd_sc_hd__a21o_1 _15773_ (.A1(_07732_),
    .A2(_07736_),
    .B1(_07734_),
    .X(_07870_));
 sky130_fd_sc_hd__o21a_1 _15774_ (.A1(_07732_),
    .A2(_07736_),
    .B1(_07870_),
    .X(_07871_));
 sky130_fd_sc_hd__o21ba_1 _15775_ (.A1(_07727_),
    .A2(_07728_),
    .B1_N(_07726_),
    .X(_07872_));
 sky130_fd_sc_hd__a21oi_2 _15776_ (.A1(_07727_),
    .A2(_07728_),
    .B1(_07872_),
    .Y(_07873_));
 sky130_fd_sc_hd__nand2_1 _15777_ (.A(net506),
    .B(net483),
    .Y(_07874_));
 sky130_fd_sc_hd__xor2_1 _15778_ (.A(net443),
    .B(_07874_),
    .X(_07875_));
 sky130_fd_sc_hd__xnor2_2 _15779_ (.A(_07873_),
    .B(_07875_),
    .Y(_07876_));
 sky130_fd_sc_hd__inv_2 _15780_ (.A(_07767_),
    .Y(_07877_));
 sky130_fd_sc_hd__and3_1 _15781_ (.A(net508),
    .B(net481),
    .C(_07877_),
    .X(_07878_));
 sky130_fd_sc_hd__xor2_1 _15782_ (.A(_07876_),
    .B(_07878_),
    .X(_07879_));
 sky130_fd_sc_hd__xnor2_2 _15783_ (.A(_07871_),
    .B(_07879_),
    .Y(_07880_));
 sky130_fd_sc_hd__xor2_1 _15784_ (.A(_07869_),
    .B(_07880_),
    .X(_07881_));
 sky130_fd_sc_hd__xnor2_1 _15785_ (.A(_07867_),
    .B(_07881_),
    .Y(_07882_));
 sky130_fd_sc_hd__nand2_1 _15786_ (.A(_07765_),
    .B(_07770_),
    .Y(_07883_));
 sky130_fd_sc_hd__or3_1 _15787_ (.A(net508),
    .B(_07618_),
    .C(_07619_),
    .X(_07884_));
 sky130_fd_sc_hd__a21oi_1 _15788_ (.A1(_07765_),
    .A2(_07884_),
    .B1(_07770_),
    .Y(_07885_));
 sky130_fd_sc_hd__a31o_1 _15789_ (.A1(net508),
    .A2(_07767_),
    .A3(_07883_),
    .B1(_07885_),
    .X(_07886_));
 sky130_fd_sc_hd__a21o_1 _15790_ (.A1(net508),
    .A2(net481),
    .B1(_07767_),
    .X(_07887_));
 sky130_fd_sc_hd__o2bb2a_1 _15791_ (.A1_N(net481),
    .A2_N(_07886_),
    .B1(_07887_),
    .B2(_07765_),
    .X(_07888_));
 sky130_fd_sc_hd__o21ba_1 _15792_ (.A1(_07718_),
    .A2(_07776_),
    .B1_N(_07775_),
    .X(_07889_));
 sky130_fd_sc_hd__xnor2_1 _15793_ (.A(_07888_),
    .B(_07889_),
    .Y(_07890_));
 sky130_fd_sc_hd__xnor2_1 _15794_ (.A(_07882_),
    .B(_07890_),
    .Y(_07891_));
 sky130_fd_sc_hd__nor2_1 _15795_ (.A(_07812_),
    .B(_07891_),
    .Y(_07892_));
 sky130_fd_sc_hd__nand2_1 _15796_ (.A(_07812_),
    .B(_07891_),
    .Y(_07893_));
 sky130_fd_sc_hd__and2b_1 _15797_ (.A_N(_07892_),
    .B(_07893_),
    .X(_07894_));
 sky130_fd_sc_hd__xor2_2 _15798_ (.A(_07810_),
    .B(_07894_),
    .X(_07895_));
 sky130_fd_sc_hd__and3_1 _15799_ (.A(net549),
    .B(_07699_),
    .C(_07895_),
    .X(_07896_));
 sky130_fd_sc_hd__a221o_1 _15800_ (.A1(\top0.pid_q.out[2] ),
    .A2(_07704_),
    .B1(_07806_),
    .B2(net544),
    .C1(_07896_),
    .X(_07897_));
 sky130_fd_sc_hd__and2_1 _15801_ (.A(_07800_),
    .B(_07897_),
    .X(_07898_));
 sky130_fd_sc_hd__clkbuf_1 _15802_ (.A(_07898_),
    .X(_00135_));
 sky130_fd_sc_hd__a22oi_2 _15803_ (.A1(\top0.pid_q.out[2] ),
    .A2(\top0.pid_q.curr_int[2] ),
    .B1(_07802_),
    .B2(_07803_),
    .Y(_07899_));
 sky130_fd_sc_hd__nor2_1 _15804_ (.A(\top0.pid_q.out[2] ),
    .B(\top0.pid_q.curr_int[2] ),
    .Y(_07900_));
 sky130_fd_sc_hd__nor2_1 _15805_ (.A(_07899_),
    .B(_07900_),
    .Y(_07901_));
 sky130_fd_sc_hd__xor2_1 _15806_ (.A(\top0.pid_q.out[3] ),
    .B(\top0.pid_q.curr_int[3] ),
    .X(_07902_));
 sky130_fd_sc_hd__or2_1 _15807_ (.A(_07901_),
    .B(_07902_),
    .X(_07903_));
 sky130_fd_sc_hd__nand2_1 _15808_ (.A(_07901_),
    .B(_07902_),
    .Y(_07904_));
 sky130_fd_sc_hd__a21o_1 _15809_ (.A1(_07810_),
    .A2(_07893_),
    .B1(_07892_),
    .X(_07905_));
 sky130_fd_sc_hd__nand2_2 _15810_ (.A(net469),
    .B(net512),
    .Y(_07906_));
 sky130_fd_sc_hd__nand2_2 _15811_ (.A(net477),
    .B(net506),
    .Y(_07907_));
 sky130_fd_sc_hd__nand2_2 _15812_ (.A(net474),
    .B(net509),
    .Y(_07908_));
 sky130_fd_sc_hd__xnor2_2 _15813_ (.A(_07907_),
    .B(_07908_),
    .Y(_07909_));
 sky130_fd_sc_hd__xnor2_4 _15814_ (.A(_07906_),
    .B(_07909_),
    .Y(_07910_));
 sky130_fd_sc_hd__nand2_1 _15815_ (.A(_07813_),
    .B(_07815_),
    .Y(_07911_));
 sky130_fd_sc_hd__nor2_1 _15816_ (.A(_07813_),
    .B(_07815_),
    .Y(_07912_));
 sky130_fd_sc_hd__a31o_1 _15817_ (.A1(net469),
    .A2(net515),
    .A3(_07911_),
    .B1(_07912_),
    .X(_07913_));
 sky130_fd_sc_hd__xor2_4 _15818_ (.A(net496),
    .B(net492),
    .X(_07914_));
 sky130_fd_sc_hd__nand2_1 _15819_ (.A(net499),
    .B(_07914_),
    .Y(_07915_));
 sky130_fd_sc_hd__nand2_1 _15820_ (.A(net488),
    .B(net502),
    .Y(_07916_));
 sky130_fd_sc_hd__xor2_2 _15821_ (.A(_07915_),
    .B(_07916_),
    .X(_07917_));
 sky130_fd_sc_hd__xor2_2 _15822_ (.A(_07913_),
    .B(_07917_),
    .X(_07918_));
 sky130_fd_sc_hd__xnor2_4 _15823_ (.A(_07910_),
    .B(_07918_),
    .Y(_07919_));
 sky130_fd_sc_hd__a21bo_1 _15824_ (.A1(_07855_),
    .A2(_07857_),
    .B1_N(_07853_),
    .X(_07920_));
 sky130_fd_sc_hd__o21ai_1 _15825_ (.A1(_07855_),
    .A2(_07857_),
    .B1(_07920_),
    .Y(_07921_));
 sky130_fd_sc_hd__o21a_1 _15826_ (.A1(_07819_),
    .A2(_07824_),
    .B1(_07817_),
    .X(_07922_));
 sky130_fd_sc_hd__a21o_1 _15827_ (.A1(_07819_),
    .A2(_07824_),
    .B1(_07922_),
    .X(_07923_));
 sky130_fd_sc_hd__nand2_1 _15828_ (.A(_07921_),
    .B(_07923_),
    .Y(_07924_));
 sky130_fd_sc_hd__nor2_1 _15829_ (.A(_07921_),
    .B(_07923_),
    .Y(_07925_));
 sky130_fd_sc_hd__inv_2 _15830_ (.A(_07925_),
    .Y(_07926_));
 sky130_fd_sc_hd__nand2_2 _15831_ (.A(_07924_),
    .B(_07926_),
    .Y(_07927_));
 sky130_fd_sc_hd__xnor2_4 _15832_ (.A(_07919_),
    .B(_07927_),
    .Y(_07928_));
 sky130_fd_sc_hd__o21a_1 _15833_ (.A1(_07847_),
    .A2(_07859_),
    .B1(_07848_),
    .X(_07929_));
 sky130_fd_sc_hd__a21o_1 _15834_ (.A1(_07847_),
    .A2(_07859_),
    .B1(_07929_),
    .X(_07930_));
 sky130_fd_sc_hd__a21bo_1 _15835_ (.A1(_07838_),
    .A2(_07842_),
    .B1_N(_07839_),
    .X(_07931_));
 sky130_fd_sc_hd__o21ai_2 _15836_ (.A1(_07838_),
    .A2(_07842_),
    .B1(_07931_),
    .Y(_07932_));
 sky130_fd_sc_hd__nand2b_2 _15837_ (.A_N(net538),
    .B(net443),
    .Y(_07933_));
 sky130_fd_sc_hd__nand2_1 _15838_ (.A(net448),
    .B(net532),
    .Y(_07934_));
 sky130_fd_sc_hd__nand2_1 _15839_ (.A(net536),
    .B(net446),
    .Y(_07935_));
 sky130_fd_sc_hd__xnor2_1 _15840_ (.A(_07934_),
    .B(_07935_),
    .Y(_07936_));
 sky130_fd_sc_hd__xnor2_1 _15841_ (.A(_07933_),
    .B(_07936_),
    .Y(_07937_));
 sky130_fd_sc_hd__nand2_2 _15842_ (.A(net455),
    .B(net523),
    .Y(_07938_));
 sky130_fd_sc_hd__nand2_1 _15843_ (.A(net451),
    .B(net529),
    .Y(_07939_));
 sky130_fd_sc_hd__nand2_1 _15844_ (.A(net454),
    .B(net526),
    .Y(_07940_));
 sky130_fd_sc_hd__xor2_1 _15845_ (.A(_07939_),
    .B(_07940_),
    .X(_07941_));
 sky130_fd_sc_hd__xnor2_2 _15846_ (.A(_07938_),
    .B(_07941_),
    .Y(_07942_));
 sky130_fd_sc_hd__xor2_1 _15847_ (.A(_07937_),
    .B(_07942_),
    .X(_07943_));
 sky130_fd_sc_hd__xnor2_2 _15848_ (.A(_07932_),
    .B(_07943_),
    .Y(_07944_));
 sky130_fd_sc_hd__and2b_1 _15849_ (.A_N(_07839_),
    .B(_07838_),
    .X(_07945_));
 sky130_fd_sc_hd__o221a_1 _15850_ (.A1(_07839_),
    .A2(_07843_),
    .B1(_07945_),
    .B2(_07182_),
    .C1(_07845_),
    .X(_07946_));
 sky130_fd_sc_hd__o32a_1 _15851_ (.A1(net536),
    .A2(_07649_),
    .A3(_07838_),
    .B1(_07946_),
    .B2(_07837_),
    .X(_07947_));
 sky130_fd_sc_hd__nand2_1 _15852_ (.A(net467),
    .B(net515),
    .Y(_07948_));
 sky130_fd_sc_hd__nand2_1 _15853_ (.A(net458),
    .B(net521),
    .Y(_07949_));
 sky130_fd_sc_hd__nand2_1 _15854_ (.A(net461),
    .B(net519),
    .Y(_07950_));
 sky130_fd_sc_hd__xnor2_1 _15855_ (.A(_07949_),
    .B(_07950_),
    .Y(_07951_));
 sky130_fd_sc_hd__xnor2_1 _15856_ (.A(_07948_),
    .B(_07951_),
    .Y(_07952_));
 sky130_fd_sc_hd__o21a_1 _15857_ (.A1(_07833_),
    .A2(_07835_),
    .B1(_07834_),
    .X(_07953_));
 sky130_fd_sc_hd__a21oi_2 _15858_ (.A1(_07833_),
    .A2(_07835_),
    .B1(_07953_),
    .Y(_07954_));
 sky130_fd_sc_hd__o21a_1 _15859_ (.A1(_07849_),
    .A2(_07851_),
    .B1(_07850_),
    .X(_07955_));
 sky130_fd_sc_hd__a21oi_2 _15860_ (.A1(_07849_),
    .A2(_07851_),
    .B1(_07955_),
    .Y(_07956_));
 sky130_fd_sc_hd__xnor2_1 _15861_ (.A(_07954_),
    .B(_07956_),
    .Y(_07957_));
 sky130_fd_sc_hd__xnor2_1 _15862_ (.A(_07952_),
    .B(_07957_),
    .Y(_07958_));
 sky130_fd_sc_hd__nor2_1 _15863_ (.A(_07947_),
    .B(_07958_),
    .Y(_07959_));
 sky130_fd_sc_hd__nand2_1 _15864_ (.A(_07947_),
    .B(_07958_),
    .Y(_07960_));
 sky130_fd_sc_hd__or2b_1 _15865_ (.A(_07959_),
    .B_N(_07960_),
    .X(_07961_));
 sky130_fd_sc_hd__xnor2_2 _15866_ (.A(_07944_),
    .B(_07961_),
    .Y(_07962_));
 sky130_fd_sc_hd__xor2_1 _15867_ (.A(_07930_),
    .B(_07962_),
    .X(_07963_));
 sky130_fd_sc_hd__xnor2_2 _15868_ (.A(_07928_),
    .B(_07963_),
    .Y(_07964_));
 sky130_fd_sc_hd__o21ba_1 _15869_ (.A1(_07832_),
    .A2(_07864_),
    .B1_N(_07865_),
    .X(_07965_));
 sky130_fd_sc_hd__o21a_1 _15870_ (.A1(_07828_),
    .A2(_07830_),
    .B1(_07826_),
    .X(_07966_));
 sky130_fd_sc_hd__a21oi_1 _15871_ (.A1(_07828_),
    .A2(_07830_),
    .B1(_07966_),
    .Y(_07967_));
 sky130_fd_sc_hd__a21bo_1 _15872_ (.A1(net443),
    .A2(_07873_),
    .B1_N(_07874_),
    .X(_07968_));
 sky130_fd_sc_hd__o21a_1 _15873_ (.A1(net443),
    .A2(_07873_),
    .B1(_07968_),
    .X(_07969_));
 sky130_fd_sc_hd__nand2_1 _15874_ (.A(net505),
    .B(net483),
    .Y(_07970_));
 sky130_fd_sc_hd__o21ai_1 _15875_ (.A1(_07821_),
    .A2(_07822_),
    .B1(_07820_),
    .Y(_07971_));
 sky130_fd_sc_hd__a21boi_2 _15876_ (.A1(_07821_),
    .A2(_07822_),
    .B1_N(_07971_),
    .Y(_07972_));
 sky130_fd_sc_hd__xnor2_2 _15877_ (.A(_07970_),
    .B(_07972_),
    .Y(_07973_));
 sky130_fd_sc_hd__xor2_1 _15878_ (.A(_07969_),
    .B(_07973_),
    .X(_07974_));
 sky130_fd_sc_hd__xnor2_1 _15879_ (.A(_07967_),
    .B(_07974_),
    .Y(_07975_));
 sky130_fd_sc_hd__nor2_1 _15880_ (.A(_07965_),
    .B(_07975_),
    .Y(_07976_));
 sky130_fd_sc_hd__nand2_1 _15881_ (.A(_07965_),
    .B(_07975_),
    .Y(_07977_));
 sky130_fd_sc_hd__or2b_1 _15882_ (.A(_07976_),
    .B_N(_07977_),
    .X(_07978_));
 sky130_fd_sc_hd__xnor2_1 _15883_ (.A(_07964_),
    .B(_07978_),
    .Y(_07979_));
 sky130_fd_sc_hd__inv_2 _15884_ (.A(_07869_),
    .Y(_07980_));
 sky130_fd_sc_hd__nand2_1 _15885_ (.A(_07980_),
    .B(_07880_),
    .Y(_07981_));
 sky130_fd_sc_hd__nor2_1 _15886_ (.A(_07980_),
    .B(_07880_),
    .Y(_07982_));
 sky130_fd_sc_hd__a21o_1 _15887_ (.A1(_07867_),
    .A2(_07981_),
    .B1(_07982_),
    .X(_07983_));
 sky130_fd_sc_hd__o21ba_1 _15888_ (.A1(_07876_),
    .A2(_07878_),
    .B1_N(_07871_),
    .X(_07984_));
 sky130_fd_sc_hd__a21o_1 _15889_ (.A1(_07876_),
    .A2(_07878_),
    .B1(_07984_),
    .X(_07985_));
 sky130_fd_sc_hd__xor2_1 _15890_ (.A(_07983_),
    .B(_07985_),
    .X(_07986_));
 sky130_fd_sc_hd__xnor2_1 _15891_ (.A(_07979_),
    .B(_07986_),
    .Y(_07987_));
 sky130_fd_sc_hd__a21o_1 _15892_ (.A1(_07888_),
    .A2(_07889_),
    .B1(_07882_),
    .X(_07988_));
 sky130_fd_sc_hd__o21ai_2 _15893_ (.A1(_07888_),
    .A2(_07889_),
    .B1(_07988_),
    .Y(_07989_));
 sky130_fd_sc_hd__xnor2_1 _15894_ (.A(_07987_),
    .B(_07989_),
    .Y(_07990_));
 sky130_fd_sc_hd__xnor2_1 _15895_ (.A(_07905_),
    .B(_07990_),
    .Y(_07991_));
 sky130_fd_sc_hd__a32o_1 _15896_ (.A1(net545),
    .A2(_07903_),
    .A3(_07904_),
    .B1(net548),
    .B2(_07991_),
    .X(_07992_));
 sky130_fd_sc_hd__inv_2 _15897_ (.A(\top0.pid_q.out[3] ),
    .Y(_07993_));
 sky130_fd_sc_hd__nand2_1 _15898_ (.A(_07993_),
    .B(_07705_),
    .Y(_07994_));
 sky130_fd_sc_hd__o211a_1 _15899_ (.A1(_07705_),
    .A2(_07992_),
    .B1(_07994_),
    .C1(_07710_),
    .X(_00136_));
 sky130_fd_sc_hd__nand2_1 _15900_ (.A(_07987_),
    .B(_07989_),
    .Y(_07995_));
 sky130_fd_sc_hd__inv_2 _15901_ (.A(_07995_),
    .Y(_07996_));
 sky130_fd_sc_hd__or2_1 _15902_ (.A(_07987_),
    .B(_07989_),
    .X(_07997_));
 sky130_fd_sc_hd__o21ai_1 _15903_ (.A1(_07905_),
    .A2(_07996_),
    .B1(_07997_),
    .Y(_07998_));
 sky130_fd_sc_hd__a21bo_1 _15904_ (.A1(_07928_),
    .A2(_07962_),
    .B1_N(_07930_),
    .X(_07999_));
 sky130_fd_sc_hd__o21ai_4 _15905_ (.A1(_07928_),
    .A2(_07962_),
    .B1(_07999_),
    .Y(_08000_));
 sky130_fd_sc_hd__o21a_1 _15906_ (.A1(_07919_),
    .A2(_07925_),
    .B1(_07924_),
    .X(_08001_));
 sky130_fd_sc_hd__or2_1 _15907_ (.A(net496),
    .B(net492),
    .X(_08002_));
 sky130_fd_sc_hd__a21o_2 _15908_ (.A1(net493),
    .A2(_07227_),
    .B1(_07228_),
    .X(_08003_));
 sky130_fd_sc_hd__nand2_1 _15909_ (.A(net499),
    .B(_08003_),
    .Y(_08004_));
 sky130_fd_sc_hd__a32o_1 _15910_ (.A1(net499),
    .A2(_07367_),
    .A3(_08002_),
    .B1(_08004_),
    .B2(net483),
    .X(_08005_));
 sky130_fd_sc_hd__a21oi_1 _15911_ (.A1(net483),
    .A2(net502),
    .B1(_07485_),
    .Y(_08006_));
 sky130_fd_sc_hd__a22o_1 _15912_ (.A1(net502),
    .A2(_08005_),
    .B1(_08006_),
    .B2(net499),
    .X(_08007_));
 sky130_fd_sc_hd__and3_1 _15913_ (.A(net505),
    .B(net483),
    .C(_07972_),
    .X(_08008_));
 sky130_fd_sc_hd__xnor2_1 _15914_ (.A(_08007_),
    .B(_08008_),
    .Y(_08009_));
 sky130_fd_sc_hd__xnor2_1 _15915_ (.A(_08001_),
    .B(_08009_),
    .Y(_08010_));
 sky130_fd_sc_hd__a21bo_1 _15916_ (.A1(_07932_),
    .A2(_07942_),
    .B1_N(_07937_),
    .X(_08011_));
 sky130_fd_sc_hd__o21a_2 _15917_ (.A1(_07932_),
    .A2(_07942_),
    .B1(_08011_),
    .X(_08012_));
 sky130_fd_sc_hd__nand2_1 _15918_ (.A(net455),
    .B(net521),
    .Y(_08013_));
 sky130_fd_sc_hd__nand2_1 _15919_ (.A(net451),
    .B(net526),
    .Y(_08014_));
 sky130_fd_sc_hd__nand2_1 _15920_ (.A(net453),
    .B(net523),
    .Y(_08015_));
 sky130_fd_sc_hd__xnor2_1 _15921_ (.A(_08014_),
    .B(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__xnor2_1 _15922_ (.A(_08013_),
    .B(_08016_),
    .Y(_08017_));
 sky130_fd_sc_hd__o21a_1 _15923_ (.A1(_07933_),
    .A2(_07935_),
    .B1(_07934_),
    .X(_08018_));
 sky130_fd_sc_hd__a21oi_2 _15924_ (.A1(_07933_),
    .A2(_07935_),
    .B1(_08018_),
    .Y(_08019_));
 sky130_fd_sc_hd__nand2b_2 _15925_ (.A_N(net536),
    .B(net443),
    .Y(_08020_));
 sky130_fd_sc_hd__nand2_1 _15926_ (.A(net448),
    .B(net529),
    .Y(_08021_));
 sky130_fd_sc_hd__nand2_1 _15927_ (.A(net532),
    .B(net446),
    .Y(_08022_));
 sky130_fd_sc_hd__xor2_2 _15928_ (.A(_08021_),
    .B(_08022_),
    .X(_08023_));
 sky130_fd_sc_hd__xnor2_2 _15929_ (.A(_08020_),
    .B(_08023_),
    .Y(_08024_));
 sky130_fd_sc_hd__xnor2_1 _15930_ (.A(_08019_),
    .B(_08024_),
    .Y(_08025_));
 sky130_fd_sc_hd__xnor2_1 _15931_ (.A(_08017_),
    .B(_08025_),
    .Y(_08026_));
 sky130_fd_sc_hd__nand2_2 _15932_ (.A(net467),
    .B(net1029),
    .Y(_08027_));
 sky130_fd_sc_hd__nand2_1 _15933_ (.A(net458),
    .B(net1028),
    .Y(_08028_));
 sky130_fd_sc_hd__nand2_1 _15934_ (.A(net461),
    .B(net516),
    .Y(_08029_));
 sky130_fd_sc_hd__xnor2_1 _15935_ (.A(_08028_),
    .B(_08029_),
    .Y(_08030_));
 sky130_fd_sc_hd__xnor2_2 _15936_ (.A(_08027_),
    .B(_08030_),
    .Y(_08031_));
 sky130_fd_sc_hd__o21a_1 _15937_ (.A1(_07938_),
    .A2(_07940_),
    .B1(_07939_),
    .X(_08032_));
 sky130_fd_sc_hd__a21oi_2 _15938_ (.A1(_07938_),
    .A2(_07940_),
    .B1(_08032_),
    .Y(_08033_));
 sky130_fd_sc_hd__o21a_1 _15939_ (.A1(_07948_),
    .A2(_07950_),
    .B1(_07949_),
    .X(_08034_));
 sky130_fd_sc_hd__a21oi_2 _15940_ (.A1(_07948_),
    .A2(_07950_),
    .B1(_08034_),
    .Y(_08035_));
 sky130_fd_sc_hd__xor2_1 _15941_ (.A(_08033_),
    .B(_08035_),
    .X(_08036_));
 sky130_fd_sc_hd__xnor2_2 _15942_ (.A(_08031_),
    .B(_08036_),
    .Y(_08037_));
 sky130_fd_sc_hd__xnor2_1 _15943_ (.A(_08026_),
    .B(_08037_),
    .Y(_08038_));
 sky130_fd_sc_hd__xnor2_2 _15944_ (.A(_08012_),
    .B(_08038_),
    .Y(_08039_));
 sky130_fd_sc_hd__o21a_1 _15945_ (.A1(_07944_),
    .A2(_07959_),
    .B1(_07960_),
    .X(_08040_));
 sky130_fd_sc_hd__nand2_1 _15946_ (.A(net468),
    .B(net509),
    .Y(_08041_));
 sky130_fd_sc_hd__nand2_1 _15947_ (.A(net477),
    .B(net505),
    .Y(_08042_));
 sky130_fd_sc_hd__nand2_1 _15948_ (.A(net474),
    .B(net506),
    .Y(_08043_));
 sky130_fd_sc_hd__xor2_1 _15949_ (.A(_08042_),
    .B(_08043_),
    .X(_08044_));
 sky130_fd_sc_hd__xnor2_2 _15950_ (.A(_08041_),
    .B(_08044_),
    .Y(_08045_));
 sky130_fd_sc_hd__o21ai_1 _15951_ (.A1(_07907_),
    .A2(_07908_),
    .B1(_07906_),
    .Y(_08046_));
 sky130_fd_sc_hd__a21bo_1 _15952_ (.A1(_07907_),
    .A2(_07908_),
    .B1_N(_08046_),
    .X(_08047_));
 sky130_fd_sc_hd__xor2_4 _15953_ (.A(net488),
    .B(_07914_),
    .X(_08048_));
 sky130_fd_sc_hd__nand2_4 _15954_ (.A(net499),
    .B(_08048_),
    .Y(_08049_));
 sky130_fd_sc_hd__nor2_1 _15955_ (.A(_08047_),
    .B(_08049_),
    .Y(_08050_));
 sky130_fd_sc_hd__nand2_1 _15956_ (.A(_08047_),
    .B(_08049_),
    .Y(_08051_));
 sky130_fd_sc_hd__and2b_1 _15957_ (.A_N(_08050_),
    .B(_08051_),
    .X(_08052_));
 sky130_fd_sc_hd__xnor2_2 _15958_ (.A(_08045_),
    .B(_08052_),
    .Y(_08053_));
 sky130_fd_sc_hd__a21bo_1 _15959_ (.A1(_07954_),
    .A2(_07956_),
    .B1_N(_07952_),
    .X(_08054_));
 sky130_fd_sc_hd__o21a_1 _15960_ (.A1(_07954_),
    .A2(_07956_),
    .B1(_08054_),
    .X(_08055_));
 sky130_fd_sc_hd__a21bo_1 _15961_ (.A1(_07913_),
    .A2(_07917_),
    .B1_N(_07910_),
    .X(_08056_));
 sky130_fd_sc_hd__o21a_1 _15962_ (.A1(_07913_),
    .A2(_07917_),
    .B1(_08056_),
    .X(_08057_));
 sky130_fd_sc_hd__xnor2_1 _15963_ (.A(_08055_),
    .B(_08057_),
    .Y(_08058_));
 sky130_fd_sc_hd__xnor2_2 _15964_ (.A(_08053_),
    .B(_08058_),
    .Y(_08059_));
 sky130_fd_sc_hd__xor2_1 _15965_ (.A(_08040_),
    .B(_08059_),
    .X(_08060_));
 sky130_fd_sc_hd__xnor2_2 _15966_ (.A(_08039_),
    .B(_08060_),
    .Y(_08061_));
 sky130_fd_sc_hd__xnor2_1 _15967_ (.A(_08010_),
    .B(_08061_),
    .Y(_08062_));
 sky130_fd_sc_hd__xnor2_2 _15968_ (.A(_08000_),
    .B(_08062_),
    .Y(_08063_));
 sky130_fd_sc_hd__o21a_1 _15969_ (.A1(_07964_),
    .A2(_07976_),
    .B1(_07977_),
    .X(_08064_));
 sky130_fd_sc_hd__a21o_1 _15970_ (.A1(_07969_),
    .A2(_07973_),
    .B1(_07967_),
    .X(_08065_));
 sky130_fd_sc_hd__o21a_1 _15971_ (.A1(_07969_),
    .A2(_07973_),
    .B1(_08065_),
    .X(_08066_));
 sky130_fd_sc_hd__xor2_1 _15972_ (.A(_08064_),
    .B(_08066_),
    .X(_08067_));
 sky130_fd_sc_hd__xnor2_1 _15973_ (.A(_08063_),
    .B(_08067_),
    .Y(_08068_));
 sky130_fd_sc_hd__or2b_1 _15974_ (.A(_07985_),
    .B_N(_07983_),
    .X(_08069_));
 sky130_fd_sc_hd__and2b_1 _15975_ (.A_N(_07983_),
    .B(_07985_),
    .X(_08070_));
 sky130_fd_sc_hd__a21oi_1 _15976_ (.A1(_07979_),
    .A2(_08069_),
    .B1(_08070_),
    .Y(_08071_));
 sky130_fd_sc_hd__nor2_1 _15977_ (.A(_08068_),
    .B(_08071_),
    .Y(_08072_));
 sky130_fd_sc_hd__nand2_1 _15978_ (.A(_08068_),
    .B(_08071_),
    .Y(_08073_));
 sky130_fd_sc_hd__or2b_1 _15979_ (.A(_08072_),
    .B_N(_08073_),
    .X(_08074_));
 sky130_fd_sc_hd__xor2_1 _15980_ (.A(_07998_),
    .B(_08074_),
    .X(_08075_));
 sky130_fd_sc_hd__inv_2 _15981_ (.A(\top0.pid_q.curr_int[3] ),
    .Y(_08076_));
 sky130_fd_sc_hd__o31a_1 _15982_ (.A1(_08076_),
    .A2(_07899_),
    .A3(_07900_),
    .B1(_07993_),
    .X(_08077_));
 sky130_fd_sc_hd__o21ba_1 _15983_ (.A1(\top0.pid_q.curr_int[3] ),
    .A2(_07901_),
    .B1_N(_08077_),
    .X(_08078_));
 sky130_fd_sc_hd__xnor2_1 _15984_ (.A(\top0.pid_q.out[4] ),
    .B(\top0.pid_q.curr_int[4] ),
    .Y(_08079_));
 sky130_fd_sc_hd__xnor2_1 _15985_ (.A(_08078_),
    .B(_08079_),
    .Y(_08080_));
 sky130_fd_sc_hd__a221o_1 _15986_ (.A1(net548),
    .A2(_08075_),
    .B1(_08080_),
    .B2(net545),
    .C1(_07705_),
    .X(_08081_));
 sky130_fd_sc_hd__o211a_1 _15987_ (.A1(\top0.pid_q.out[4] ),
    .A2(_07700_),
    .B1(_08081_),
    .C1(_07710_),
    .X(_00137_));
 sky130_fd_sc_hd__a21o_1 _15988_ (.A1(\top0.pid_q.curr_int[4] ),
    .A2(_08078_),
    .B1(\top0.pid_q.out[4] ),
    .X(_08082_));
 sky130_fd_sc_hd__o21a_1 _15989_ (.A1(\top0.pid_q.curr_int[4] ),
    .A2(_08078_),
    .B1(_08082_),
    .X(_08083_));
 sky130_fd_sc_hd__xor2_1 _15990_ (.A(\top0.pid_q.out[5] ),
    .B(\top0.pid_q.curr_int[5] ),
    .X(_08084_));
 sky130_fd_sc_hd__or2_1 _15991_ (.A(_08083_),
    .B(_08084_),
    .X(_08085_));
 sky130_fd_sc_hd__nand2_1 _15992_ (.A(_08083_),
    .B(_08084_),
    .Y(_08086_));
 sky130_fd_sc_hd__a21bo_1 _15993_ (.A1(_07905_),
    .A2(_07997_),
    .B1_N(_07995_),
    .X(_08087_));
 sky130_fd_sc_hd__a21o_1 _15994_ (.A1(_08073_),
    .A2(_08087_),
    .B1(_08072_),
    .X(_08088_));
 sky130_fd_sc_hd__o21ba_1 _15995_ (.A1(_08000_),
    .A2(_08061_),
    .B1_N(_08010_),
    .X(_08089_));
 sky130_fd_sc_hd__a21oi_2 _15996_ (.A1(_08000_),
    .A2(_08061_),
    .B1(_08089_),
    .Y(_08090_));
 sky130_fd_sc_hd__a21bo_1 _15997_ (.A1(_08012_),
    .A2(_08037_),
    .B1_N(_08026_),
    .X(_08091_));
 sky130_fd_sc_hd__o21ai_2 _15998_ (.A1(_08012_),
    .A2(_08037_),
    .B1(_08091_),
    .Y(_08092_));
 sky130_fd_sc_hd__nand2b_2 _15999_ (.A_N(net532),
    .B(\top0.pid_q.mult0.b[15] ),
    .Y(_08093_));
 sky130_fd_sc_hd__nand2_1 _16000_ (.A(net448),
    .B(net526),
    .Y(_08094_));
 sky130_fd_sc_hd__nand2_1 _16001_ (.A(net529),
    .B(net446),
    .Y(_08095_));
 sky130_fd_sc_hd__xnor2_1 _16002_ (.A(_08094_),
    .B(_08095_),
    .Y(_08096_));
 sky130_fd_sc_hd__xnor2_2 _16003_ (.A(_08093_),
    .B(_08096_),
    .Y(_08097_));
 sky130_fd_sc_hd__o21a_1 _16004_ (.A1(_08020_),
    .A2(_08022_),
    .B1(_08021_),
    .X(_08098_));
 sky130_fd_sc_hd__a21oi_1 _16005_ (.A1(_08020_),
    .A2(_08022_),
    .B1(_08098_),
    .Y(_08099_));
 sky130_fd_sc_hd__nand2_2 _16006_ (.A(net456),
    .B(net1028),
    .Y(_08100_));
 sky130_fd_sc_hd__nand2_1 _16007_ (.A(net449),
    .B(net523),
    .Y(_08101_));
 sky130_fd_sc_hd__nand2_1 _16008_ (.A(net453),
    .B(net521),
    .Y(_08102_));
 sky130_fd_sc_hd__xnor2_1 _16009_ (.A(_08101_),
    .B(_08102_),
    .Y(_08103_));
 sky130_fd_sc_hd__xnor2_2 _16010_ (.A(_08100_),
    .B(_08103_),
    .Y(_08104_));
 sky130_fd_sc_hd__xor2_1 _16011_ (.A(_08099_),
    .B(_08104_),
    .X(_08105_));
 sky130_fd_sc_hd__xnor2_1 _16012_ (.A(_08097_),
    .B(_08105_),
    .Y(_08106_));
 sky130_fd_sc_hd__a21bo_1 _16013_ (.A1(_08019_),
    .A2(_08024_),
    .B1_N(_08017_),
    .X(_08107_));
 sky130_fd_sc_hd__o21a_1 _16014_ (.A1(_08019_),
    .A2(_08024_),
    .B1(_08107_),
    .X(_08108_));
 sky130_fd_sc_hd__nand2_1 _16015_ (.A(net461),
    .B(net1029),
    .Y(_08109_));
 sky130_fd_sc_hd__nand2_1 _16016_ (.A(net458),
    .B(net516),
    .Y(_08110_));
 sky130_fd_sc_hd__nand2_1 _16017_ (.A(net467),
    .B(net510),
    .Y(_08111_));
 sky130_fd_sc_hd__xnor2_1 _16018_ (.A(_08110_),
    .B(_08111_),
    .Y(_08112_));
 sky130_fd_sc_hd__xnor2_1 _16019_ (.A(_08109_),
    .B(_08112_),
    .Y(_08113_));
 sky130_fd_sc_hd__o21a_1 _16020_ (.A1(_08013_),
    .A2(_08015_),
    .B1(_08014_),
    .X(_08114_));
 sky130_fd_sc_hd__a21oi_2 _16021_ (.A1(_08013_),
    .A2(_08015_),
    .B1(_08114_),
    .Y(_08115_));
 sky130_fd_sc_hd__o21a_1 _16022_ (.A1(_08027_),
    .A2(_08029_),
    .B1(_08028_),
    .X(_08116_));
 sky130_fd_sc_hd__a21oi_2 _16023_ (.A1(_08027_),
    .A2(_08029_),
    .B1(_08116_),
    .Y(_08117_));
 sky130_fd_sc_hd__xor2_1 _16024_ (.A(_08115_),
    .B(_08117_),
    .X(_08118_));
 sky130_fd_sc_hd__xnor2_1 _16025_ (.A(_08113_),
    .B(_08118_),
    .Y(_08119_));
 sky130_fd_sc_hd__xor2_1 _16026_ (.A(_08108_),
    .B(_08119_),
    .X(_08120_));
 sky130_fd_sc_hd__xnor2_1 _16027_ (.A(_08106_),
    .B(_08120_),
    .Y(_08121_));
 sky130_fd_sc_hd__o21ai_1 _16028_ (.A1(_08042_),
    .A2(_08043_),
    .B1(_08041_),
    .Y(_08122_));
 sky130_fd_sc_hd__a21bo_1 _16029_ (.A1(_08042_),
    .A2(_08043_),
    .B1_N(_08122_),
    .X(_08123_));
 sky130_fd_sc_hd__nand2_1 _16030_ (.A(net476),
    .B(net502),
    .Y(_08124_));
 sky130_fd_sc_hd__nand2_1 _16031_ (.A(net474),
    .B(net503),
    .Y(_08125_));
 sky130_fd_sc_hd__nand2_1 _16032_ (.A(net468),
    .B(net507),
    .Y(_08126_));
 sky130_fd_sc_hd__xnor2_1 _16033_ (.A(_08125_),
    .B(_08126_),
    .Y(_08127_));
 sky130_fd_sc_hd__xnor2_1 _16034_ (.A(_08124_),
    .B(_08127_),
    .Y(_08128_));
 sky130_fd_sc_hd__xnor2_1 _16035_ (.A(_08123_),
    .B(_08128_),
    .Y(_08129_));
 sky130_fd_sc_hd__xnor2_1 _16036_ (.A(_08049_),
    .B(_08129_),
    .Y(_08130_));
 sky130_fd_sc_hd__a21bo_1 _16037_ (.A1(_08033_),
    .A2(_08035_),
    .B1_N(_08031_),
    .X(_08131_));
 sky130_fd_sc_hd__o21a_1 _16038_ (.A1(_08033_),
    .A2(_08035_),
    .B1(_08131_),
    .X(_08132_));
 sky130_fd_sc_hd__o21a_1 _16039_ (.A1(_08045_),
    .A2(_08050_),
    .B1(_08051_),
    .X(_08133_));
 sky130_fd_sc_hd__xnor2_1 _16040_ (.A(_08132_),
    .B(_08133_),
    .Y(_08134_));
 sky130_fd_sc_hd__xnor2_1 _16041_ (.A(_08130_),
    .B(_08134_),
    .Y(_08135_));
 sky130_fd_sc_hd__xnor2_1 _16042_ (.A(_08121_),
    .B(_08135_),
    .Y(_08136_));
 sky130_fd_sc_hd__xnor2_2 _16043_ (.A(_08092_),
    .B(_08136_),
    .Y(_08137_));
 sky130_fd_sc_hd__nor2_1 _16044_ (.A(_08039_),
    .B(_08059_),
    .Y(_08138_));
 sky130_fd_sc_hd__nand2_1 _16045_ (.A(_08039_),
    .B(_08059_),
    .Y(_08139_));
 sky130_fd_sc_hd__o21a_1 _16046_ (.A1(_08040_),
    .A2(_08138_),
    .B1(_08139_),
    .X(_08140_));
 sky130_fd_sc_hd__inv_2 _16047_ (.A(net502),
    .Y(_08141_));
 sky130_fd_sc_hd__o21ai_4 _16048_ (.A1(net483),
    .A2(_08003_),
    .B1(net499),
    .Y(_08142_));
 sky130_fd_sc_hd__a31o_1 _16049_ (.A1(net483),
    .A2(_08141_),
    .A3(_08003_),
    .B1(_08142_),
    .X(_08143_));
 sky130_fd_sc_hd__a21bo_1 _16050_ (.A1(_08055_),
    .A2(_08057_),
    .B1_N(_08053_),
    .X(_08144_));
 sky130_fd_sc_hd__o21ai_2 _16051_ (.A1(_08055_),
    .A2(_08057_),
    .B1(_08144_),
    .Y(_08145_));
 sky130_fd_sc_hd__xnor2_1 _16052_ (.A(_08143_),
    .B(_08145_),
    .Y(_08146_));
 sky130_fd_sc_hd__inv_2 _16053_ (.A(_08146_),
    .Y(_08147_));
 sky130_fd_sc_hd__xnor2_1 _16054_ (.A(_08140_),
    .B(_08147_),
    .Y(_08148_));
 sky130_fd_sc_hd__xnor2_2 _16055_ (.A(_08137_),
    .B(_08148_),
    .Y(_08149_));
 sky130_fd_sc_hd__a21o_1 _16056_ (.A1(_08001_),
    .A2(_08007_),
    .B1(_08008_),
    .X(_08150_));
 sky130_fd_sc_hd__o21ai_1 _16057_ (.A1(_08001_),
    .A2(_08007_),
    .B1(_08150_),
    .Y(_08151_));
 sky130_fd_sc_hd__xnor2_1 _16058_ (.A(_08149_),
    .B(_08151_),
    .Y(_08152_));
 sky130_fd_sc_hd__xnor2_2 _16059_ (.A(_08090_),
    .B(_08152_),
    .Y(_08153_));
 sky130_fd_sc_hd__a21o_1 _16060_ (.A1(_08063_),
    .A2(_08066_),
    .B1(_08064_),
    .X(_08154_));
 sky130_fd_sc_hd__o21ai_2 _16061_ (.A1(_08063_),
    .A2(_08066_),
    .B1(_08154_),
    .Y(_08155_));
 sky130_fd_sc_hd__xnor2_1 _16062_ (.A(_08153_),
    .B(_08155_),
    .Y(_08156_));
 sky130_fd_sc_hd__xnor2_1 _16063_ (.A(_08088_),
    .B(_08156_),
    .Y(_08157_));
 sky130_fd_sc_hd__a32o_1 _16064_ (.A1(net545),
    .A2(_08085_),
    .A3(_08086_),
    .B1(net548),
    .B2(_08157_),
    .X(_08158_));
 sky130_fd_sc_hd__mux2_1 _16065_ (.A0(\top0.pid_q.out[5] ),
    .A1(_08158_),
    .S(_07700_),
    .X(_08159_));
 sky130_fd_sc_hd__and2_1 _16066_ (.A(_07800_),
    .B(_08159_),
    .X(_08160_));
 sky130_fd_sc_hd__clkbuf_1 _16067_ (.A(_08160_),
    .X(_00138_));
 sky130_fd_sc_hd__nand2_1 _16068_ (.A(_08153_),
    .B(_08155_),
    .Y(_08161_));
 sky130_fd_sc_hd__nor2_1 _16069_ (.A(_08153_),
    .B(_08155_),
    .Y(_08162_));
 sky130_fd_sc_hd__a21oi_1 _16070_ (.A1(_08088_),
    .A2(_08161_),
    .B1(_08162_),
    .Y(_08163_));
 sky130_fd_sc_hd__a21bo_1 _16071_ (.A1(_08090_),
    .A2(_08149_),
    .B1_N(_08151_),
    .X(_08164_));
 sky130_fd_sc_hd__o21ai_1 _16072_ (.A1(_08090_),
    .A2(_08149_),
    .B1(_08164_),
    .Y(_08165_));
 sky130_fd_sc_hd__o21ai_1 _16073_ (.A1(_08124_),
    .A2(_08125_),
    .B1(_08126_),
    .Y(_08166_));
 sky130_fd_sc_hd__a21bo_1 _16074_ (.A1(_08124_),
    .A2(_08125_),
    .B1_N(_08166_),
    .X(_08167_));
 sky130_fd_sc_hd__nand2_2 _16075_ (.A(net476),
    .B(net499),
    .Y(_08168_));
 sky130_fd_sc_hd__nand2_1 _16076_ (.A(net468),
    .B(net503),
    .Y(_08169_));
 sky130_fd_sc_hd__nand2_2 _16077_ (.A(net473),
    .B(net500),
    .Y(_08170_));
 sky130_fd_sc_hd__xnor2_1 _16078_ (.A(_08169_),
    .B(_08170_),
    .Y(_08171_));
 sky130_fd_sc_hd__xnor2_2 _16079_ (.A(_08168_),
    .B(_08171_),
    .Y(_08172_));
 sky130_fd_sc_hd__xnor2_1 _16080_ (.A(_08167_),
    .B(_08172_),
    .Y(_08173_));
 sky130_fd_sc_hd__xnor2_2 _16081_ (.A(_08049_),
    .B(_08173_),
    .Y(_08174_));
 sky130_fd_sc_hd__a21bo_1 _16082_ (.A1(_08115_),
    .A2(_08117_),
    .B1_N(_08113_),
    .X(_08175_));
 sky130_fd_sc_hd__o21ai_1 _16083_ (.A1(_08115_),
    .A2(_08117_),
    .B1(_08175_),
    .Y(_08176_));
 sky130_fd_sc_hd__o21a_1 _16084_ (.A1(_08123_),
    .A2(_08128_),
    .B1(_08049_),
    .X(_08177_));
 sky130_fd_sc_hd__a21o_1 _16085_ (.A1(_08123_),
    .A2(_08128_),
    .B1(_08177_),
    .X(_08178_));
 sky130_fd_sc_hd__and2_1 _16086_ (.A(_08176_),
    .B(_08178_),
    .X(_08179_));
 sky130_fd_sc_hd__nor2_1 _16087_ (.A(_08176_),
    .B(_08178_),
    .Y(_08180_));
 sky130_fd_sc_hd__or2_1 _16088_ (.A(_08179_),
    .B(_08180_),
    .X(_08181_));
 sky130_fd_sc_hd__xnor2_2 _16089_ (.A(_08174_),
    .B(_08181_),
    .Y(_08182_));
 sky130_fd_sc_hd__a21bo_1 _16090_ (.A1(_08108_),
    .A2(_08119_),
    .B1_N(_08106_),
    .X(_08183_));
 sky130_fd_sc_hd__o21a_1 _16091_ (.A1(_08108_),
    .A2(_08119_),
    .B1(_08183_),
    .X(_08184_));
 sky130_fd_sc_hd__nand2b_1 _16092_ (.A_N(net529),
    .B(net443),
    .Y(_08185_));
 sky130_fd_sc_hd__nand2_1 _16093_ (.A(\top0.pid_q.mult0.b[13] ),
    .B(net523),
    .Y(_08186_));
 sky130_fd_sc_hd__nand2_1 _16094_ (.A(net526),
    .B(net446),
    .Y(_08187_));
 sky130_fd_sc_hd__xnor2_1 _16095_ (.A(_08186_),
    .B(_08187_),
    .Y(_08188_));
 sky130_fd_sc_hd__xnor2_1 _16096_ (.A(_08185_),
    .B(_08188_),
    .Y(_08189_));
 sky130_fd_sc_hd__o21a_1 _16097_ (.A1(_08093_),
    .A2(_08095_),
    .B1(_08094_),
    .X(_08190_));
 sky130_fd_sc_hd__a21oi_2 _16098_ (.A1(_08093_),
    .A2(_08095_),
    .B1(_08190_),
    .Y(_08191_));
 sky130_fd_sc_hd__nand2_2 _16099_ (.A(net456),
    .B(net516),
    .Y(_08192_));
 sky130_fd_sc_hd__nand2_1 _16100_ (.A(net450),
    .B(net521),
    .Y(_08193_));
 sky130_fd_sc_hd__nand2_1 _16101_ (.A(net453),
    .B(net1028),
    .Y(_08194_));
 sky130_fd_sc_hd__xor2_1 _16102_ (.A(_08193_),
    .B(_08194_),
    .X(_08195_));
 sky130_fd_sc_hd__xnor2_2 _16103_ (.A(_08192_),
    .B(_08195_),
    .Y(_08196_));
 sky130_fd_sc_hd__xnor2_1 _16104_ (.A(_08191_),
    .B(_08196_),
    .Y(_08197_));
 sky130_fd_sc_hd__xnor2_1 _16105_ (.A(_08189_),
    .B(_08197_),
    .Y(_08198_));
 sky130_fd_sc_hd__o21ba_1 _16106_ (.A1(_08097_),
    .A2(_08104_),
    .B1_N(_08099_),
    .X(_08199_));
 sky130_fd_sc_hd__a21o_1 _16107_ (.A1(_08097_),
    .A2(_08104_),
    .B1(_08199_),
    .X(_08200_));
 sky130_fd_sc_hd__and2_1 _16108_ (.A(net458),
    .B(net1029),
    .X(_08201_));
 sky130_fd_sc_hd__nand2_1 _16109_ (.A(net466),
    .B(net507),
    .Y(_08202_));
 sky130_fd_sc_hd__nand2_1 _16110_ (.A(net463),
    .B(net510),
    .Y(_08203_));
 sky130_fd_sc_hd__xor2_1 _16111_ (.A(_08202_),
    .B(_08203_),
    .X(_08204_));
 sky130_fd_sc_hd__xnor2_2 _16112_ (.A(_08201_),
    .B(_08204_),
    .Y(_08205_));
 sky130_fd_sc_hd__o21a_1 _16113_ (.A1(_08100_),
    .A2(_08102_),
    .B1(_08101_),
    .X(_08206_));
 sky130_fd_sc_hd__a21oi_2 _16114_ (.A1(_08100_),
    .A2(_08102_),
    .B1(_08206_),
    .Y(_08207_));
 sky130_fd_sc_hd__o21a_1 _16115_ (.A1(_08109_),
    .A2(_08111_),
    .B1(_08110_),
    .X(_08208_));
 sky130_fd_sc_hd__a21oi_2 _16116_ (.A1(_08109_),
    .A2(_08111_),
    .B1(_08208_),
    .Y(_08209_));
 sky130_fd_sc_hd__xnor2_1 _16117_ (.A(_08207_),
    .B(_08209_),
    .Y(_08210_));
 sky130_fd_sc_hd__xnor2_2 _16118_ (.A(_08205_),
    .B(_08210_),
    .Y(_08211_));
 sky130_fd_sc_hd__xor2_1 _16119_ (.A(_08200_),
    .B(_08211_),
    .X(_08212_));
 sky130_fd_sc_hd__xnor2_1 _16120_ (.A(_08198_),
    .B(_08212_),
    .Y(_08213_));
 sky130_fd_sc_hd__nor2_1 _16121_ (.A(_08184_),
    .B(_08213_),
    .Y(_08214_));
 sky130_fd_sc_hd__nand2_1 _16122_ (.A(_08184_),
    .B(_08213_),
    .Y(_08215_));
 sky130_fd_sc_hd__or2b_1 _16123_ (.A(_08214_),
    .B_N(_08215_),
    .X(_08216_));
 sky130_fd_sc_hd__xnor2_2 _16124_ (.A(_08182_),
    .B(_08216_),
    .Y(_08217_));
 sky130_fd_sc_hd__a21bo_1 _16125_ (.A1(_08092_),
    .A2(_08135_),
    .B1_N(_08121_),
    .X(_08218_));
 sky130_fd_sc_hd__o21a_1 _16126_ (.A1(_08092_),
    .A2(_08135_),
    .B1(_08218_),
    .X(_08219_));
 sky130_fd_sc_hd__o21a_2 _16127_ (.A1(net483),
    .A2(_08003_),
    .B1(net499),
    .X(_08220_));
 sky130_fd_sc_hd__a21bo_1 _16128_ (.A1(_08132_),
    .A2(_08133_),
    .B1_N(_08130_),
    .X(_08221_));
 sky130_fd_sc_hd__o21a_1 _16129_ (.A1(_08132_),
    .A2(_08133_),
    .B1(_08221_),
    .X(_08222_));
 sky130_fd_sc_hd__xnor2_2 _16130_ (.A(_08220_),
    .B(_08222_),
    .Y(_08223_));
 sky130_fd_sc_hd__xnor2_1 _16131_ (.A(_08219_),
    .B(_08223_),
    .Y(_08224_));
 sky130_fd_sc_hd__xor2_2 _16132_ (.A(_08217_),
    .B(_08224_),
    .X(_08225_));
 sky130_fd_sc_hd__a21o_1 _16133_ (.A1(_08140_),
    .A2(_08147_),
    .B1(_08137_),
    .X(_08226_));
 sky130_fd_sc_hd__o21a_1 _16134_ (.A1(_08140_),
    .A2(_08147_),
    .B1(_08226_),
    .X(_08227_));
 sky130_fd_sc_hd__nor2_1 _16135_ (.A(_08143_),
    .B(_08145_),
    .Y(_08228_));
 sky130_fd_sc_hd__xnor2_1 _16136_ (.A(_08227_),
    .B(_08228_),
    .Y(_08229_));
 sky130_fd_sc_hd__xor2_1 _16137_ (.A(_08225_),
    .B(_08229_),
    .X(_08230_));
 sky130_fd_sc_hd__nand2_1 _16138_ (.A(_08165_),
    .B(_08230_),
    .Y(_08231_));
 sky130_fd_sc_hd__nor2_1 _16139_ (.A(_08165_),
    .B(_08230_),
    .Y(_08232_));
 sky130_fd_sc_hd__inv_2 _16140_ (.A(_08232_),
    .Y(_08233_));
 sky130_fd_sc_hd__nand2_1 _16141_ (.A(_08231_),
    .B(_08233_),
    .Y(_08234_));
 sky130_fd_sc_hd__xnor2_1 _16142_ (.A(_08163_),
    .B(_08234_),
    .Y(_08235_));
 sky130_fd_sc_hd__nor2_1 _16143_ (.A(_07701_),
    .B(_08235_),
    .Y(_08236_));
 sky130_fd_sc_hd__nor2_1 _16144_ (.A(\top0.pid_q.out[6] ),
    .B(_07704_),
    .Y(_08237_));
 sky130_fd_sc_hd__a21o_1 _16145_ (.A1(\top0.pid_q.curr_int[5] ),
    .A2(_08083_),
    .B1(\top0.pid_q.out[5] ),
    .X(_08238_));
 sky130_fd_sc_hd__o21ai_2 _16146_ (.A1(\top0.pid_q.curr_int[5] ),
    .A2(_08083_),
    .B1(_08238_),
    .Y(_08239_));
 sky130_fd_sc_hd__xnor2_1 _16147_ (.A(\top0.pid_q.curr_int[6] ),
    .B(_08239_),
    .Y(_08240_));
 sky130_fd_sc_hd__mux2_1 _16148_ (.A0(\top0.pid_q.out[6] ),
    .A1(_08237_),
    .S(_08240_),
    .X(_08241_));
 sky130_fd_sc_hd__a22o_1 _16149_ (.A1(\top0.pid_q.out[6] ),
    .A2(_07705_),
    .B1(_08241_),
    .B2(net545),
    .X(_08242_));
 sky130_fd_sc_hd__o21a_1 _16150_ (.A1(_08236_),
    .A2(_08242_),
    .B1(_07710_),
    .X(_00139_));
 sky130_fd_sc_hd__inv_2 _16151_ (.A(\top0.pid_q.curr_int[6] ),
    .Y(_08243_));
 sky130_fd_sc_hd__o21ba_1 _16152_ (.A1(_08243_),
    .A2(_08239_),
    .B1_N(\top0.pid_q.out[6] ),
    .X(_08244_));
 sky130_fd_sc_hd__a21o_1 _16153_ (.A1(_08243_),
    .A2(_08239_),
    .B1(_08244_),
    .X(_08245_));
 sky130_fd_sc_hd__xnor2_1 _16154_ (.A(\top0.pid_q.out[7] ),
    .B(\top0.pid_q.curr_int[7] ),
    .Y(_08246_));
 sky130_fd_sc_hd__nand2_1 _16155_ (.A(_08245_),
    .B(_08246_),
    .Y(_08247_));
 sky130_fd_sc_hd__or2_1 _16156_ (.A(_08245_),
    .B(_08246_),
    .X(_08248_));
 sky130_fd_sc_hd__a211o_1 _16157_ (.A1(_08088_),
    .A2(_08161_),
    .B1(_08162_),
    .C1(_08232_),
    .X(_08249_));
 sky130_fd_sc_hd__nand2_1 _16158_ (.A(_08231_),
    .B(_08249_),
    .Y(_08250_));
 sky130_fd_sc_hd__a21o_1 _16159_ (.A1(_08227_),
    .A2(_08225_),
    .B1(_08228_),
    .X(_08251_));
 sky130_fd_sc_hd__or2_1 _16160_ (.A(_08227_),
    .B(_08225_),
    .X(_08252_));
 sky130_fd_sc_hd__a21o_1 _16161_ (.A1(_08219_),
    .A2(_08223_),
    .B1(_08217_),
    .X(_08253_));
 sky130_fd_sc_hd__o21ai_2 _16162_ (.A1(_08219_),
    .A2(_08223_),
    .B1(_08253_),
    .Y(_08254_));
 sky130_fd_sc_hd__nand2_2 _16163_ (.A(_07320_),
    .B(net444),
    .Y(_08255_));
 sky130_fd_sc_hd__nand2_1 _16164_ (.A(net447),
    .B(net521),
    .Y(_08256_));
 sky130_fd_sc_hd__nand2_2 _16165_ (.A(net523),
    .B(net446),
    .Y(_08257_));
 sky130_fd_sc_hd__xnor2_2 _16166_ (.A(_08256_),
    .B(_08257_),
    .Y(_08258_));
 sky130_fd_sc_hd__xnor2_4 _16167_ (.A(_08255_),
    .B(_08258_),
    .Y(_08259_));
 sky130_fd_sc_hd__o21a_1 _16168_ (.A1(_08185_),
    .A2(_08187_),
    .B1(_08186_),
    .X(_08260_));
 sky130_fd_sc_hd__a21oi_2 _16169_ (.A1(_08185_),
    .A2(_08187_),
    .B1(_08260_),
    .Y(_08261_));
 sky130_fd_sc_hd__nand2_2 _16170_ (.A(net456),
    .B(net1029),
    .Y(_08262_));
 sky130_fd_sc_hd__nand2_1 _16171_ (.A(net450),
    .B(net1028),
    .Y(_08263_));
 sky130_fd_sc_hd__nand2_1 _16172_ (.A(net453),
    .B(net516),
    .Y(_08264_));
 sky130_fd_sc_hd__xor2_1 _16173_ (.A(_08263_),
    .B(_08264_),
    .X(_08265_));
 sky130_fd_sc_hd__xnor2_2 _16174_ (.A(_08262_),
    .B(_08265_),
    .Y(_08266_));
 sky130_fd_sc_hd__xnor2_2 _16175_ (.A(_08261_),
    .B(_08266_),
    .Y(_08267_));
 sky130_fd_sc_hd__xnor2_4 _16176_ (.A(_08259_),
    .B(_08267_),
    .Y(_08268_));
 sky130_fd_sc_hd__a21bo_1 _16177_ (.A1(_08191_),
    .A2(_08196_),
    .B1_N(_08189_),
    .X(_08269_));
 sky130_fd_sc_hd__o21a_1 _16178_ (.A1(_08191_),
    .A2(_08196_),
    .B1(_08269_),
    .X(_08270_));
 sky130_fd_sc_hd__and2_1 _16179_ (.A(net458),
    .B(net510),
    .X(_08271_));
 sky130_fd_sc_hd__nand2_1 _16180_ (.A(net466),
    .B(net503),
    .Y(_08272_));
 sky130_fd_sc_hd__nand2_1 _16181_ (.A(net463),
    .B(net507),
    .Y(_08273_));
 sky130_fd_sc_hd__xor2_1 _16182_ (.A(_08272_),
    .B(_08273_),
    .X(_08274_));
 sky130_fd_sc_hd__xnor2_2 _16183_ (.A(_08271_),
    .B(_08274_),
    .Y(_08275_));
 sky130_fd_sc_hd__o21a_1 _16184_ (.A1(_08192_),
    .A2(_08194_),
    .B1(_08193_),
    .X(_08276_));
 sky130_fd_sc_hd__a21oi_2 _16185_ (.A1(_08192_),
    .A2(_08194_),
    .B1(_08276_),
    .Y(_08277_));
 sky130_fd_sc_hd__o21ba_1 _16186_ (.A1(_08202_),
    .A2(_08203_),
    .B1_N(_08201_),
    .X(_08278_));
 sky130_fd_sc_hd__a21oi_2 _16187_ (.A1(_08202_),
    .A2(_08203_),
    .B1(_08278_),
    .Y(_08279_));
 sky130_fd_sc_hd__xor2_1 _16188_ (.A(_08277_),
    .B(_08279_),
    .X(_08280_));
 sky130_fd_sc_hd__xnor2_2 _16189_ (.A(_08275_),
    .B(_08280_),
    .Y(_08281_));
 sky130_fd_sc_hd__xor2_2 _16190_ (.A(_08270_),
    .B(_08281_),
    .X(_08282_));
 sky130_fd_sc_hd__xnor2_4 _16191_ (.A(_08268_),
    .B(_08282_),
    .Y(_08283_));
 sky130_fd_sc_hd__o21a_1 _16192_ (.A1(_08200_),
    .A2(_08211_),
    .B1(_08198_),
    .X(_08284_));
 sky130_fd_sc_hd__a21o_1 _16193_ (.A1(_08200_),
    .A2(_08211_),
    .B1(_08284_),
    .X(_08285_));
 sky130_fd_sc_hd__inv_2 _16194_ (.A(_08049_),
    .Y(_08286_));
 sky130_fd_sc_hd__inv_2 _16195_ (.A(net504),
    .Y(_08287_));
 sky130_fd_sc_hd__and2_1 _16196_ (.A(net476),
    .B(_08287_),
    .X(_08288_));
 sky130_fd_sc_hd__o22ai_1 _16197_ (.A1(net503),
    .A2(net497),
    .B1(_08288_),
    .B2(net473),
    .Y(_08289_));
 sky130_fd_sc_hd__nor2_1 _16198_ (.A(net473),
    .B(net501),
    .Y(_08290_));
 sky130_fd_sc_hd__a21o_1 _16199_ (.A1(_08287_),
    .A2(net500),
    .B1(net476),
    .X(_08291_));
 sky130_fd_sc_hd__o21ai_1 _16200_ (.A1(net500),
    .A2(_08169_),
    .B1(_08291_),
    .Y(_08292_));
 sky130_fd_sc_hd__a21oi_1 _16201_ (.A1(_07493_),
    .A2(_08170_),
    .B1(net468),
    .Y(_08293_));
 sky130_fd_sc_hd__a221o_1 _16202_ (.A1(_08288_),
    .A2(_08290_),
    .B1(_08292_),
    .B2(net473),
    .C1(_08293_),
    .X(_08294_));
 sky130_fd_sc_hd__a32o_2 _16203_ (.A1(net468),
    .A2(net501),
    .A3(_08289_),
    .B1(_08294_),
    .B2(net497),
    .X(_08295_));
 sky130_fd_sc_hd__xnor2_2 _16204_ (.A(_08286_),
    .B(_08295_),
    .Y(_08296_));
 sky130_fd_sc_hd__a21bo_1 _16205_ (.A1(_08207_),
    .A2(_08209_),
    .B1_N(_08205_),
    .X(_08297_));
 sky130_fd_sc_hd__o21ai_1 _16206_ (.A1(_08207_),
    .A2(_08209_),
    .B1(_08297_),
    .Y(_08298_));
 sky130_fd_sc_hd__o21a_1 _16207_ (.A1(_08167_),
    .A2(_08172_),
    .B1(_08049_),
    .X(_08299_));
 sky130_fd_sc_hd__a21o_1 _16208_ (.A1(_08167_),
    .A2(_08172_),
    .B1(_08299_),
    .X(_08300_));
 sky130_fd_sc_hd__xor2_1 _16209_ (.A(_08298_),
    .B(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__xnor2_2 _16210_ (.A(_08296_),
    .B(_08301_),
    .Y(_08302_));
 sky130_fd_sc_hd__xor2_1 _16211_ (.A(_08285_),
    .B(_08302_),
    .X(_08303_));
 sky130_fd_sc_hd__xnor2_2 _16212_ (.A(_08283_),
    .B(_08303_),
    .Y(_08304_));
 sky130_fd_sc_hd__a21o_1 _16213_ (.A1(_08182_),
    .A2(_08215_),
    .B1(_08214_),
    .X(_08305_));
 sky130_fd_sc_hd__nor2_1 _16214_ (.A(_08174_),
    .B(_08179_),
    .Y(_08306_));
 sky130_fd_sc_hd__o21ai_1 _16215_ (.A1(_08180_),
    .A2(_08306_),
    .B1(_08220_),
    .Y(_08307_));
 sky130_fd_sc_hd__or3_1 _16216_ (.A(_08220_),
    .B(_08180_),
    .C(_08306_),
    .X(_08308_));
 sky130_fd_sc_hd__and2_1 _16217_ (.A(_08307_),
    .B(_08308_),
    .X(_08309_));
 sky130_fd_sc_hd__xor2_1 _16218_ (.A(_08305_),
    .B(_08309_),
    .X(_08310_));
 sky130_fd_sc_hd__xnor2_2 _16219_ (.A(_08304_),
    .B(_08310_),
    .Y(_08311_));
 sky130_fd_sc_hd__clkbuf_4 _16220_ (.A(_08220_),
    .X(_08312_));
 sky130_fd_sc_hd__and2_1 _16221_ (.A(_08312_),
    .B(_08222_),
    .X(_08313_));
 sky130_fd_sc_hd__xnor2_1 _16222_ (.A(_08311_),
    .B(_08313_),
    .Y(_08314_));
 sky130_fd_sc_hd__xnor2_1 _16223_ (.A(_08254_),
    .B(_08314_),
    .Y(_08315_));
 sky130_fd_sc_hd__a21o_1 _16224_ (.A1(_08251_),
    .A2(_08252_),
    .B1(_08315_),
    .X(_08316_));
 sky130_fd_sc_hd__and3_1 _16225_ (.A(_08315_),
    .B(_08251_),
    .C(_08252_),
    .X(_08317_));
 sky130_fd_sc_hd__inv_2 _16226_ (.A(_08317_),
    .Y(_08318_));
 sky130_fd_sc_hd__nand2_1 _16227_ (.A(_08316_),
    .B(_08318_),
    .Y(_08319_));
 sky130_fd_sc_hd__xor2_1 _16228_ (.A(_08250_),
    .B(_08319_),
    .X(_08320_));
 sky130_fd_sc_hd__a32o_1 _16229_ (.A1(net545),
    .A2(_08247_),
    .A3(_08248_),
    .B1(net548),
    .B2(_08320_),
    .X(_08321_));
 sky130_fd_sc_hd__mux2_1 _16230_ (.A0(\top0.pid_q.out[7] ),
    .A1(_08321_),
    .S(_07700_),
    .X(_08322_));
 sky130_fd_sc_hd__and2_1 _16231_ (.A(_07800_),
    .B(_08322_),
    .X(_08323_));
 sky130_fd_sc_hd__clkbuf_1 _16232_ (.A(_08323_),
    .X(_00140_));
 sky130_fd_sc_hd__inv_2 _16233_ (.A(\top0.pid_q.curr_int[7] ),
    .Y(_08324_));
 sky130_fd_sc_hd__o21ba_1 _16234_ (.A1(_08324_),
    .A2(_08245_),
    .B1_N(\top0.pid_q.out[7] ),
    .X(_08325_));
 sky130_fd_sc_hd__a21o_1 _16235_ (.A1(_08324_),
    .A2(_08245_),
    .B1(_08325_),
    .X(_08326_));
 sky130_fd_sc_hd__xnor2_1 _16236_ (.A(\top0.pid_q.out[8] ),
    .B(\top0.pid_q.curr_int[8] ),
    .Y(_08327_));
 sky130_fd_sc_hd__nand2_1 _16237_ (.A(_08326_),
    .B(_08327_),
    .Y(_08328_));
 sky130_fd_sc_hd__or2_1 _16238_ (.A(_08326_),
    .B(_08327_),
    .X(_08329_));
 sky130_fd_sc_hd__a21o_1 _16239_ (.A1(_08231_),
    .A2(_08249_),
    .B1(_08317_),
    .X(_08330_));
 sky130_fd_sc_hd__inv_2 _16240_ (.A(_08309_),
    .Y(_08331_));
 sky130_fd_sc_hd__nor2_1 _16241_ (.A(_08305_),
    .B(_08331_),
    .Y(_08332_));
 sky130_fd_sc_hd__nand2_1 _16242_ (.A(_08305_),
    .B(_08331_),
    .Y(_08333_));
 sky130_fd_sc_hd__o21a_1 _16243_ (.A1(_08304_),
    .A2(_08332_),
    .B1(_08333_),
    .X(_08334_));
 sky130_fd_sc_hd__a21boi_1 _16244_ (.A1(net503),
    .A2(_08290_),
    .B1_N(_08170_),
    .Y(_08335_));
 sky130_fd_sc_hd__o32ai_4 _16245_ (.A1(_08287_),
    .A2(net497),
    .A3(_08170_),
    .B1(_08335_),
    .B2(_08168_),
    .Y(_08336_));
 sky130_fd_sc_hd__a22oi_4 _16246_ (.A1(_08286_),
    .A2(_08295_),
    .B1(_08336_),
    .B2(net468),
    .Y(_08337_));
 sky130_fd_sc_hd__a21bo_1 _16247_ (.A1(_08277_),
    .A2(_08279_),
    .B1_N(_08275_),
    .X(_08338_));
 sky130_fd_sc_hd__o21ai_2 _16248_ (.A1(_08277_),
    .A2(_08279_),
    .B1(_08338_),
    .Y(_08339_));
 sky130_fd_sc_hd__or3_1 _16249_ (.A(net468),
    .B(net473),
    .C(net477),
    .X(_08340_));
 sky130_fd_sc_hd__o21a_1 _16250_ (.A1(net476),
    .A2(_08141_),
    .B1(net473),
    .X(_08341_));
 sky130_fd_sc_hd__a21o_1 _16251_ (.A1(net476),
    .A2(_08141_),
    .B1(_08341_),
    .X(_08342_));
 sky130_fd_sc_hd__nand2_1 _16252_ (.A(net469),
    .B(_08342_),
    .Y(_08343_));
 sky130_fd_sc_hd__and3_1 _16253_ (.A(_08048_),
    .B(_08340_),
    .C(_08343_),
    .X(_08344_));
 sky130_fd_sc_hd__a21oi_1 _16254_ (.A1(_08340_),
    .A2(_08343_),
    .B1(_08048_),
    .Y(_08345_));
 sky130_fd_sc_hd__or3b_2 _16255_ (.A(_08344_),
    .B(_08345_),
    .C_N(net497),
    .X(_08346_));
 sky130_fd_sc_hd__xnor2_1 _16256_ (.A(_08339_),
    .B(_08346_),
    .Y(_08347_));
 sky130_fd_sc_hd__xnor2_2 _16257_ (.A(_08337_),
    .B(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__o21a_1 _16258_ (.A1(_08255_),
    .A2(_08257_),
    .B1(_08256_),
    .X(_08349_));
 sky130_fd_sc_hd__a21oi_2 _16259_ (.A1(_08255_),
    .A2(_08257_),
    .B1(_08349_),
    .Y(_08350_));
 sky130_fd_sc_hd__nand2_1 _16260_ (.A(_07241_),
    .B(net444),
    .Y(_08351_));
 sky130_fd_sc_hd__nand2_1 _16261_ (.A(net447),
    .B(net1028),
    .Y(_08352_));
 sky130_fd_sc_hd__nand2_1 _16262_ (.A(net521),
    .B(net446),
    .Y(_08353_));
 sky130_fd_sc_hd__xnor2_1 _16263_ (.A(_08352_),
    .B(_08353_),
    .Y(_08354_));
 sky130_fd_sc_hd__xnor2_1 _16264_ (.A(_08351_),
    .B(_08354_),
    .Y(_08355_));
 sky130_fd_sc_hd__nand2_1 _16265_ (.A(net453),
    .B(net1029),
    .Y(_08356_));
 sky130_fd_sc_hd__nand2_1 _16266_ (.A(net449),
    .B(net516),
    .Y(_08357_));
 sky130_fd_sc_hd__nand2_1 _16267_ (.A(net456),
    .B(net510),
    .Y(_08358_));
 sky130_fd_sc_hd__xor2_1 _16268_ (.A(_08357_),
    .B(_08358_),
    .X(_08359_));
 sky130_fd_sc_hd__xnor2_1 _16269_ (.A(_08356_),
    .B(_08359_),
    .Y(_08360_));
 sky130_fd_sc_hd__xnor2_1 _16270_ (.A(_08355_),
    .B(_08360_),
    .Y(_08361_));
 sky130_fd_sc_hd__xnor2_2 _16271_ (.A(_08350_),
    .B(_08361_),
    .Y(_08362_));
 sky130_fd_sc_hd__a21bo_1 _16272_ (.A1(_08261_),
    .A2(_08266_),
    .B1_N(_08259_),
    .X(_08363_));
 sky130_fd_sc_hd__o21a_1 _16273_ (.A1(_08261_),
    .A2(_08266_),
    .B1(_08363_),
    .X(_08364_));
 sky130_fd_sc_hd__nand2_2 _16274_ (.A(net467),
    .B(net500),
    .Y(_08365_));
 sky130_fd_sc_hd__nand2_1 _16275_ (.A(net463),
    .B(net503),
    .Y(_08366_));
 sky130_fd_sc_hd__nand2_1 _16276_ (.A(net458),
    .B(net507),
    .Y(_08367_));
 sky130_fd_sc_hd__xnor2_1 _16277_ (.A(_08366_),
    .B(_08367_),
    .Y(_08368_));
 sky130_fd_sc_hd__xnor2_2 _16278_ (.A(_08365_),
    .B(_08368_),
    .Y(_08369_));
 sky130_fd_sc_hd__o21a_1 _16279_ (.A1(_08262_),
    .A2(_08264_),
    .B1(_08263_),
    .X(_08370_));
 sky130_fd_sc_hd__a21oi_2 _16280_ (.A1(_08262_),
    .A2(_08264_),
    .B1(_08370_),
    .Y(_08371_));
 sky130_fd_sc_hd__o21ba_1 _16281_ (.A1(_08272_),
    .A2(_08273_),
    .B1_N(_08271_),
    .X(_08372_));
 sky130_fd_sc_hd__a21oi_2 _16282_ (.A1(_08272_),
    .A2(_08273_),
    .B1(_08372_),
    .Y(_08373_));
 sky130_fd_sc_hd__xor2_1 _16283_ (.A(_08371_),
    .B(_08373_),
    .X(_08374_));
 sky130_fd_sc_hd__xnor2_2 _16284_ (.A(_08369_),
    .B(_08374_),
    .Y(_08375_));
 sky130_fd_sc_hd__xor2_1 _16285_ (.A(_08364_),
    .B(_08375_),
    .X(_08376_));
 sky130_fd_sc_hd__xnor2_2 _16286_ (.A(_08362_),
    .B(_08376_),
    .Y(_08377_));
 sky130_fd_sc_hd__a21bo_1 _16287_ (.A1(_08270_),
    .A2(_08281_),
    .B1_N(_08268_),
    .X(_08378_));
 sky130_fd_sc_hd__o21a_1 _16288_ (.A1(_08270_),
    .A2(_08281_),
    .B1(_08378_),
    .X(_08379_));
 sky130_fd_sc_hd__xnor2_1 _16289_ (.A(_08377_),
    .B(_08379_),
    .Y(_08380_));
 sky130_fd_sc_hd__xnor2_2 _16290_ (.A(_08348_),
    .B(_08380_),
    .Y(_08381_));
 sky130_fd_sc_hd__a21o_1 _16291_ (.A1(_08296_),
    .A2(_08300_),
    .B1(_08298_),
    .X(_08382_));
 sky130_fd_sc_hd__o21a_1 _16292_ (.A1(_08296_),
    .A2(_08300_),
    .B1(_08382_),
    .X(_08383_));
 sky130_fd_sc_hd__xnor2_1 _16293_ (.A(_08142_),
    .B(_08383_),
    .Y(_08384_));
 sky130_fd_sc_hd__a21bo_1 _16294_ (.A1(_08283_),
    .A2(_08302_),
    .B1_N(_08285_),
    .X(_08385_));
 sky130_fd_sc_hd__o21ai_2 _16295_ (.A1(_08283_),
    .A2(_08302_),
    .B1(_08385_),
    .Y(_08386_));
 sky130_fd_sc_hd__xnor2_1 _16296_ (.A(_08384_),
    .B(_08386_),
    .Y(_08387_));
 sky130_fd_sc_hd__xnor2_1 _16297_ (.A(_08381_),
    .B(_08387_),
    .Y(_08388_));
 sky130_fd_sc_hd__xnor2_1 _16298_ (.A(_08307_),
    .B(_08388_),
    .Y(_08389_));
 sky130_fd_sc_hd__xnor2_1 _16299_ (.A(_08334_),
    .B(_08389_),
    .Y(_08390_));
 sky130_fd_sc_hd__a21o_1 _16300_ (.A1(_08254_),
    .A2(_08311_),
    .B1(_08313_),
    .X(_08391_));
 sky130_fd_sc_hd__o21ai_1 _16301_ (.A1(_08254_),
    .A2(_08311_),
    .B1(_08391_),
    .Y(_08392_));
 sky130_fd_sc_hd__or2b_1 _16302_ (.A(_08390_),
    .B_N(_08392_),
    .X(_08393_));
 sky130_fd_sc_hd__and2b_1 _16303_ (.A_N(_08392_),
    .B(_08390_),
    .X(_08394_));
 sky130_fd_sc_hd__inv_2 _16304_ (.A(_08394_),
    .Y(_08395_));
 sky130_fd_sc_hd__nand2_1 _16305_ (.A(_08393_),
    .B(_08395_),
    .Y(_08396_));
 sky130_fd_sc_hd__a21oi_1 _16306_ (.A1(_08316_),
    .A2(_08330_),
    .B1(_08396_),
    .Y(_08397_));
 sky130_fd_sc_hd__and3_1 _16307_ (.A(_08316_),
    .B(_08330_),
    .C(_08396_),
    .X(_08398_));
 sky130_fd_sc_hd__or2_1 _16308_ (.A(_08397_),
    .B(_08398_),
    .X(_08399_));
 sky130_fd_sc_hd__a32o_1 _16309_ (.A1(net545),
    .A2(_08328_),
    .A3(_08329_),
    .B1(net548),
    .B2(_08399_),
    .X(_08400_));
 sky130_fd_sc_hd__mux2_1 _16310_ (.A0(\top0.pid_q.out[8] ),
    .A1(_08400_),
    .S(_07700_),
    .X(_08401_));
 sky130_fd_sc_hd__and2_1 _16311_ (.A(_07800_),
    .B(_08401_),
    .X(_08402_));
 sky130_fd_sc_hd__clkbuf_1 _16312_ (.A(_08402_),
    .X(_00141_));
 sky130_fd_sc_hd__clkbuf_2 _16313_ (.A(_05443_),
    .X(_08403_));
 sky130_fd_sc_hd__inv_2 _16314_ (.A(\top0.pid_q.curr_int[8] ),
    .Y(_08404_));
 sky130_fd_sc_hd__o21ba_1 _16315_ (.A1(_08404_),
    .A2(_08326_),
    .B1_N(\top0.pid_q.out[8] ),
    .X(_08405_));
 sky130_fd_sc_hd__a21o_1 _16316_ (.A1(_08404_),
    .A2(_08326_),
    .B1(_08405_),
    .X(_08406_));
 sky130_fd_sc_hd__xnor2_1 _16317_ (.A(\top0.pid_q.out[9] ),
    .B(\top0.pid_q.curr_int[9] ),
    .Y(_08407_));
 sky130_fd_sc_hd__nand2_1 _16318_ (.A(_08406_),
    .B(_08407_),
    .Y(_08408_));
 sky130_fd_sc_hd__or2_1 _16319_ (.A(_08406_),
    .B(_08407_),
    .X(_08409_));
 sky130_fd_sc_hd__a21o_1 _16320_ (.A1(_08316_),
    .A2(_08330_),
    .B1(_08394_),
    .X(_08410_));
 sky130_fd_sc_hd__nand2_1 _16321_ (.A(_08393_),
    .B(_08410_),
    .Y(_08411_));
 sky130_fd_sc_hd__o21ba_1 _16322_ (.A1(_08377_),
    .A2(_08379_),
    .B1_N(_08348_),
    .X(_08412_));
 sky130_fd_sc_hd__a21o_1 _16323_ (.A1(_08377_),
    .A2(_08379_),
    .B1(_08412_),
    .X(_08413_));
 sky130_fd_sc_hd__o21a_1 _16324_ (.A1(_08351_),
    .A2(_08353_),
    .B1(_08352_),
    .X(_08414_));
 sky130_fd_sc_hd__a21oi_2 _16325_ (.A1(_08351_),
    .A2(_08353_),
    .B1(_08414_),
    .Y(_08415_));
 sky130_fd_sc_hd__nand2_2 _16326_ (.A(_07230_),
    .B(net444),
    .Y(_08416_));
 sky130_fd_sc_hd__nand2_1 _16327_ (.A(net447),
    .B(net516),
    .Y(_08417_));
 sky130_fd_sc_hd__nand2_1 _16328_ (.A(net1028),
    .B(net446),
    .Y(_08418_));
 sky130_fd_sc_hd__xnor2_1 _16329_ (.A(_08417_),
    .B(_08418_),
    .Y(_08419_));
 sky130_fd_sc_hd__xnor2_2 _16330_ (.A(_08416_),
    .B(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__nand2_1 _16331_ (.A(net449),
    .B(net1029),
    .Y(_08421_));
 sky130_fd_sc_hd__nand2_1 _16332_ (.A(net456),
    .B(net507),
    .Y(_08422_));
 sky130_fd_sc_hd__nand2_1 _16333_ (.A(net453),
    .B(net510),
    .Y(_08423_));
 sky130_fd_sc_hd__xnor2_1 _16334_ (.A(_08422_),
    .B(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__xnor2_2 _16335_ (.A(_08421_),
    .B(_08424_),
    .Y(_08425_));
 sky130_fd_sc_hd__xor2_1 _16336_ (.A(_08420_),
    .B(_08425_),
    .X(_08426_));
 sky130_fd_sc_hd__xnor2_2 _16337_ (.A(_08415_),
    .B(_08426_),
    .Y(_08427_));
 sky130_fd_sc_hd__a21bo_1 _16338_ (.A1(_08350_),
    .A2(_08360_),
    .B1_N(_08355_),
    .X(_08428_));
 sky130_fd_sc_hd__o21a_1 _16339_ (.A1(_08350_),
    .A2(_08360_),
    .B1(_08428_),
    .X(_08429_));
 sky130_fd_sc_hd__nand2_2 _16340_ (.A(net466),
    .B(net497),
    .Y(_08430_));
 sky130_fd_sc_hd__nand2_1 _16341_ (.A(net458),
    .B(net503),
    .Y(_08431_));
 sky130_fd_sc_hd__nand2_1 _16342_ (.A(net463),
    .B(net501),
    .Y(_08432_));
 sky130_fd_sc_hd__xnor2_1 _16343_ (.A(_08431_),
    .B(_08432_),
    .Y(_08433_));
 sky130_fd_sc_hd__xnor2_2 _16344_ (.A(_08430_),
    .B(_08433_),
    .Y(_08434_));
 sky130_fd_sc_hd__o21a_1 _16345_ (.A1(_08356_),
    .A2(_08358_),
    .B1(_08357_),
    .X(_08435_));
 sky130_fd_sc_hd__a21oi_2 _16346_ (.A1(_08356_),
    .A2(_08358_),
    .B1(_08435_),
    .Y(_08436_));
 sky130_fd_sc_hd__o21a_1 _16347_ (.A1(_08365_),
    .A2(_08366_),
    .B1(_08367_),
    .X(_08437_));
 sky130_fd_sc_hd__a21oi_2 _16348_ (.A1(_08365_),
    .A2(_08366_),
    .B1(_08437_),
    .Y(_08438_));
 sky130_fd_sc_hd__xor2_1 _16349_ (.A(_08436_),
    .B(_08438_),
    .X(_08439_));
 sky130_fd_sc_hd__xnor2_2 _16350_ (.A(_08434_),
    .B(_08439_),
    .Y(_08440_));
 sky130_fd_sc_hd__xnor2_1 _16351_ (.A(_08429_),
    .B(_08440_),
    .Y(_08441_));
 sky130_fd_sc_hd__xnor2_2 _16352_ (.A(_08427_),
    .B(_08441_),
    .Y(_08442_));
 sky130_fd_sc_hd__a21bo_1 _16353_ (.A1(_08364_),
    .A2(_08375_),
    .B1_N(_08362_),
    .X(_08443_));
 sky130_fd_sc_hd__o21a_1 _16354_ (.A1(_08364_),
    .A2(_08375_),
    .B1(_08443_),
    .X(_08444_));
 sky130_fd_sc_hd__a21bo_1 _16355_ (.A1(_08371_),
    .A2(_08373_),
    .B1_N(_08369_),
    .X(_08445_));
 sky130_fd_sc_hd__o21ai_2 _16356_ (.A1(_08371_),
    .A2(_08373_),
    .B1(_08445_),
    .Y(_08446_));
 sky130_fd_sc_hd__or2_1 _16357_ (.A(_08048_),
    .B(_08340_),
    .X(_08447_));
 sky130_fd_sc_hd__or2b_1 _16358_ (.A(net476),
    .B_N(net473),
    .X(_08448_));
 sky130_fd_sc_hd__nand2_1 _16359_ (.A(_07493_),
    .B(_08448_),
    .Y(_08449_));
 sky130_fd_sc_hd__nand4_1 _16360_ (.A(net469),
    .B(_08141_),
    .C(_08048_),
    .D(_08449_),
    .Y(_08450_));
 sky130_fd_sc_hd__nand3_1 _16361_ (.A(net497),
    .B(_08447_),
    .C(_08450_),
    .Y(_08451_));
 sky130_fd_sc_hd__and4_1 _16362_ (.A(net468),
    .B(net473),
    .C(net476),
    .D(_08286_),
    .X(_08452_));
 sky130_fd_sc_hd__buf_2 _16363_ (.A(_08452_),
    .X(_08453_));
 sky130_fd_sc_hd__nor2_1 _16364_ (.A(_08451_),
    .B(_08453_),
    .Y(_08454_));
 sky130_fd_sc_hd__xnor2_1 _16365_ (.A(_08446_),
    .B(_08454_),
    .Y(_08455_));
 sky130_fd_sc_hd__nor2_1 _16366_ (.A(_08444_),
    .B(_08455_),
    .Y(_08456_));
 sky130_fd_sc_hd__nand2_1 _16367_ (.A(_08444_),
    .B(_08455_),
    .Y(_08457_));
 sky130_fd_sc_hd__or2b_1 _16368_ (.A(_08456_),
    .B_N(_08457_),
    .X(_08458_));
 sky130_fd_sc_hd__xnor2_1 _16369_ (.A(_08442_),
    .B(_08458_),
    .Y(_08459_));
 sky130_fd_sc_hd__o21a_1 _16370_ (.A1(_08339_),
    .A2(_08346_),
    .B1(_08337_),
    .X(_08460_));
 sky130_fd_sc_hd__a21o_1 _16371_ (.A1(_08339_),
    .A2(_08346_),
    .B1(_08460_),
    .X(_08461_));
 sky130_fd_sc_hd__xnor2_1 _16372_ (.A(_08142_),
    .B(_08461_),
    .Y(_08462_));
 sky130_fd_sc_hd__nand2_1 _16373_ (.A(_08459_),
    .B(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__nor2_1 _16374_ (.A(_08459_),
    .B(_08462_),
    .Y(_08464_));
 sky130_fd_sc_hd__inv_2 _16375_ (.A(_08464_),
    .Y(_08465_));
 sky130_fd_sc_hd__nand2_1 _16376_ (.A(_08463_),
    .B(_08465_),
    .Y(_08466_));
 sky130_fd_sc_hd__xnor2_2 _16377_ (.A(_08413_),
    .B(_08466_),
    .Y(_08467_));
 sky130_fd_sc_hd__inv_2 _16378_ (.A(_08386_),
    .Y(_08468_));
 sky130_fd_sc_hd__nand2_1 _16379_ (.A(_08383_),
    .B(_08381_),
    .Y(_08469_));
 sky130_fd_sc_hd__nor2_1 _16380_ (.A(_08383_),
    .B(_08381_),
    .Y(_08470_));
 sky130_fd_sc_hd__a21o_1 _16381_ (.A1(_08468_),
    .A2(_08469_),
    .B1(_08470_),
    .X(_08471_));
 sky130_fd_sc_hd__or4_1 _16382_ (.A(_08142_),
    .B(_08383_),
    .C(_08381_),
    .D(_08386_),
    .X(_08472_));
 sky130_fd_sc_hd__o221a_1 _16383_ (.A1(_08468_),
    .A2(_08469_),
    .B1(_08471_),
    .B2(_08312_),
    .C1(_08472_),
    .X(_08473_));
 sky130_fd_sc_hd__xnor2_2 _16384_ (.A(_08467_),
    .B(_08473_),
    .Y(_08474_));
 sky130_fd_sc_hd__inv_2 _16385_ (.A(_08388_),
    .Y(_08475_));
 sky130_fd_sc_hd__o21ba_1 _16386_ (.A1(_08334_),
    .A2(_08475_),
    .B1_N(_08307_),
    .X(_08476_));
 sky130_fd_sc_hd__a21oi_2 _16387_ (.A1(_08334_),
    .A2(_08475_),
    .B1(_08476_),
    .Y(_08477_));
 sky130_fd_sc_hd__xor2_1 _16388_ (.A(_08474_),
    .B(_08477_),
    .X(_08478_));
 sky130_fd_sc_hd__xnor2_2 _16389_ (.A(_08411_),
    .B(_08478_),
    .Y(_08479_));
 sky130_fd_sc_hd__a32o_1 _16390_ (.A1(net545),
    .A2(_08408_),
    .A3(_08409_),
    .B1(net549),
    .B2(_08479_),
    .X(_08480_));
 sky130_fd_sc_hd__mux2_1 _16391_ (.A0(\top0.pid_q.out[9] ),
    .A1(_08480_),
    .S(net13),
    .X(_08481_));
 sky130_fd_sc_hd__and2_1 _16392_ (.A(net1018),
    .B(_08481_),
    .X(_08482_));
 sky130_fd_sc_hd__clkbuf_1 _16393_ (.A(_08482_),
    .X(_00142_));
 sky130_fd_sc_hd__xor2_1 _16394_ (.A(\top0.pid_q.out[10] ),
    .B(\top0.pid_q.curr_int[10] ),
    .X(_08483_));
 sky130_fd_sc_hd__nor2_1 _16395_ (.A(\top0.pid_q.out[9] ),
    .B(\top0.pid_q.curr_int[9] ),
    .Y(_08484_));
 sky130_fd_sc_hd__nand2_1 _16396_ (.A(\top0.pid_q.out[9] ),
    .B(\top0.pid_q.curr_int[9] ),
    .Y(_08485_));
 sky130_fd_sc_hd__o21ai_2 _16397_ (.A1(_08406_),
    .A2(_08484_),
    .B1(_08485_),
    .Y(_08486_));
 sky130_fd_sc_hd__nand2_1 _16398_ (.A(_08483_),
    .B(_08486_),
    .Y(_08487_));
 sky130_fd_sc_hd__or2_1 _16399_ (.A(_08483_),
    .B(_08486_),
    .X(_08488_));
 sky130_fd_sc_hd__nand2_1 _16400_ (.A(_08474_),
    .B(_08477_),
    .Y(_08489_));
 sky130_fd_sc_hd__nor2_1 _16401_ (.A(_08474_),
    .B(_08477_),
    .Y(_08490_));
 sky130_fd_sc_hd__a31o_1 _16402_ (.A1(_08393_),
    .A2(_08410_),
    .A3(_08489_),
    .B1(_08490_),
    .X(_08491_));
 sky130_fd_sc_hd__a21oi_2 _16403_ (.A1(_08413_),
    .A2(_08463_),
    .B1(_08464_),
    .Y(_08492_));
 sky130_fd_sc_hd__nor2_1 _16404_ (.A(_08142_),
    .B(_08461_),
    .Y(_08493_));
 sky130_fd_sc_hd__o21a_1 _16405_ (.A1(_08416_),
    .A2(_08418_),
    .B1(_08417_),
    .X(_08494_));
 sky130_fd_sc_hd__a21oi_2 _16406_ (.A1(_08416_),
    .A2(_08418_),
    .B1(_08494_),
    .Y(_08495_));
 sky130_fd_sc_hd__nand2_1 _16407_ (.A(net450),
    .B(net510),
    .Y(_08496_));
 sky130_fd_sc_hd__nand2_1 _16408_ (.A(net456),
    .B(net503),
    .Y(_08497_));
 sky130_fd_sc_hd__nand2_1 _16409_ (.A(net452),
    .B(net506),
    .Y(_08498_));
 sky130_fd_sc_hd__xnor2_1 _16410_ (.A(_08497_),
    .B(_08498_),
    .Y(_08499_));
 sky130_fd_sc_hd__xnor2_2 _16411_ (.A(_08496_),
    .B(_08499_),
    .Y(_08500_));
 sky130_fd_sc_hd__nand2b_2 _16412_ (.A_N(net1028),
    .B(net444),
    .Y(_08501_));
 sky130_fd_sc_hd__nand2_1 _16413_ (.A(net447),
    .B(net1029),
    .Y(_08502_));
 sky130_fd_sc_hd__nand2_1 _16414_ (.A(net516),
    .B(net445),
    .Y(_08503_));
 sky130_fd_sc_hd__xnor2_1 _16415_ (.A(_08502_),
    .B(_08503_),
    .Y(_08504_));
 sky130_fd_sc_hd__xnor2_2 _16416_ (.A(_08501_),
    .B(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__xnor2_1 _16417_ (.A(_08500_),
    .B(_08505_),
    .Y(_08506_));
 sky130_fd_sc_hd__xnor2_2 _16418_ (.A(_08495_),
    .B(_08506_),
    .Y(_08507_));
 sky130_fd_sc_hd__o21ba_1 _16419_ (.A1(_08420_),
    .A2(_08425_),
    .B1_N(_08415_),
    .X(_08508_));
 sky130_fd_sc_hd__a21o_1 _16420_ (.A1(_08420_),
    .A2(_08425_),
    .B1(_08508_),
    .X(_08509_));
 sky130_fd_sc_hd__nand2_1 _16421_ (.A(net458),
    .B(net501),
    .Y(_08510_));
 sky130_fd_sc_hd__xor2_1 _16422_ (.A(net461),
    .B(net466),
    .X(_08511_));
 sky130_fd_sc_hd__nand2_1 _16423_ (.A(net498),
    .B(_08511_),
    .Y(_08512_));
 sky130_fd_sc_hd__xor2_1 _16424_ (.A(_08510_),
    .B(_08512_),
    .X(_08513_));
 sky130_fd_sc_hd__o21ai_1 _16425_ (.A1(_08422_),
    .A2(_08423_),
    .B1(_08421_),
    .Y(_08514_));
 sky130_fd_sc_hd__a21bo_1 _16426_ (.A1(_08422_),
    .A2(_08423_),
    .B1_N(_08514_),
    .X(_08515_));
 sky130_fd_sc_hd__o21ai_1 _16427_ (.A1(_08430_),
    .A2(_08432_),
    .B1(_08431_),
    .Y(_08516_));
 sky130_fd_sc_hd__a21bo_1 _16428_ (.A1(_08430_),
    .A2(_08432_),
    .B1_N(_08516_),
    .X(_08517_));
 sky130_fd_sc_hd__xnor2_1 _16429_ (.A(_08515_),
    .B(_08517_),
    .Y(_08518_));
 sky130_fd_sc_hd__xnor2_1 _16430_ (.A(_08513_),
    .B(_08518_),
    .Y(_08519_));
 sky130_fd_sc_hd__xnor2_1 _16431_ (.A(_08509_),
    .B(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__xnor2_2 _16432_ (.A(_08507_),
    .B(_08520_),
    .Y(_08521_));
 sky130_fd_sc_hd__a21bo_1 _16433_ (.A1(_08429_),
    .A2(_08440_),
    .B1_N(_08427_),
    .X(_08522_));
 sky130_fd_sc_hd__o21a_1 _16434_ (.A1(_08429_),
    .A2(_08440_),
    .B1(_08522_),
    .X(_08523_));
 sky130_fd_sc_hd__a21bo_1 _16435_ (.A1(_08436_),
    .A2(_08438_),
    .B1_N(_08434_),
    .X(_08524_));
 sky130_fd_sc_hd__o21a_1 _16436_ (.A1(_08436_),
    .A2(_08438_),
    .B1(_08524_),
    .X(_08525_));
 sky130_fd_sc_hd__nand2_2 _16437_ (.A(net498),
    .B(_08447_),
    .Y(_08526_));
 sky130_fd_sc_hd__nor2_4 _16438_ (.A(_08453_),
    .B(_08526_),
    .Y(_08527_));
 sky130_fd_sc_hd__xnor2_1 _16439_ (.A(_08525_),
    .B(_08527_),
    .Y(_08528_));
 sky130_fd_sc_hd__and2b_1 _16440_ (.A_N(_08523_),
    .B(_08528_),
    .X(_08529_));
 sky130_fd_sc_hd__or2b_1 _16441_ (.A(_08528_),
    .B_N(_08523_),
    .X(_08530_));
 sky130_fd_sc_hd__or2b_1 _16442_ (.A(_08529_),
    .B_N(_08530_),
    .X(_08531_));
 sky130_fd_sc_hd__xnor2_2 _16443_ (.A(_08521_),
    .B(_08531_),
    .Y(_08532_));
 sky130_fd_sc_hd__a21o_1 _16444_ (.A1(_08442_),
    .A2(_08457_),
    .B1(_08456_),
    .X(_08533_));
 sky130_fd_sc_hd__nand4_2 _16445_ (.A(net468),
    .B(net473),
    .C(net476),
    .D(_08286_),
    .Y(_08534_));
 sky130_fd_sc_hd__a21oi_1 _16446_ (.A1(_08446_),
    .A2(_08534_),
    .B1(_08451_),
    .Y(_08535_));
 sky130_fd_sc_hd__xnor2_1 _16447_ (.A(_08220_),
    .B(_08535_),
    .Y(_08536_));
 sky130_fd_sc_hd__and2_1 _16448_ (.A(_08533_),
    .B(_08536_),
    .X(_08537_));
 sky130_fd_sc_hd__or2_1 _16449_ (.A(_08533_),
    .B(_08536_),
    .X(_08538_));
 sky130_fd_sc_hd__or2b_1 _16450_ (.A(_08537_),
    .B_N(_08538_),
    .X(_08539_));
 sky130_fd_sc_hd__xnor2_2 _16451_ (.A(_08532_),
    .B(_08539_),
    .Y(_08540_));
 sky130_fd_sc_hd__xnor2_1 _16452_ (.A(_08493_),
    .B(_08540_),
    .Y(_08541_));
 sky130_fd_sc_hd__xnor2_2 _16453_ (.A(_08492_),
    .B(_08541_),
    .Y(_08542_));
 sky130_fd_sc_hd__inv_2 _16454_ (.A(_08542_),
    .Y(_08543_));
 sky130_fd_sc_hd__nor2_1 _16455_ (.A(_08467_),
    .B(_08470_),
    .Y(_08544_));
 sky130_fd_sc_hd__o2bb2a_1 _16456_ (.A1_N(_08467_),
    .A2_N(_08469_),
    .B1(_08544_),
    .B2(_08386_),
    .X(_08545_));
 sky130_fd_sc_hd__o2bb2a_1 _16457_ (.A1_N(_08467_),
    .A2_N(_08471_),
    .B1(_08545_),
    .B2(_08142_),
    .X(_08546_));
 sky130_fd_sc_hd__nor2_1 _16458_ (.A(_08543_),
    .B(_08546_),
    .Y(_08547_));
 sky130_fd_sc_hd__nand2_1 _16459_ (.A(_08543_),
    .B(_08546_),
    .Y(_08548_));
 sky130_fd_sc_hd__or2b_1 _16460_ (.A(_08547_),
    .B_N(_08548_),
    .X(_08549_));
 sky130_fd_sc_hd__xnor2_2 _16461_ (.A(_08491_),
    .B(_08549_),
    .Y(_08550_));
 sky130_fd_sc_hd__a32o_1 _16462_ (.A1(net545),
    .A2(_08487_),
    .A3(_08488_),
    .B1(net549),
    .B2(_08550_),
    .X(_08551_));
 sky130_fd_sc_hd__mux2_1 _16463_ (.A0(\top0.pid_q.out[10] ),
    .A1(_08551_),
    .S(net13),
    .X(_08552_));
 sky130_fd_sc_hd__and2_1 _16464_ (.A(net1018),
    .B(_08552_),
    .X(_08553_));
 sky130_fd_sc_hd__clkbuf_1 _16465_ (.A(_08553_),
    .X(_00143_));
 sky130_fd_sc_hd__nand2_2 _16466_ (.A(net455),
    .B(net500),
    .Y(_08554_));
 sky130_fd_sc_hd__nand2_1 _16467_ (.A(net452),
    .B(net503),
    .Y(_08555_));
 sky130_fd_sc_hd__nand2_1 _16468_ (.A(net450),
    .B(net506),
    .Y(_08556_));
 sky130_fd_sc_hd__xnor2_1 _16469_ (.A(_08555_),
    .B(_08556_),
    .Y(_08557_));
 sky130_fd_sc_hd__xnor2_2 _16470_ (.A(_08554_),
    .B(_08557_),
    .Y(_08558_));
 sky130_fd_sc_hd__o21a_1 _16471_ (.A1(_08501_),
    .A2(_08503_),
    .B1(_08502_),
    .X(_08559_));
 sky130_fd_sc_hd__a21oi_2 _16472_ (.A1(_08501_),
    .A2(_08503_),
    .B1(_08559_),
    .Y(_08560_));
 sky130_fd_sc_hd__nand2b_2 _16473_ (.A_N(net516),
    .B(\top0.pid_q.mult0.b[15] ),
    .Y(_08561_));
 sky130_fd_sc_hd__nand2_1 _16474_ (.A(net1029),
    .B(\top0.pid_q.mult0.b[14] ),
    .Y(_08562_));
 sky130_fd_sc_hd__nand2_1 _16475_ (.A(net447),
    .B(net510),
    .Y(_08563_));
 sky130_fd_sc_hd__xor2_1 _16476_ (.A(_08562_),
    .B(_08563_),
    .X(_08564_));
 sky130_fd_sc_hd__xnor2_2 _16477_ (.A(_08561_),
    .B(_08564_),
    .Y(_08565_));
 sky130_fd_sc_hd__xnor2_1 _16478_ (.A(_08560_),
    .B(_08565_),
    .Y(_08566_));
 sky130_fd_sc_hd__xnor2_2 _16479_ (.A(_08558_),
    .B(_08566_),
    .Y(_08567_));
 sky130_fd_sc_hd__o21ba_1 _16480_ (.A1(_08500_),
    .A2(_08505_),
    .B1_N(_08495_),
    .X(_08568_));
 sky130_fd_sc_hd__a21o_1 _16481_ (.A1(_08500_),
    .A2(_08505_),
    .B1(_08568_),
    .X(_08569_));
 sky130_fd_sc_hd__o21ai_1 _16482_ (.A1(_08497_),
    .A2(_08498_),
    .B1(_08496_),
    .Y(_08570_));
 sky130_fd_sc_hd__a21boi_2 _16483_ (.A1(_08497_),
    .A2(_08498_),
    .B1_N(_08570_),
    .Y(_08571_));
 sky130_fd_sc_hd__o21a_1 _16484_ (.A1(net466),
    .A2(_08141_),
    .B1(net461),
    .X(_08572_));
 sky130_fd_sc_hd__a21o_1 _16485_ (.A1(net466),
    .A2(_08141_),
    .B1(_08572_),
    .X(_08573_));
 sky130_fd_sc_hd__or3_1 _16486_ (.A(net458),
    .B(net461),
    .C(net466),
    .X(_08574_));
 sky130_fd_sc_hd__nand2_1 _16487_ (.A(net497),
    .B(_08574_),
    .Y(_08575_));
 sky130_fd_sc_hd__a21oi_1 _16488_ (.A1(net459),
    .A2(_08573_),
    .B1(_08575_),
    .Y(_08576_));
 sky130_fd_sc_hd__xnor2_2 _16489_ (.A(_08571_),
    .B(_08576_),
    .Y(_08577_));
 sky130_fd_sc_hd__xor2_1 _16490_ (.A(_08569_),
    .B(_08577_),
    .X(_08578_));
 sky130_fd_sc_hd__xnor2_2 _16491_ (.A(_08567_),
    .B(_08578_),
    .Y(_08579_));
 sky130_fd_sc_hd__inv_2 _16492_ (.A(_08519_),
    .Y(_08580_));
 sky130_fd_sc_hd__o21ba_1 _16493_ (.A1(_08509_),
    .A2(_08580_),
    .B1_N(_08507_),
    .X(_08581_));
 sky130_fd_sc_hd__a21oi_2 _16494_ (.A1(_08509_),
    .A2(_08580_),
    .B1(_08581_),
    .Y(_08582_));
 sky130_fd_sc_hd__a21bo_1 _16495_ (.A1(_08515_),
    .A2(_08517_),
    .B1_N(_08513_),
    .X(_08583_));
 sky130_fd_sc_hd__o21a_1 _16496_ (.A1(_08515_),
    .A2(_08517_),
    .B1(_08583_),
    .X(_08584_));
 sky130_fd_sc_hd__xnor2_2 _16497_ (.A(_08527_),
    .B(_08584_),
    .Y(_08585_));
 sky130_fd_sc_hd__xor2_1 _16498_ (.A(_08582_),
    .B(_08585_),
    .X(_08586_));
 sky130_fd_sc_hd__xnor2_2 _16499_ (.A(_08579_),
    .B(_08586_),
    .Y(_08587_));
 sky130_fd_sc_hd__a21o_1 _16500_ (.A1(_08521_),
    .A2(_08530_),
    .B1(_08529_),
    .X(_08588_));
 sky130_fd_sc_hd__o21ba_1 _16501_ (.A1(_08453_),
    .A2(_08525_),
    .B1_N(_08526_),
    .X(_08589_));
 sky130_fd_sc_hd__xnor2_2 _16502_ (.A(_08312_),
    .B(_08589_),
    .Y(_08590_));
 sky130_fd_sc_hd__xnor2_1 _16503_ (.A(_08588_),
    .B(_08590_),
    .Y(_08591_));
 sky130_fd_sc_hd__xnor2_2 _16504_ (.A(_08587_),
    .B(_08591_),
    .Y(_08592_));
 sky130_fd_sc_hd__o21a_1 _16505_ (.A1(_08532_),
    .A2(_08537_),
    .B1(_08538_),
    .X(_08593_));
 sky130_fd_sc_hd__nand2_1 _16506_ (.A(_08312_),
    .B(_08535_),
    .Y(_08594_));
 sky130_fd_sc_hd__xnor2_1 _16507_ (.A(_08593_),
    .B(_08594_),
    .Y(_08595_));
 sky130_fd_sc_hd__xnor2_1 _16508_ (.A(_08592_),
    .B(_08595_),
    .Y(_08596_));
 sky130_fd_sc_hd__a21bo_1 _16509_ (.A1(_08492_),
    .A2(_08540_),
    .B1_N(_08493_),
    .X(_08597_));
 sky130_fd_sc_hd__o21a_1 _16510_ (.A1(_08492_),
    .A2(_08540_),
    .B1(_08597_),
    .X(_08598_));
 sky130_fd_sc_hd__nand2_1 _16511_ (.A(_08596_),
    .B(_08598_),
    .Y(_08599_));
 sky130_fd_sc_hd__inv_2 _16512_ (.A(_08599_),
    .Y(_08600_));
 sky130_fd_sc_hd__nor2_1 _16513_ (.A(_08596_),
    .B(_08598_),
    .Y(_08601_));
 sky130_fd_sc_hd__or2_1 _16514_ (.A(_08600_),
    .B(_08601_),
    .X(_08602_));
 sky130_fd_sc_hd__a31o_1 _16515_ (.A1(_08316_),
    .A2(_08330_),
    .A3(_08393_),
    .B1(_08394_),
    .X(_08603_));
 sky130_fd_sc_hd__a21oi_1 _16516_ (.A1(_08489_),
    .A2(_08603_),
    .B1(_08490_),
    .Y(_08604_));
 sky130_fd_sc_hd__nor2_1 _16517_ (.A(_08546_),
    .B(_08604_),
    .Y(_08605_));
 sky130_fd_sc_hd__a21o_1 _16518_ (.A1(_08393_),
    .A2(_08410_),
    .B1(_08490_),
    .X(_08606_));
 sky130_fd_sc_hd__a21bo_1 _16519_ (.A1(_08489_),
    .A2(_08606_),
    .B1_N(_08546_),
    .X(_08607_));
 sky130_fd_sc_hd__o21ai_2 _16520_ (.A1(_08542_),
    .A2(_08605_),
    .B1(_08607_),
    .Y(_08608_));
 sky130_fd_sc_hd__xnor2_2 _16521_ (.A(_08602_),
    .B(_08608_),
    .Y(_08609_));
 sky130_fd_sc_hd__nor2_1 _16522_ (.A(_07701_),
    .B(_08609_),
    .Y(_08610_));
 sky130_fd_sc_hd__nor2_1 _16523_ (.A(\top0.pid_q.out[11] ),
    .B(_07704_),
    .Y(_08611_));
 sky130_fd_sc_hd__and2_1 _16524_ (.A(\top0.pid_q.out[10] ),
    .B(\top0.pid_q.curr_int[10] ),
    .X(_08612_));
 sky130_fd_sc_hd__or2_1 _16525_ (.A(\top0.pid_q.out[10] ),
    .B(\top0.pid_q.curr_int[10] ),
    .X(_08613_));
 sky130_fd_sc_hd__o21ai_2 _16526_ (.A1(_08486_),
    .A2(_08612_),
    .B1(_08613_),
    .Y(_08614_));
 sky130_fd_sc_hd__xnor2_1 _16527_ (.A(\top0.pid_q.curr_int[11] ),
    .B(_08614_),
    .Y(_08615_));
 sky130_fd_sc_hd__mux2_1 _16528_ (.A0(\top0.pid_q.out[11] ),
    .A1(_08611_),
    .S(_08615_),
    .X(_08616_));
 sky130_fd_sc_hd__a22o_1 _16529_ (.A1(\top0.pid_q.out[11] ),
    .A2(_07705_),
    .B1(_08616_),
    .B2(net544),
    .X(_08617_));
 sky130_fd_sc_hd__o21a_1 _16530_ (.A1(_08610_),
    .A2(_08617_),
    .B1(_07710_),
    .X(_00144_));
 sky130_fd_sc_hd__nor2_1 _16531_ (.A(\top0.pid_q.out[12] ),
    .B(\top0.pid_q.curr_int[12] ),
    .Y(_08618_));
 sky130_fd_sc_hd__nand2_1 _16532_ (.A(\top0.pid_q.out[12] ),
    .B(\top0.pid_q.curr_int[12] ),
    .Y(_08619_));
 sky130_fd_sc_hd__a21bo_1 _16533_ (.A1(net13),
    .A2(_08618_),
    .B1_N(_08619_),
    .X(_08620_));
 sky130_fd_sc_hd__inv_2 _16534_ (.A(\top0.pid_q.curr_int[12] ),
    .Y(_08621_));
 sky130_fd_sc_hd__nor2_1 _16535_ (.A(_08621_),
    .B(_07703_),
    .Y(_08622_));
 sky130_fd_sc_hd__mux2_1 _16536_ (.A0(_08622_),
    .A1(_08621_),
    .S(\top0.pid_q.out[12] ),
    .X(_08623_));
 sky130_fd_sc_hd__inv_2 _16537_ (.A(\top0.pid_q.curr_int[11] ),
    .Y(_08624_));
 sky130_fd_sc_hd__a21bo_1 _16538_ (.A1(_08624_),
    .A2(_08614_),
    .B1_N(\top0.pid_q.out[11] ),
    .X(_08625_));
 sky130_fd_sc_hd__o21a_1 _16539_ (.A1(_08624_),
    .A2(_08614_),
    .B1(_08625_),
    .X(_08626_));
 sky130_fd_sc_hd__mux2_1 _16540_ (.A0(_08620_),
    .A1(_08623_),
    .S(_08626_),
    .X(_08627_));
 sky130_fd_sc_hd__o21a_1 _16541_ (.A1(_08567_),
    .A2(_08577_),
    .B1(_08569_),
    .X(_08628_));
 sky130_fd_sc_hd__a21o_1 _16542_ (.A1(_08567_),
    .A2(_08577_),
    .B1(_08628_),
    .X(_08629_));
 sky130_fd_sc_hd__nand2b_2 _16543_ (.A_N(net1029),
    .B(net444),
    .Y(_08630_));
 sky130_fd_sc_hd__nand2_1 _16544_ (.A(net510),
    .B(net445),
    .Y(_08631_));
 sky130_fd_sc_hd__nand2_1 _16545_ (.A(net447),
    .B(net507),
    .Y(_08632_));
 sky130_fd_sc_hd__xnor2_1 _16546_ (.A(_08631_),
    .B(_08632_),
    .Y(_08633_));
 sky130_fd_sc_hd__xnor2_2 _16547_ (.A(_08630_),
    .B(_08633_),
    .Y(_08634_));
 sky130_fd_sc_hd__o21a_1 _16548_ (.A1(_08561_),
    .A2(_08562_),
    .B1(_08563_),
    .X(_08635_));
 sky130_fd_sc_hd__a21oi_2 _16549_ (.A1(_08561_),
    .A2(_08562_),
    .B1(_08635_),
    .Y(_08636_));
 sky130_fd_sc_hd__nand2_2 _16550_ (.A(net456),
    .B(net497),
    .Y(_08637_));
 sky130_fd_sc_hd__nand2_1 _16551_ (.A(net450),
    .B(net503),
    .Y(_08638_));
 sky130_fd_sc_hd__nand2_1 _16552_ (.A(net452),
    .B(net501),
    .Y(_08639_));
 sky130_fd_sc_hd__xor2_1 _16553_ (.A(_08638_),
    .B(_08639_),
    .X(_08640_));
 sky130_fd_sc_hd__xnor2_2 _16554_ (.A(_08637_),
    .B(_08640_),
    .Y(_08641_));
 sky130_fd_sc_hd__xnor2_1 _16555_ (.A(_08636_),
    .B(_08641_),
    .Y(_08642_));
 sky130_fd_sc_hd__xnor2_2 _16556_ (.A(_08634_),
    .B(_08642_),
    .Y(_08643_));
 sky130_fd_sc_hd__a21bo_1 _16557_ (.A1(_08560_),
    .A2(_08565_),
    .B1_N(_08558_),
    .X(_08644_));
 sky130_fd_sc_hd__o21a_1 _16558_ (.A1(_08560_),
    .A2(_08565_),
    .B1(_08644_),
    .X(_08645_));
 sky130_fd_sc_hd__o21a_1 _16559_ (.A1(_08554_),
    .A2(_08555_),
    .B1(_08556_),
    .X(_08646_));
 sky130_fd_sc_hd__a21o_1 _16560_ (.A1(_08554_),
    .A2(_08555_),
    .B1(_08646_),
    .X(_08647_));
 sky130_fd_sc_hd__a21oi_4 _16561_ (.A1(net458),
    .A2(_07213_),
    .B1(_08575_),
    .Y(_08648_));
 sky130_fd_sc_hd__xnor2_1 _16562_ (.A(_08647_),
    .B(_08648_),
    .Y(_08649_));
 sky130_fd_sc_hd__nor2_1 _16563_ (.A(_08645_),
    .B(_08649_),
    .Y(_08650_));
 sky130_fd_sc_hd__nand2_1 _16564_ (.A(_08645_),
    .B(_08649_),
    .Y(_08651_));
 sky130_fd_sc_hd__and2b_1 _16565_ (.A_N(_08650_),
    .B(_08651_),
    .X(_08652_));
 sky130_fd_sc_hd__xor2_2 _16566_ (.A(_08643_),
    .B(_08652_),
    .X(_08653_));
 sky130_fd_sc_hd__nor2_1 _16567_ (.A(net461),
    .B(net466),
    .Y(_08654_));
 sky130_fd_sc_hd__or3b_1 _16568_ (.A(net501),
    .B(_08654_),
    .C_N(net459),
    .X(_08655_));
 sky130_fd_sc_hd__a32o_1 _16569_ (.A1(_08571_),
    .A2(_08574_),
    .A3(_08655_),
    .B1(_07213_),
    .B2(net459),
    .X(_08656_));
 sky130_fd_sc_hd__nand2_1 _16570_ (.A(net497),
    .B(_08656_),
    .Y(_08657_));
 sky130_fd_sc_hd__xor2_2 _16571_ (.A(_08527_),
    .B(_08657_),
    .X(_08658_));
 sky130_fd_sc_hd__xnor2_1 _16572_ (.A(_08653_),
    .B(_08658_),
    .Y(_08659_));
 sky130_fd_sc_hd__xnor2_2 _16573_ (.A(_08629_),
    .B(_08659_),
    .Y(_08660_));
 sky130_fd_sc_hd__a21o_1 _16574_ (.A1(_08582_),
    .A2(_08585_),
    .B1(_08579_),
    .X(_08661_));
 sky130_fd_sc_hd__o21ai_2 _16575_ (.A1(_08582_),
    .A2(_08585_),
    .B1(_08661_),
    .Y(_08662_));
 sky130_fd_sc_hd__o21ai_1 _16576_ (.A1(_08526_),
    .A2(_08584_),
    .B1(_08534_),
    .Y(_08663_));
 sky130_fd_sc_hd__nand2_1 _16577_ (.A(_08312_),
    .B(_08663_),
    .Y(_08664_));
 sky130_fd_sc_hd__or2_1 _16578_ (.A(_08312_),
    .B(_08663_),
    .X(_08665_));
 sky130_fd_sc_hd__nand2_1 _16579_ (.A(_08664_),
    .B(_08665_),
    .Y(_08666_));
 sky130_fd_sc_hd__xor2_1 _16580_ (.A(_08662_),
    .B(_08666_),
    .X(_08667_));
 sky130_fd_sc_hd__xnor2_2 _16581_ (.A(_08660_),
    .B(_08667_),
    .Y(_08668_));
 sky130_fd_sc_hd__o21a_1 _16582_ (.A1(_08588_),
    .A2(_08590_),
    .B1(_08587_),
    .X(_08669_));
 sky130_fd_sc_hd__a21oi_2 _16583_ (.A1(_08588_),
    .A2(_08590_),
    .B1(_08669_),
    .Y(_08670_));
 sky130_fd_sc_hd__nand2_1 _16584_ (.A(_08312_),
    .B(_08589_),
    .Y(_08671_));
 sky130_fd_sc_hd__xor2_1 _16585_ (.A(_08670_),
    .B(_08671_),
    .X(_08672_));
 sky130_fd_sc_hd__xnor2_1 _16586_ (.A(_08668_),
    .B(_08672_),
    .Y(_08673_));
 sky130_fd_sc_hd__a21oi_1 _16587_ (.A1(_08593_),
    .A2(_08592_),
    .B1(_08594_),
    .Y(_08674_));
 sky130_fd_sc_hd__nor2_1 _16588_ (.A(_08593_),
    .B(_08592_),
    .Y(_08675_));
 sky130_fd_sc_hd__or3_1 _16589_ (.A(_08673_),
    .B(_08674_),
    .C(_08675_),
    .X(_08676_));
 sky130_fd_sc_hd__o21ai_2 _16590_ (.A1(_08674_),
    .A2(_08675_),
    .B1(_08673_),
    .Y(_08677_));
 sky130_fd_sc_hd__nand2_1 _16591_ (.A(_08676_),
    .B(_08677_),
    .Y(_08678_));
 sky130_fd_sc_hd__mux2_1 _16592_ (.A0(_08600_),
    .A1(_08601_),
    .S(_08678_),
    .X(_08679_));
 sky130_fd_sc_hd__and3_1 _16593_ (.A(net549),
    .B(net13),
    .C(_08679_),
    .X(_08680_));
 sky130_fd_sc_hd__a221o_1 _16594_ (.A1(\top0.pid_q.out[12] ),
    .A2(_07705_),
    .B1(_08627_),
    .B2(net544),
    .C1(_08680_),
    .X(_08681_));
 sky130_fd_sc_hd__or2_1 _16595_ (.A(_08601_),
    .B(_08678_),
    .X(_08682_));
 sky130_fd_sc_hd__nand2_1 _16596_ (.A(_08599_),
    .B(_08678_),
    .Y(_08683_));
 sky130_fd_sc_hd__a21o_1 _16597_ (.A1(_08542_),
    .A2(_08607_),
    .B1(_08605_),
    .X(_08684_));
 sky130_fd_sc_hd__mux2_2 _16598_ (.A0(_08682_),
    .A1(_08683_),
    .S(_08684_),
    .X(_08685_));
 sky130_fd_sc_hd__nor2_1 _16599_ (.A(_07701_),
    .B(_08685_),
    .Y(_08686_));
 sky130_fd_sc_hd__o21a_1 _16600_ (.A1(_08681_),
    .A2(_08686_),
    .B1(_07710_),
    .X(_00145_));
 sky130_fd_sc_hd__a21oi_2 _16601_ (.A1(_08491_),
    .A2(_08548_),
    .B1(_08547_),
    .Y(_08687_));
 sky130_fd_sc_hd__nand2_1 _16602_ (.A(_08599_),
    .B(_08676_),
    .Y(_08688_));
 sky130_fd_sc_hd__nand2_1 _16603_ (.A(_08601_),
    .B(_08676_),
    .Y(_08689_));
 sky130_fd_sc_hd__o211ai_4 _16604_ (.A1(_08687_),
    .A2(_08688_),
    .B1(_08689_),
    .C1(_08677_),
    .Y(_08690_));
 sky130_fd_sc_hd__o21a_1 _16605_ (.A1(_08653_),
    .A2(_08658_),
    .B1(_08629_),
    .X(_08691_));
 sky130_fd_sc_hd__a21oi_2 _16606_ (.A1(_08653_),
    .A2(_08658_),
    .B1(_08691_),
    .Y(_08692_));
 sky130_fd_sc_hd__a21oi_1 _16607_ (.A1(_08534_),
    .A2(_08657_),
    .B1(_08526_),
    .Y(_08693_));
 sky130_fd_sc_hd__xnor2_1 _16608_ (.A(_08312_),
    .B(_08693_),
    .Y(_08694_));
 sky130_fd_sc_hd__nand2_1 _16609_ (.A(net449),
    .B(net500),
    .Y(_08695_));
 sky130_fd_sc_hd__xor2_1 _16610_ (.A(net452),
    .B(net455),
    .X(_08696_));
 sky130_fd_sc_hd__nand2_1 _16611_ (.A(net498),
    .B(_08696_),
    .Y(_08697_));
 sky130_fd_sc_hd__xor2_1 _16612_ (.A(_08695_),
    .B(_08697_),
    .X(_08698_));
 sky130_fd_sc_hd__o21a_1 _16613_ (.A1(_08630_),
    .A2(_08631_),
    .B1(_08632_),
    .X(_08699_));
 sky130_fd_sc_hd__a21oi_2 _16614_ (.A1(_08630_),
    .A2(_08631_),
    .B1(_08699_),
    .Y(_08700_));
 sky130_fd_sc_hd__nand2b_1 _16615_ (.A_N(net510),
    .B(net444),
    .Y(_08701_));
 sky130_fd_sc_hd__nand2_1 _16616_ (.A(net507),
    .B(net445),
    .Y(_08702_));
 sky130_fd_sc_hd__nand2_1 _16617_ (.A(net447),
    .B(net504),
    .Y(_08703_));
 sky130_fd_sc_hd__xor2_1 _16618_ (.A(_08702_),
    .B(_08703_),
    .X(_08704_));
 sky130_fd_sc_hd__xnor2_1 _16619_ (.A(_08701_),
    .B(_08704_),
    .Y(_08705_));
 sky130_fd_sc_hd__xor2_1 _16620_ (.A(_08700_),
    .B(_08705_),
    .X(_08706_));
 sky130_fd_sc_hd__xnor2_1 _16621_ (.A(_08698_),
    .B(_08706_),
    .Y(_08707_));
 sky130_fd_sc_hd__a21bo_1 _16622_ (.A1(_08636_),
    .A2(_08641_),
    .B1_N(_08634_),
    .X(_08708_));
 sky130_fd_sc_hd__o21a_1 _16623_ (.A1(_08636_),
    .A2(_08641_),
    .B1(_08708_),
    .X(_08709_));
 sky130_fd_sc_hd__o21a_1 _16624_ (.A1(_08637_),
    .A2(_08639_),
    .B1(_08638_),
    .X(_08710_));
 sky130_fd_sc_hd__a21oi_2 _16625_ (.A1(_08637_),
    .A2(_08639_),
    .B1(_08710_),
    .Y(_08711_));
 sky130_fd_sc_hd__xor2_1 _16626_ (.A(_08648_),
    .B(_08711_),
    .X(_08712_));
 sky130_fd_sc_hd__nor2_1 _16627_ (.A(_08709_),
    .B(_08712_),
    .Y(_08713_));
 sky130_fd_sc_hd__nand2_1 _16628_ (.A(_08709_),
    .B(_08712_),
    .Y(_08714_));
 sky130_fd_sc_hd__or2b_1 _16629_ (.A(_08713_),
    .B_N(_08714_),
    .X(_08715_));
 sky130_fd_sc_hd__xnor2_1 _16630_ (.A(_08707_),
    .B(_08715_),
    .Y(_08716_));
 sky130_fd_sc_hd__a21o_1 _16631_ (.A1(_08643_),
    .A2(_08651_),
    .B1(_08650_),
    .X(_08717_));
 sky130_fd_sc_hd__nand2_1 _16632_ (.A(net461),
    .B(net466),
    .Y(_08718_));
 sky130_fd_sc_hd__nand2_1 _16633_ (.A(_08718_),
    .B(_08647_),
    .Y(_08719_));
 sky130_fd_sc_hd__a2bb2o_1 _16634_ (.A1_N(_08654_),
    .A2_N(_08647_),
    .B1(_08719_),
    .B2(net459),
    .X(_08720_));
 sky130_fd_sc_hd__and2_1 _16635_ (.A(net498),
    .B(_08720_),
    .X(_08721_));
 sky130_fd_sc_hd__xnor2_2 _16636_ (.A(_08527_),
    .B(_08721_),
    .Y(_08722_));
 sky130_fd_sc_hd__xnor2_1 _16637_ (.A(_08717_),
    .B(_08722_),
    .Y(_08723_));
 sky130_fd_sc_hd__xnor2_1 _16638_ (.A(_08716_),
    .B(_08723_),
    .Y(_08724_));
 sky130_fd_sc_hd__nand2_1 _16639_ (.A(_08694_),
    .B(_08724_),
    .Y(_08725_));
 sky130_fd_sc_hd__or2_1 _16640_ (.A(_08694_),
    .B(_08724_),
    .X(_08726_));
 sky130_fd_sc_hd__nand2_1 _16641_ (.A(_08725_),
    .B(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__xnor2_2 _16642_ (.A(_08692_),
    .B(_08727_),
    .Y(_08728_));
 sky130_fd_sc_hd__a21o_1 _16643_ (.A1(_08662_),
    .A2(_08666_),
    .B1(_08660_),
    .X(_08729_));
 sky130_fd_sc_hd__o21ai_2 _16644_ (.A1(_08662_),
    .A2(_08666_),
    .B1(_08729_),
    .Y(_08730_));
 sky130_fd_sc_hd__xnor2_1 _16645_ (.A(_08664_),
    .B(_08730_),
    .Y(_08731_));
 sky130_fd_sc_hd__xnor2_1 _16646_ (.A(_08728_),
    .B(_08731_),
    .Y(_08732_));
 sky130_fd_sc_hd__a21bo_1 _16647_ (.A1(_08670_),
    .A2(_08668_),
    .B1_N(_08671_),
    .X(_08733_));
 sky130_fd_sc_hd__o21ai_1 _16648_ (.A1(_08670_),
    .A2(_08668_),
    .B1(_08733_),
    .Y(_08734_));
 sky130_fd_sc_hd__nand2_1 _16649_ (.A(_08732_),
    .B(_08734_),
    .Y(_08735_));
 sky130_fd_sc_hd__or2_1 _16650_ (.A(_08732_),
    .B(_08734_),
    .X(_08736_));
 sky130_fd_sc_hd__nand2_1 _16651_ (.A(_08735_),
    .B(_08736_),
    .Y(_08737_));
 sky130_fd_sc_hd__xnor2_2 _16652_ (.A(_08690_),
    .B(_08737_),
    .Y(_08738_));
 sky130_fd_sc_hd__nor2_1 _16653_ (.A(\top0.pid_q.out[13] ),
    .B(_07704_),
    .Y(_08739_));
 sky130_fd_sc_hd__a21oi_2 _16654_ (.A1(_08619_),
    .A2(_08626_),
    .B1(_08618_),
    .Y(_08740_));
 sky130_fd_sc_hd__xor2_1 _16655_ (.A(\top0.pid_q.curr_int[13] ),
    .B(_08740_),
    .X(_08741_));
 sky130_fd_sc_hd__mux2_1 _16656_ (.A0(\top0.pid_q.out[13] ),
    .A1(_08739_),
    .S(_08741_),
    .X(_08742_));
 sky130_fd_sc_hd__a22o_1 _16657_ (.A1(\top0.pid_q.out[13] ),
    .A2(_07705_),
    .B1(_08742_),
    .B2(net544),
    .X(_08743_));
 sky130_fd_sc_hd__a31oi_1 _16658_ (.A1(net549),
    .A2(_07700_),
    .A3(_08738_),
    .B1(_08743_),
    .Y(_08744_));
 sky130_fd_sc_hd__nor2_1 _16659_ (.A(net16),
    .B(_08744_),
    .Y(_00146_));
 sky130_fd_sc_hd__a21bo_1 _16660_ (.A1(_08690_),
    .A2(_08735_),
    .B1_N(_08736_),
    .X(_08745_));
 sky130_fd_sc_hd__nand2_1 _16661_ (.A(_08312_),
    .B(_08693_),
    .Y(_08746_));
 sky130_fd_sc_hd__a21boi_2 _16662_ (.A1(_08692_),
    .A2(_08725_),
    .B1_N(_08726_),
    .Y(_08747_));
 sky130_fd_sc_hd__o21a_1 _16663_ (.A1(_08717_),
    .A2(_08722_),
    .B1(_08716_),
    .X(_08748_));
 sky130_fd_sc_hd__a21o_1 _16664_ (.A1(_08717_),
    .A2(_08722_),
    .B1(_08748_),
    .X(_08749_));
 sky130_fd_sc_hd__a21o_1 _16665_ (.A1(_08707_),
    .A2(_08714_),
    .B1(_08713_),
    .X(_08750_));
 sky130_fd_sc_hd__o21a_1 _16666_ (.A1(_07213_),
    .A2(_08711_),
    .B1(net459),
    .X(_08751_));
 sky130_fd_sc_hd__and2b_1 _16667_ (.A_N(_08654_),
    .B(_08711_),
    .X(_08752_));
 sky130_fd_sc_hd__o21a_1 _16668_ (.A1(_08751_),
    .A2(_08752_),
    .B1(net497),
    .X(_08753_));
 sky130_fd_sc_hd__xnor2_2 _16669_ (.A(_08527_),
    .B(_08753_),
    .Y(_08754_));
 sky130_fd_sc_hd__xnor2_1 _16670_ (.A(_08750_),
    .B(_08754_),
    .Y(_08755_));
 sky130_fd_sc_hd__o211a_1 _16671_ (.A1(_08453_),
    .A2(_08720_),
    .B1(net498),
    .C1(_08447_),
    .X(_08756_));
 sky130_fd_sc_hd__xnor2_1 _16672_ (.A(_08220_),
    .B(_08756_),
    .Y(_08757_));
 sky130_fd_sc_hd__nand2_1 _16673_ (.A(_07781_),
    .B(net444),
    .Y(_08758_));
 sky130_fd_sc_hd__nand2_1 _16674_ (.A(net447),
    .B(net500),
    .Y(_08759_));
 sky130_fd_sc_hd__nand2_1 _16675_ (.A(net504),
    .B(net445),
    .Y(_08760_));
 sky130_fd_sc_hd__xor2_1 _16676_ (.A(_08759_),
    .B(_08760_),
    .X(_08761_));
 sky130_fd_sc_hd__xnor2_2 _16677_ (.A(_08758_),
    .B(_08761_),
    .Y(_08762_));
 sky130_fd_sc_hd__o21a_1 _16678_ (.A1(_08701_),
    .A2(_08702_),
    .B1(_08703_),
    .X(_08763_));
 sky130_fd_sc_hd__a21oi_2 _16679_ (.A1(_08701_),
    .A2(_08702_),
    .B1(_08763_),
    .Y(_08764_));
 sky130_fd_sc_hd__nor2_1 _16680_ (.A(net449),
    .B(_08696_),
    .Y(_08765_));
 sky130_fd_sc_hd__and2_1 _16681_ (.A(net449),
    .B(_08696_),
    .X(_08766_));
 sky130_fd_sc_hd__or3b_1 _16682_ (.A(_08765_),
    .B(_08766_),
    .C_N(net498),
    .X(_08767_));
 sky130_fd_sc_hd__xnor2_1 _16683_ (.A(_08764_),
    .B(_08767_),
    .Y(_08768_));
 sky130_fd_sc_hd__xnor2_2 _16684_ (.A(_08762_),
    .B(_08768_),
    .Y(_08769_));
 sky130_fd_sc_hd__a21o_1 _16685_ (.A1(_08700_),
    .A2(_08705_),
    .B1(_08698_),
    .X(_08770_));
 sky130_fd_sc_hd__o21a_1 _16686_ (.A1(_08700_),
    .A2(_08705_),
    .B1(_08770_),
    .X(_08771_));
 sky130_fd_sc_hd__a22o_1 _16687_ (.A1(net452),
    .A2(net455),
    .B1(net500),
    .B2(net449),
    .X(_08772_));
 sky130_fd_sc_hd__o211a_1 _16688_ (.A1(net452),
    .A2(net455),
    .B1(net498),
    .C1(_08772_),
    .X(_08773_));
 sky130_fd_sc_hd__xnor2_2 _16689_ (.A(_08648_),
    .B(_08773_),
    .Y(_08774_));
 sky130_fd_sc_hd__xor2_1 _16690_ (.A(_08771_),
    .B(_08774_),
    .X(_08775_));
 sky130_fd_sc_hd__xnor2_1 _16691_ (.A(_08769_),
    .B(_08775_),
    .Y(_08776_));
 sky130_fd_sc_hd__or2_1 _16692_ (.A(_08757_),
    .B(_08776_),
    .X(_08777_));
 sky130_fd_sc_hd__and2_1 _16693_ (.A(_08757_),
    .B(_08776_),
    .X(_08778_));
 sky130_fd_sc_hd__inv_2 _16694_ (.A(_08778_),
    .Y(_08779_));
 sky130_fd_sc_hd__nand2_1 _16695_ (.A(_08777_),
    .B(_08779_),
    .Y(_08780_));
 sky130_fd_sc_hd__xnor2_1 _16696_ (.A(_08755_),
    .B(_08780_),
    .Y(_08781_));
 sky130_fd_sc_hd__xnor2_2 _16697_ (.A(_08749_),
    .B(_08781_),
    .Y(_08782_));
 sky130_fd_sc_hd__xor2_1 _16698_ (.A(_08747_),
    .B(_08782_),
    .X(_08783_));
 sky130_fd_sc_hd__xnor2_1 _16699_ (.A(_08746_),
    .B(_08783_),
    .Y(_08784_));
 sky130_fd_sc_hd__a21bo_1 _16700_ (.A1(_08730_),
    .A2(_08728_),
    .B1_N(_08664_),
    .X(_08785_));
 sky130_fd_sc_hd__o21a_1 _16701_ (.A1(_08730_),
    .A2(_08728_),
    .B1(_08785_),
    .X(_08786_));
 sky130_fd_sc_hd__and2_1 _16702_ (.A(_08784_),
    .B(_08786_),
    .X(_08787_));
 sky130_fd_sc_hd__or2_1 _16703_ (.A(_08784_),
    .B(_08786_),
    .X(_08788_));
 sky130_fd_sc_hd__inv_2 _16704_ (.A(_08788_),
    .Y(_08789_));
 sky130_fd_sc_hd__or2_1 _16705_ (.A(_08787_),
    .B(_08789_),
    .X(_08790_));
 sky130_fd_sc_hd__xnor2_2 _16706_ (.A(_08745_),
    .B(_08790_),
    .Y(_08791_));
 sky130_fd_sc_hd__nor2_1 _16707_ (.A(\top0.pid_q.out[14] ),
    .B(_07704_),
    .Y(_08792_));
 sky130_fd_sc_hd__a21o_1 _16708_ (.A1(\top0.pid_q.curr_int[13] ),
    .A2(_08740_),
    .B1(\top0.pid_q.out[13] ),
    .X(_08793_));
 sky130_fd_sc_hd__o21ai_1 _16709_ (.A1(\top0.pid_q.curr_int[13] ),
    .A2(_08740_),
    .B1(_08793_),
    .Y(_08794_));
 sky130_fd_sc_hd__xnor2_1 _16710_ (.A(\top0.pid_q.curr_int[14] ),
    .B(_08794_),
    .Y(_08795_));
 sky130_fd_sc_hd__mux2_1 _16711_ (.A0(\top0.pid_q.out[14] ),
    .A1(_08792_),
    .S(_08795_),
    .X(_08796_));
 sky130_fd_sc_hd__a22o_1 _16712_ (.A1(\top0.pid_q.out[14] ),
    .A2(_07705_),
    .B1(_08796_),
    .B2(net544),
    .X(_08797_));
 sky130_fd_sc_hd__a32o_1 _16713_ (.A1(_00011_),
    .A2(_07700_),
    .A3(_08791_),
    .B1(_08797_),
    .B2(_07800_),
    .X(_00147_));
 sky130_fd_sc_hd__o21a_1 _16714_ (.A1(_08747_),
    .A2(_08782_),
    .B1(_08746_),
    .X(_08798_));
 sky130_fd_sc_hd__a21oi_1 _16715_ (.A1(_08747_),
    .A2(_08782_),
    .B1(_08798_),
    .Y(_08799_));
 sky130_fd_sc_hd__and3_1 _16716_ (.A(_08757_),
    .B(_08754_),
    .C(_08776_),
    .X(_08800_));
 sky130_fd_sc_hd__nand2_1 _16717_ (.A(_08750_),
    .B(_08800_),
    .Y(_08801_));
 sky130_fd_sc_hd__a21o_1 _16718_ (.A1(_08754_),
    .A2(_08777_),
    .B1(_08778_),
    .X(_08802_));
 sky130_fd_sc_hd__o22a_1 _16719_ (.A1(_08754_),
    .A2(_08777_),
    .B1(_08802_),
    .B2(_08750_),
    .X(_08803_));
 sky130_fd_sc_hd__a21oi_1 _16720_ (.A1(_08750_),
    .A2(_08802_),
    .B1(_08800_),
    .Y(_08804_));
 sky130_fd_sc_hd__mux2_1 _16721_ (.A0(_08803_),
    .A1(_08804_),
    .S(_08749_),
    .X(_08805_));
 sky130_fd_sc_hd__o311a_1 _16722_ (.A1(_08750_),
    .A2(_08754_),
    .A3(_08777_),
    .B1(_08801_),
    .C1(_08805_),
    .X(_08806_));
 sky130_fd_sc_hd__a21bo_1 _16723_ (.A1(_08769_),
    .A2(_08774_),
    .B1_N(_08771_),
    .X(_08807_));
 sky130_fd_sc_hd__o21a_1 _16724_ (.A1(_08769_),
    .A2(_08774_),
    .B1(_08807_),
    .X(_08808_));
 sky130_fd_sc_hd__and3_1 _16725_ (.A(net449),
    .B(net452),
    .C(net455),
    .X(_08809_));
 sky130_fd_sc_hd__nor3_1 _16726_ (.A(net449),
    .B(net452),
    .C(net455),
    .Y(_08810_));
 sky130_fd_sc_hd__nor2_1 _16727_ (.A(_08809_),
    .B(_08810_),
    .Y(_08811_));
 sky130_fd_sc_hd__xnor2_1 _16728_ (.A(net447),
    .B(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__o21ai_1 _16729_ (.A1(net452),
    .A2(net455),
    .B1(_08772_),
    .Y(_08813_));
 sky130_fd_sc_hd__nand2_1 _16730_ (.A(_08718_),
    .B(_08813_),
    .Y(_08814_));
 sky130_fd_sc_hd__a2bb2o_1 _16731_ (.A1_N(_08654_),
    .A2_N(_08813_),
    .B1(_08814_),
    .B2(net459),
    .X(_08815_));
 sky130_fd_sc_hd__xnor2_1 _16732_ (.A(_08812_),
    .B(_08815_),
    .Y(_08816_));
 sky130_fd_sc_hd__nand2_1 _16733_ (.A(net498),
    .B(_08816_),
    .Y(_08817_));
 sky130_fd_sc_hd__a21bo_1 _16734_ (.A1(_08764_),
    .A2(_08762_),
    .B1_N(_08767_),
    .X(_08818_));
 sky130_fd_sc_hd__o21a_1 _16735_ (.A1(_08764_),
    .A2(_08762_),
    .B1(_08818_),
    .X(_08819_));
 sky130_fd_sc_hd__xnor2_1 _16736_ (.A(_08817_),
    .B(_08819_),
    .Y(_08820_));
 sky130_fd_sc_hd__o21ai_1 _16737_ (.A1(_08287_),
    .A2(_07781_),
    .B1(net444),
    .Y(_08821_));
 sky130_fd_sc_hd__and2_1 _16738_ (.A(net447),
    .B(_07781_),
    .X(_08822_));
 sky130_fd_sc_hd__and3b_1 _16739_ (.A_N(net445),
    .B(net444),
    .C(net504),
    .X(_08823_));
 sky130_fd_sc_hd__a21o_1 _16740_ (.A1(_08287_),
    .A2(net445),
    .B1(_08823_),
    .X(_08824_));
 sky130_fd_sc_hd__a32o_1 _16741_ (.A1(net445),
    .A2(_08703_),
    .A3(_08821_),
    .B1(_08822_),
    .B2(_08824_),
    .X(_08825_));
 sky130_fd_sc_hd__o21ai_1 _16742_ (.A1(net445),
    .A2(_08822_),
    .B1(net500),
    .Y(_08826_));
 sky130_fd_sc_hd__a32o_1 _16743_ (.A1(_07781_),
    .A2(net445),
    .A3(_08141_),
    .B1(_08826_),
    .B2(_08287_),
    .X(_08827_));
 sky130_fd_sc_hd__a22o_1 _16744_ (.A1(net500),
    .A2(_08825_),
    .B1(_08827_),
    .B2(net444),
    .X(_08828_));
 sky130_fd_sc_hd__xor2_1 _16745_ (.A(_08648_),
    .B(_08828_),
    .X(_08829_));
 sky130_fd_sc_hd__xnor2_1 _16746_ (.A(_08820_),
    .B(_08829_),
    .Y(_08830_));
 sky130_fd_sc_hd__xnor2_1 _16747_ (.A(_08808_),
    .B(_08830_),
    .Y(_08831_));
 sky130_fd_sc_hd__nor3_1 _16748_ (.A(_08142_),
    .B(_08721_),
    .C(_08753_),
    .Y(_08832_));
 sky130_fd_sc_hd__a21oi_1 _16749_ (.A1(_08721_),
    .A2(_08753_),
    .B1(_08832_),
    .Y(_08833_));
 sky130_fd_sc_hd__nor2_1 _16750_ (.A(_08526_),
    .B(_08753_),
    .Y(_08834_));
 sky130_fd_sc_hd__o22a_1 _16751_ (.A1(_08526_),
    .A2(_08833_),
    .B1(_08834_),
    .B2(_08312_),
    .X(_08835_));
 sky130_fd_sc_hd__nor2_1 _16752_ (.A(_08453_),
    .B(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__xnor2_1 _16753_ (.A(_08831_),
    .B(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__xnor2_1 _16754_ (.A(_08806_),
    .B(_08837_),
    .Y(_08838_));
 sky130_fd_sc_hd__xnor2_1 _16755_ (.A(_08799_),
    .B(_08838_),
    .Y(_08839_));
 sky130_fd_sc_hd__nor2_1 _16756_ (.A(_08787_),
    .B(_08839_),
    .Y(_08840_));
 sky130_fd_sc_hd__and2_1 _16757_ (.A(_08788_),
    .B(_08839_),
    .X(_08841_));
 sky130_fd_sc_hd__mux2_2 _16758_ (.A0(_08840_),
    .A1(_08841_),
    .S(_08745_),
    .X(_08842_));
 sky130_fd_sc_hd__nor2_1 _16759_ (.A(\top0.pid_q.out[15] ),
    .B(_07704_),
    .Y(_08843_));
 sky130_fd_sc_hd__nand2_1 _16760_ (.A(\top0.pid_q.out[14] ),
    .B(\top0.pid_q.curr_int[14] ),
    .Y(_08844_));
 sky130_fd_sc_hd__nor2_1 _16761_ (.A(\top0.pid_q.out[14] ),
    .B(\top0.pid_q.curr_int[14] ),
    .Y(_08845_));
 sky130_fd_sc_hd__a21o_1 _16762_ (.A1(_08794_),
    .A2(_08844_),
    .B1(_08845_),
    .X(_08846_));
 sky130_fd_sc_hd__xnor2_1 _16763_ (.A(\top0.pid_q.curr_int[15] ),
    .B(_08846_),
    .Y(_08847_));
 sky130_fd_sc_hd__mux2_1 _16764_ (.A0(\top0.pid_q.out[15] ),
    .A1(_08843_),
    .S(_08847_),
    .X(_08848_));
 sky130_fd_sc_hd__mux2_2 _16765_ (.A0(_08789_),
    .A1(_08787_),
    .S(_08839_),
    .X(_08849_));
 sky130_fd_sc_hd__and3_1 _16766_ (.A(\top0.pid_q.out[15] ),
    .B(_05442_),
    .C(_07704_),
    .X(_08850_));
 sky130_fd_sc_hd__a31o_1 _16767_ (.A1(_05448_),
    .A2(_07700_),
    .A3(_08849_),
    .B1(_08850_),
    .X(_08851_));
 sky130_fd_sc_hd__a31o_1 _16768_ (.A1(net544),
    .A2(net1019),
    .A3(_08848_),
    .B1(_08851_),
    .X(_08852_));
 sky130_fd_sc_hd__a31o_1 _16769_ (.A1(_00011_),
    .A2(_07700_),
    .A3(_08842_),
    .B1(_08852_),
    .X(_00148_));
 sky130_fd_sc_hd__or2_2 _16770_ (.A(\top0.pid_q.state[0] ),
    .B(net544),
    .X(_08853_));
 sky130_fd_sc_hd__nor2_4 _16771_ (.A(_07698_),
    .B(_08853_),
    .Y(_08854_));
 sky130_fd_sc_hd__nor2_4 _16772_ (.A(net15),
    .B(_08854_),
    .Y(_08855_));
 sky130_fd_sc_hd__buf_2 _16773_ (.A(_08855_),
    .X(_08856_));
 sky130_fd_sc_hd__and3_1 _16774_ (.A(net547),
    .B(_05442_),
    .C(_08854_),
    .X(_08857_));
 sky130_fd_sc_hd__clkbuf_2 _16775_ (.A(_08857_),
    .X(_08858_));
 sky130_fd_sc_hd__buf_2 _16776_ (.A(_08858_),
    .X(_08859_));
 sky130_fd_sc_hd__buf_2 _16777_ (.A(_05448_),
    .X(_08860_));
 sky130_fd_sc_hd__clkbuf_4 _16778_ (.A(_08854_),
    .X(_08861_));
 sky130_fd_sc_hd__and3_1 _16779_ (.A(\top0.kiq[0] ),
    .B(_08860_),
    .C(_08861_),
    .X(_08862_));
 sky130_fd_sc_hd__a221o_1 _16780_ (.A1(net542),
    .A2(_08856_),
    .B1(_08859_),
    .B2(net843),
    .C1(_08862_),
    .X(_00149_));
 sky130_fd_sc_hd__clkbuf_2 _16781_ (.A(_05448_),
    .X(_08863_));
 sky130_fd_sc_hd__and3_1 _16782_ (.A(\top0.kiq[1] ),
    .B(_08863_),
    .C(_08861_),
    .X(_08864_));
 sky130_fd_sc_hd__a221o_1 _16783_ (.A1(net539),
    .A2(_08856_),
    .B1(_08859_),
    .B2(net757),
    .C1(_08864_),
    .X(_00150_));
 sky130_fd_sc_hd__and3_1 _16784_ (.A(\top0.kiq[2] ),
    .B(_08863_),
    .C(_08861_),
    .X(_08865_));
 sky130_fd_sc_hd__a221o_1 _16785_ (.A1(\top0.pid_q.mult0.a[2] ),
    .A2(_08856_),
    .B1(_08859_),
    .B2(net787),
    .C1(_08865_),
    .X(_00151_));
 sky130_fd_sc_hd__clkbuf_2 _16786_ (.A(_08854_),
    .X(_08866_));
 sky130_fd_sc_hd__and3_1 _16787_ (.A(\top0.kiq[3] ),
    .B(_08863_),
    .C(_08866_),
    .X(_08867_));
 sky130_fd_sc_hd__a221o_1 _16788_ (.A1(net533),
    .A2(_08856_),
    .B1(_08859_),
    .B2(net789),
    .C1(_08867_),
    .X(_00152_));
 sky130_fd_sc_hd__and3_1 _16789_ (.A(\top0.kiq[4] ),
    .B(_08863_),
    .C(_08866_),
    .X(_08868_));
 sky130_fd_sc_hd__a221o_1 _16790_ (.A1(net1026),
    .A2(_08856_),
    .B1(_08859_),
    .B2(net751),
    .C1(_08868_),
    .X(_00153_));
 sky130_fd_sc_hd__and3_1 _16791_ (.A(\top0.kiq[5] ),
    .B(_08863_),
    .C(_08866_),
    .X(_08869_));
 sky130_fd_sc_hd__a221o_1 _16792_ (.A1(net527),
    .A2(_08856_),
    .B1(_08859_),
    .B2(net793),
    .C1(_08869_),
    .X(_00154_));
 sky130_fd_sc_hd__and3_1 _16793_ (.A(\top0.kiq[6] ),
    .B(_08863_),
    .C(_08866_),
    .X(_08870_));
 sky130_fd_sc_hd__a221o_1 _16794_ (.A1(net524),
    .A2(_08856_),
    .B1(_08859_),
    .B2(net719),
    .C1(_08870_),
    .X(_00155_));
 sky130_fd_sc_hd__and3_1 _16795_ (.A(\top0.kiq[7] ),
    .B(_08863_),
    .C(_08866_),
    .X(_08871_));
 sky130_fd_sc_hd__a221o_1 _16796_ (.A1(\top0.pid_q.mult0.a[7] ),
    .A2(_08856_),
    .B1(_08859_),
    .B2(net775),
    .C1(_08871_),
    .X(_00156_));
 sky130_fd_sc_hd__and3_1 _16797_ (.A(\top0.kiq[8] ),
    .B(_08863_),
    .C(_08866_),
    .X(_08872_));
 sky130_fd_sc_hd__a221o_1 _16798_ (.A1(net1028),
    .A2(_08856_),
    .B1(_08859_),
    .B2(net827),
    .C1(_08872_),
    .X(_00157_));
 sky130_fd_sc_hd__and3_1 _16799_ (.A(\top0.kiq[9] ),
    .B(_08863_),
    .C(_08866_),
    .X(_08873_));
 sky130_fd_sc_hd__a221o_1 _16800_ (.A1(net515),
    .A2(_08856_),
    .B1(_08859_),
    .B2(net734),
    .C1(_08873_),
    .X(_00158_));
 sky130_fd_sc_hd__and3_1 _16801_ (.A(\top0.kiq[10] ),
    .B(_08863_),
    .C(_08866_),
    .X(_08874_));
 sky130_fd_sc_hd__a221o_1 _16802_ (.A1(net512),
    .A2(_08855_),
    .B1(_08858_),
    .B2(net796),
    .C1(_08874_),
    .X(_00159_));
 sky130_fd_sc_hd__and3_1 _16803_ (.A(\top0.kiq[11] ),
    .B(_05448_),
    .C(_08866_),
    .X(_08875_));
 sky130_fd_sc_hd__a221o_1 _16804_ (.A1(net509),
    .A2(_08855_),
    .B1(_08858_),
    .B2(net713),
    .C1(_08875_),
    .X(_00160_));
 sky130_fd_sc_hd__and3_1 _16805_ (.A(\top0.kiq[12] ),
    .B(_05448_),
    .C(_08866_),
    .X(_08876_));
 sky130_fd_sc_hd__a221o_1 _16806_ (.A1(net506),
    .A2(_08855_),
    .B1(_08858_),
    .B2(net710),
    .C1(_08876_),
    .X(_00161_));
 sky130_fd_sc_hd__and3_1 _16807_ (.A(\top0.kiq[13] ),
    .B(_05448_),
    .C(_08854_),
    .X(_08877_));
 sky130_fd_sc_hd__a221o_1 _16808_ (.A1(net505),
    .A2(_08855_),
    .B1(_08858_),
    .B2(net703),
    .C1(_08877_),
    .X(_00162_));
 sky130_fd_sc_hd__and3_1 _16809_ (.A(\top0.kiq[14] ),
    .B(_05448_),
    .C(_08854_),
    .X(_08878_));
 sky130_fd_sc_hd__a221o_1 _16810_ (.A1(\top0.pid_q.mult0.a[14] ),
    .A2(_08855_),
    .B1(_08858_),
    .B2(net803),
    .C1(_08878_),
    .X(_00163_));
 sky130_fd_sc_hd__and3_1 _16811_ (.A(\top0.kiq[15] ),
    .B(_05448_),
    .C(_08854_),
    .X(_08879_));
 sky130_fd_sc_hd__a221o_1 _16812_ (.A1(\top0.pid_q.mult0.a[15] ),
    .A2(_08855_),
    .B1(_08858_),
    .B2(net937),
    .C1(_08879_),
    .X(_00164_));
 sky130_fd_sc_hd__or2_1 _16813_ (.A(_07698_),
    .B(_08853_),
    .X(_08880_));
 sky130_fd_sc_hd__buf_2 _16814_ (.A(_08880_),
    .X(_08881_));
 sky130_fd_sc_hd__clkbuf_4 _16815_ (.A(_08881_),
    .X(_08882_));
 sky130_fd_sc_hd__nand2_1 _16816_ (.A(\top0.matmul0.beta_pass[0] ),
    .B(_05438_),
    .Y(_08883_));
 sky130_fd_sc_hd__xnor2_1 _16817_ (.A(\top0.currT_r[0] ),
    .B(_08883_),
    .Y(_08884_));
 sky130_fd_sc_hd__and2_1 _16818_ (.A(net547),
    .B(_08884_),
    .X(_08885_));
 sky130_fd_sc_hd__xor2_1 _16819_ (.A(\top0.pid_q.prev_error[0] ),
    .B(\top0.pid_q.curr_error[0] ),
    .X(_08886_));
 sky130_fd_sc_hd__and2_1 _16820_ (.A(net550),
    .B(_08886_),
    .X(_08887_));
 sky130_fd_sc_hd__or2_1 _16821_ (.A(net496),
    .B(_08861_),
    .X(_08888_));
 sky130_fd_sc_hd__buf_4 _16822_ (.A(net1019),
    .X(_08889_));
 sky130_fd_sc_hd__o311a_1 _16823_ (.A1(_08882_),
    .A2(_08885_),
    .A3(_08887_),
    .B1(_08888_),
    .C1(_08889_),
    .X(_00165_));
 sky130_fd_sc_hd__buf_2 _16824_ (.A(_08861_),
    .X(_08890_));
 sky130_fd_sc_hd__and2b_1 _16825_ (.A_N(\top0.currT_r[0] ),
    .B(\top0.matmul0.beta_pass[0] ),
    .X(_08891_));
 sky130_fd_sc_hd__xor2_1 _16826_ (.A(\top0.matmul0.beta_pass[1] ),
    .B(_08891_),
    .X(_08892_));
 sky130_fd_sc_hd__nand2_1 _16827_ (.A(_05439_),
    .B(_08892_),
    .Y(_08893_));
 sky130_fd_sc_hd__xnor2_2 _16828_ (.A(\top0.currT_r[1] ),
    .B(_08893_),
    .Y(_08894_));
 sky130_fd_sc_hd__nand2_1 _16829_ (.A(\top0.pid_q.prev_error[0] ),
    .B(\top0.pid_q.curr_error[0] ),
    .Y(_08895_));
 sky130_fd_sc_hd__xor2_1 _16830_ (.A(\top0.pid_q.prev_error[1] ),
    .B(\top0.pid_q.curr_error[1] ),
    .X(_08896_));
 sky130_fd_sc_hd__xnor2_2 _16831_ (.A(_08895_),
    .B(_08896_),
    .Y(_08897_));
 sky130_fd_sc_hd__a221o_1 _16832_ (.A1(net547),
    .A2(_08894_),
    .B1(_08897_),
    .B2(net550),
    .C1(_08881_),
    .X(_08898_));
 sky130_fd_sc_hd__o211a_1 _16833_ (.A1(net492),
    .A2(_08890_),
    .B1(_08898_),
    .C1(_07710_),
    .X(_00166_));
 sky130_fd_sc_hd__buf_2 _16834_ (.A(_05601_),
    .X(_08899_));
 sky130_fd_sc_hd__buf_4 _16835_ (.A(_08899_),
    .X(_08900_));
 sky130_fd_sc_hd__or2b_1 _16836_ (.A(\top0.matmul0.beta_pass[1] ),
    .B_N(\top0.currT_r[1] ),
    .X(_08901_));
 sky130_fd_sc_hd__and2b_1 _16837_ (.A_N(\top0.currT_r[1] ),
    .B(\top0.matmul0.beta_pass[1] ),
    .X(_08902_));
 sky130_fd_sc_hd__a21oi_1 _16838_ (.A1(_08891_),
    .A2(_08901_),
    .B1(_08902_),
    .Y(_08903_));
 sky130_fd_sc_hd__xor2_1 _16839_ (.A(\top0.matmul0.beta_pass[2] ),
    .B(_08903_),
    .X(_08904_));
 sky130_fd_sc_hd__o21ai_1 _16840_ (.A1(_08900_),
    .A2(_08904_),
    .B1(\top0.currT_r[2] ),
    .Y(_08905_));
 sky130_fd_sc_hd__or3_1 _16841_ (.A(\top0.currT_r[2] ),
    .B(_08900_),
    .C(_08904_),
    .X(_08906_));
 sky130_fd_sc_hd__a21boi_2 _16842_ (.A1(_08905_),
    .A2(_08906_),
    .B1_N(net547),
    .Y(_08907_));
 sky130_fd_sc_hd__nand2_1 _16843_ (.A(\top0.pid_q.prev_error[1] ),
    .B(\top0.pid_q.curr_error[1] ),
    .Y(_08908_));
 sky130_fd_sc_hd__o211ai_2 _16844_ (.A1(\top0.pid_q.prev_error[1] ),
    .A2(\top0.pid_q.curr_error[1] ),
    .B1(\top0.pid_q.prev_error[0] ),
    .C1(\top0.pid_q.curr_error[0] ),
    .Y(_08909_));
 sky130_fd_sc_hd__xor2_1 _16845_ (.A(\top0.pid_q.prev_error[2] ),
    .B(\top0.pid_q.curr_error[2] ),
    .X(_08910_));
 sky130_fd_sc_hd__and3_1 _16846_ (.A(_08908_),
    .B(_08909_),
    .C(_08910_),
    .X(_08911_));
 sky130_fd_sc_hd__a21oi_1 _16847_ (.A1(_08908_),
    .A2(_08909_),
    .B1(_08910_),
    .Y(_08912_));
 sky130_fd_sc_hd__o21a_1 _16848_ (.A1(_08911_),
    .A2(_08912_),
    .B1(net550),
    .X(_08913_));
 sky130_fd_sc_hd__or2_1 _16849_ (.A(net488),
    .B(_08861_),
    .X(_08914_));
 sky130_fd_sc_hd__o311a_1 _16850_ (.A1(_08882_),
    .A2(_08907_),
    .A3(_08913_),
    .B1(_08914_),
    .C1(_08889_),
    .X(_00167_));
 sky130_fd_sc_hd__a21bo_1 _16851_ (.A1(\top0.currT_r[2] ),
    .A2(_08903_),
    .B1_N(\top0.matmul0.beta_pass[2] ),
    .X(_08915_));
 sky130_fd_sc_hd__or2_1 _16852_ (.A(\top0.currT_r[2] ),
    .B(_08903_),
    .X(_08916_));
 sky130_fd_sc_hd__a21o_1 _16853_ (.A1(_08915_),
    .A2(_08916_),
    .B1(_05601_),
    .X(_08917_));
 sky130_fd_sc_hd__nand2_1 _16854_ (.A(\top0.matmul0.beta_pass[3] ),
    .B(_05438_),
    .Y(_08918_));
 sky130_fd_sc_hd__xnor2_1 _16855_ (.A(\top0.currT_r[3] ),
    .B(_08918_),
    .Y(_08919_));
 sky130_fd_sc_hd__xnor2_2 _16856_ (.A(_08917_),
    .B(_08919_),
    .Y(_08920_));
 sky130_fd_sc_hd__inv_2 _16857_ (.A(\top0.pid_q.curr_error[2] ),
    .Y(_08921_));
 sky130_fd_sc_hd__a21o_1 _16858_ (.A1(_08908_),
    .A2(_08909_),
    .B1(_08921_),
    .X(_08922_));
 sky130_fd_sc_hd__inv_2 _16859_ (.A(\top0.pid_q.prev_error[2] ),
    .Y(_08923_));
 sky130_fd_sc_hd__a31o_1 _16860_ (.A1(_08921_),
    .A2(_08908_),
    .A3(_08909_),
    .B1(_08923_),
    .X(_08924_));
 sky130_fd_sc_hd__and2_1 _16861_ (.A(_08922_),
    .B(_08924_),
    .X(_08925_));
 sky130_fd_sc_hd__xnor2_1 _16862_ (.A(\top0.pid_q.prev_error[3] ),
    .B(\top0.pid_q.curr_error[3] ),
    .Y(_08926_));
 sky130_fd_sc_hd__xnor2_1 _16863_ (.A(_08925_),
    .B(_08926_),
    .Y(_08927_));
 sky130_fd_sc_hd__inv_2 _16864_ (.A(_08927_),
    .Y(_08928_));
 sky130_fd_sc_hd__a221o_1 _16865_ (.A1(net546),
    .A2(_08920_),
    .B1(_08928_),
    .B2(net550),
    .C1(_08881_),
    .X(_08929_));
 sky130_fd_sc_hd__buf_2 _16866_ (.A(net1019),
    .X(_08930_));
 sky130_fd_sc_hd__o211a_1 _16867_ (.A1(net483),
    .A2(_08890_),
    .B1(_08929_),
    .C1(_08930_),
    .X(_00168_));
 sky130_fd_sc_hd__a21bo_1 _16868_ (.A1(\top0.currT_r[3] ),
    .A2(_08917_),
    .B1_N(\top0.matmul0.beta_pass[3] ),
    .X(_08931_));
 sky130_fd_sc_hd__o21a_1 _16869_ (.A1(\top0.currT_r[3] ),
    .A2(_08917_),
    .B1(_08931_),
    .X(_08932_));
 sky130_fd_sc_hd__xnor2_1 _16870_ (.A(\top0.matmul0.beta_pass[4] ),
    .B(_08932_),
    .Y(_08933_));
 sky130_fd_sc_hd__nand2_1 _16871_ (.A(_05438_),
    .B(_08933_),
    .Y(_08934_));
 sky130_fd_sc_hd__xnor2_2 _16872_ (.A(\top0.currT_r[4] ),
    .B(_08934_),
    .Y(_08935_));
 sky130_fd_sc_hd__inv_2 _16873_ (.A(\top0.pid_q.curr_error[3] ),
    .Y(_08936_));
 sky130_fd_sc_hd__inv_2 _16874_ (.A(\top0.pid_q.prev_error[3] ),
    .Y(_08937_));
 sky130_fd_sc_hd__a31o_1 _16875_ (.A1(_08936_),
    .A2(_08922_),
    .A3(_08924_),
    .B1(_08937_),
    .X(_08938_));
 sky130_fd_sc_hd__o21ai_2 _16876_ (.A1(_08936_),
    .A2(_08925_),
    .B1(_08938_),
    .Y(_08939_));
 sky130_fd_sc_hd__xor2_1 _16877_ (.A(\top0.pid_q.prev_error[4] ),
    .B(\top0.pid_q.curr_error[4] ),
    .X(_08940_));
 sky130_fd_sc_hd__xnor2_1 _16878_ (.A(_08939_),
    .B(_08940_),
    .Y(_08941_));
 sky130_fd_sc_hd__inv_2 _16879_ (.A(_08941_),
    .Y(_08942_));
 sky130_fd_sc_hd__a221o_1 _16880_ (.A1(net546),
    .A2(_08935_),
    .B1(_08942_),
    .B2(net550),
    .C1(_08881_),
    .X(_08943_));
 sky130_fd_sc_hd__o211a_1 _16881_ (.A1(net476),
    .A2(_08890_),
    .B1(_08943_),
    .C1(_08930_),
    .X(_00169_));
 sky130_fd_sc_hd__inv_2 _16882_ (.A(\top0.matmul0.beta_pass[4] ),
    .Y(_08944_));
 sky130_fd_sc_hd__o221a_1 _16883_ (.A1(_08944_),
    .A2(\top0.currT_r[4] ),
    .B1(_08917_),
    .B2(\top0.currT_r[3] ),
    .C1(_08931_),
    .X(_08945_));
 sky130_fd_sc_hd__a21o_1 _16884_ (.A1(_08944_),
    .A2(\top0.currT_r[4] ),
    .B1(_08945_),
    .X(_08946_));
 sky130_fd_sc_hd__xnor2_1 _16885_ (.A(\top0.matmul0.beta_pass[5] ),
    .B(_08946_),
    .Y(_08947_));
 sky130_fd_sc_hd__nand2_1 _16886_ (.A(_05439_),
    .B(_08947_),
    .Y(_08948_));
 sky130_fd_sc_hd__xnor2_2 _16887_ (.A(\top0.currT_r[5] ),
    .B(_08948_),
    .Y(_08949_));
 sky130_fd_sc_hd__a21o_1 _16888_ (.A1(\top0.pid_q.curr_error[4] ),
    .A2(_08939_),
    .B1(\top0.pid_q.prev_error[4] ),
    .X(_08950_));
 sky130_fd_sc_hd__o21a_1 _16889_ (.A1(\top0.pid_q.curr_error[4] ),
    .A2(_08939_),
    .B1(_08950_),
    .X(_08951_));
 sky130_fd_sc_hd__xor2_1 _16890_ (.A(\top0.pid_q.prev_error[5] ),
    .B(\top0.pid_q.curr_error[5] ),
    .X(_08952_));
 sky130_fd_sc_hd__or2_1 _16891_ (.A(_08951_),
    .B(_08952_),
    .X(_08953_));
 sky130_fd_sc_hd__nand2_1 _16892_ (.A(_08951_),
    .B(_08952_),
    .Y(_08954_));
 sky130_fd_sc_hd__and3_1 _16893_ (.A(net550),
    .B(_08953_),
    .C(_08954_),
    .X(_08955_));
 sky130_fd_sc_hd__a211o_1 _16894_ (.A1(net546),
    .A2(_08949_),
    .B1(_08955_),
    .C1(_08882_),
    .X(_08956_));
 sky130_fd_sc_hd__o211a_1 _16895_ (.A1(net473),
    .A2(_08890_),
    .B1(_08956_),
    .C1(_08930_),
    .X(_00170_));
 sky130_fd_sc_hd__a21bo_1 _16896_ (.A1(\top0.currT_r[5] ),
    .A2(_08946_),
    .B1_N(\top0.matmul0.beta_pass[5] ),
    .X(_08957_));
 sky130_fd_sc_hd__or2_1 _16897_ (.A(\top0.currT_r[5] ),
    .B(_08946_),
    .X(_08958_));
 sky130_fd_sc_hd__a21o_1 _16898_ (.A1(_08957_),
    .A2(_08958_),
    .B1(_05601_),
    .X(_08959_));
 sky130_fd_sc_hd__and3_1 _16899_ (.A(\top0.matmul0.done_pass ),
    .B(\top0.matmul0.state[1] ),
    .C(\top0.matmul0.beta_pass[6] ),
    .X(_08960_));
 sky130_fd_sc_hd__xor2_1 _16900_ (.A(\top0.currT_r[6] ),
    .B(_08960_),
    .X(_08961_));
 sky130_fd_sc_hd__xnor2_2 _16901_ (.A(_08959_),
    .B(_08961_),
    .Y(_08962_));
 sky130_fd_sc_hd__or2_1 _16902_ (.A(\top0.pid_q.curr_error[5] ),
    .B(_08951_),
    .X(_08963_));
 sky130_fd_sc_hd__a21o_1 _16903_ (.A1(\top0.pid_q.curr_error[5] ),
    .A2(_08951_),
    .B1(\top0.pid_q.prev_error[5] ),
    .X(_08964_));
 sky130_fd_sc_hd__and2_1 _16904_ (.A(_08963_),
    .B(_08964_),
    .X(_08965_));
 sky130_fd_sc_hd__xor2_1 _16905_ (.A(\top0.pid_q.prev_error[6] ),
    .B(\top0.pid_q.curr_error[6] ),
    .X(_08966_));
 sky130_fd_sc_hd__xnor2_1 _16906_ (.A(_08965_),
    .B(_08966_),
    .Y(_08967_));
 sky130_fd_sc_hd__and2b_1 _16907_ (.A_N(_08967_),
    .B(net550),
    .X(_08968_));
 sky130_fd_sc_hd__a211o_1 _16908_ (.A1(net546),
    .A2(_08962_),
    .B1(_08968_),
    .C1(_08882_),
    .X(_08969_));
 sky130_fd_sc_hd__o211a_1 _16909_ (.A1(net468),
    .A2(_08890_),
    .B1(_08969_),
    .C1(_08930_),
    .X(_00171_));
 sky130_fd_sc_hd__o21ba_1 _16910_ (.A1(\top0.currT_r[6] ),
    .A2(_08959_),
    .B1_N(_08960_),
    .X(_08970_));
 sky130_fd_sc_hd__a21o_1 _16911_ (.A1(\top0.currT_r[6] ),
    .A2(_08959_),
    .B1(_08970_),
    .X(_08971_));
 sky130_fd_sc_hd__nand2_1 _16912_ (.A(\top0.matmul0.beta_pass[7] ),
    .B(_05436_),
    .Y(_08972_));
 sky130_fd_sc_hd__xnor2_1 _16913_ (.A(\top0.currT_r[7] ),
    .B(_08972_),
    .Y(_08973_));
 sky130_fd_sc_hd__xnor2_2 _16914_ (.A(_08971_),
    .B(_08973_),
    .Y(_08974_));
 sky130_fd_sc_hd__a21o_1 _16915_ (.A1(_08963_),
    .A2(_08964_),
    .B1(\top0.pid_q.curr_error[6] ),
    .X(_08975_));
 sky130_fd_sc_hd__and3_1 _16916_ (.A(\top0.pid_q.curr_error[6] ),
    .B(_08963_),
    .C(_08964_),
    .X(_08976_));
 sky130_fd_sc_hd__a21oi_2 _16917_ (.A1(\top0.pid_q.prev_error[6] ),
    .A2(_08975_),
    .B1(_08976_),
    .Y(_08977_));
 sky130_fd_sc_hd__xnor2_1 _16918_ (.A(\top0.pid_q.prev_error[7] ),
    .B(\top0.pid_q.curr_error[7] ),
    .Y(_08978_));
 sky130_fd_sc_hd__nand2_1 _16919_ (.A(_08977_),
    .B(_08978_),
    .Y(_08979_));
 sky130_fd_sc_hd__or2_1 _16920_ (.A(_08977_),
    .B(_08978_),
    .X(_08980_));
 sky130_fd_sc_hd__and3_1 _16921_ (.A(net550),
    .B(_08979_),
    .C(_08980_),
    .X(_08981_));
 sky130_fd_sc_hd__a211o_1 _16922_ (.A1(net546),
    .A2(_08974_),
    .B1(_08981_),
    .C1(_08882_),
    .X(_08982_));
 sky130_fd_sc_hd__o211a_1 _16923_ (.A1(net466),
    .A2(_08890_),
    .B1(_08982_),
    .C1(_08930_),
    .X(_00172_));
 sky130_fd_sc_hd__o21a_1 _16924_ (.A1(\top0.currT_r[7] ),
    .A2(_08971_),
    .B1(_08972_),
    .X(_08983_));
 sky130_fd_sc_hd__a21o_1 _16925_ (.A1(\top0.currT_r[7] ),
    .A2(_08971_),
    .B1(_08983_),
    .X(_08984_));
 sky130_fd_sc_hd__nand2_1 _16926_ (.A(\top0.matmul0.beta_pass[8] ),
    .B(_05436_),
    .Y(_08985_));
 sky130_fd_sc_hd__xnor2_1 _16927_ (.A(\top0.currT_r[8] ),
    .B(_08985_),
    .Y(_08986_));
 sky130_fd_sc_hd__xnor2_2 _16928_ (.A(_08984_),
    .B(_08986_),
    .Y(_08987_));
 sky130_fd_sc_hd__inv_2 _16929_ (.A(\top0.pid_q.curr_error[7] ),
    .Y(_08988_));
 sky130_fd_sc_hd__o21ba_1 _16930_ (.A1(_08988_),
    .A2(_08977_),
    .B1_N(\top0.pid_q.prev_error[7] ),
    .X(_08989_));
 sky130_fd_sc_hd__a21o_1 _16931_ (.A1(_08988_),
    .A2(_08977_),
    .B1(_08989_),
    .X(_08990_));
 sky130_fd_sc_hd__xnor2_1 _16932_ (.A(\top0.pid_q.prev_error[8] ),
    .B(\top0.pid_q.curr_error[8] ),
    .Y(_08991_));
 sky130_fd_sc_hd__nand2_1 _16933_ (.A(_08990_),
    .B(_08991_),
    .Y(_08992_));
 sky130_fd_sc_hd__or2_1 _16934_ (.A(_08990_),
    .B(_08991_),
    .X(_08993_));
 sky130_fd_sc_hd__and3_1 _16935_ (.A(net550),
    .B(_08992_),
    .C(_08993_),
    .X(_08994_));
 sky130_fd_sc_hd__a211o_1 _16936_ (.A1(\top0.pid_q.state[3] ),
    .A2(_08987_),
    .B1(_08994_),
    .C1(_08882_),
    .X(_08995_));
 sky130_fd_sc_hd__o211a_1 _16937_ (.A1(net461),
    .A2(_08890_),
    .B1(_08995_),
    .C1(_08930_),
    .X(_00173_));
 sky130_fd_sc_hd__o21a_1 _16938_ (.A1(\top0.currT_r[8] ),
    .A2(_08984_),
    .B1(_08985_),
    .X(_08996_));
 sky130_fd_sc_hd__a21o_1 _16939_ (.A1(\top0.currT_r[8] ),
    .A2(_08984_),
    .B1(_08996_),
    .X(_08997_));
 sky130_fd_sc_hd__a21bo_1 _16940_ (.A1(\top0.matmul0.beta_pass[9] ),
    .A2(_05437_),
    .B1_N(\top0.currT_r[9] ),
    .X(_08998_));
 sky130_fd_sc_hd__or3b_1 _16941_ (.A(\top0.currT_r[9] ),
    .B(_08899_),
    .C_N(\top0.matmul0.beta_pass[9] ),
    .X(_08999_));
 sky130_fd_sc_hd__and3_1 _16942_ (.A(_08997_),
    .B(_08998_),
    .C(_08999_),
    .X(_09000_));
 sky130_fd_sc_hd__a21o_1 _16943_ (.A1(_08998_),
    .A2(_08999_),
    .B1(_08997_),
    .X(_09001_));
 sky130_fd_sc_hd__and3b_1 _16944_ (.A_N(_09000_),
    .B(_09001_),
    .C(net547),
    .X(_09002_));
 sky130_fd_sc_hd__inv_2 _16945_ (.A(\top0.pid_q.curr_error[8] ),
    .Y(_09003_));
 sky130_fd_sc_hd__o21ba_1 _16946_ (.A1(_09003_),
    .A2(_08990_),
    .B1_N(\top0.pid_q.prev_error[8] ),
    .X(_09004_));
 sky130_fd_sc_hd__a21o_1 _16947_ (.A1(_09003_),
    .A2(_08990_),
    .B1(_09004_),
    .X(_09005_));
 sky130_fd_sc_hd__xnor2_1 _16948_ (.A(\top0.pid_q.prev_error[9] ),
    .B(\top0.pid_q.curr_error[9] ),
    .Y(_09006_));
 sky130_fd_sc_hd__nand2_1 _16949_ (.A(_09005_),
    .B(_09006_),
    .Y(_09007_));
 sky130_fd_sc_hd__or2_1 _16950_ (.A(_09005_),
    .B(_09006_),
    .X(_09008_));
 sky130_fd_sc_hd__and3_1 _16951_ (.A(net550),
    .B(_09007_),
    .C(_09008_),
    .X(_09009_));
 sky130_fd_sc_hd__or2_1 _16952_ (.A(net459),
    .B(_08861_),
    .X(_09010_));
 sky130_fd_sc_hd__o311a_1 _16953_ (.A1(_08882_),
    .A2(_09002_),
    .A3(_09009_),
    .B1(_09010_),
    .C1(_08889_),
    .X(_00174_));
 sky130_fd_sc_hd__a21bo_1 _16954_ (.A1(\top0.currT_r[9] ),
    .A2(_08997_),
    .B1_N(\top0.matmul0.beta_pass[9] ),
    .X(_09011_));
 sky130_fd_sc_hd__o21ai_1 _16955_ (.A1(\top0.currT_r[9] ),
    .A2(_08997_),
    .B1(_09011_),
    .Y(_09012_));
 sky130_fd_sc_hd__xnor2_1 _16956_ (.A(net429),
    .B(_09012_),
    .Y(_09013_));
 sky130_fd_sc_hd__o21ai_1 _16957_ (.A1(_08900_),
    .A2(_09013_),
    .B1(\top0.currT_r[10] ),
    .Y(_09014_));
 sky130_fd_sc_hd__or3_1 _16958_ (.A(\top0.currT_r[10] ),
    .B(_08900_),
    .C(_09013_),
    .X(_09015_));
 sky130_fd_sc_hd__a21boi_2 _16959_ (.A1(_09014_),
    .A2(_09015_),
    .B1_N(net547),
    .Y(_09016_));
 sky130_fd_sc_hd__inv_2 _16960_ (.A(\top0.pid_q.curr_error[9] ),
    .Y(_09017_));
 sky130_fd_sc_hd__o21ba_1 _16961_ (.A1(_09017_),
    .A2(_09005_),
    .B1_N(\top0.pid_q.prev_error[9] ),
    .X(_09018_));
 sky130_fd_sc_hd__a21o_1 _16962_ (.A1(_09017_),
    .A2(_09005_),
    .B1(_09018_),
    .X(_09019_));
 sky130_fd_sc_hd__xnor2_1 _16963_ (.A(\top0.pid_q.prev_error[10] ),
    .B(\top0.pid_q.curr_error[10] ),
    .Y(_09020_));
 sky130_fd_sc_hd__nand2_1 _16964_ (.A(_09019_),
    .B(_09020_),
    .Y(_09021_));
 sky130_fd_sc_hd__or2_1 _16965_ (.A(_09019_),
    .B(_09020_),
    .X(_09022_));
 sky130_fd_sc_hd__and3_1 _16966_ (.A(net552),
    .B(_09021_),
    .C(_09022_),
    .X(_09023_));
 sky130_fd_sc_hd__or2_1 _16967_ (.A(net455),
    .B(_08861_),
    .X(_09024_));
 sky130_fd_sc_hd__o311a_1 _16968_ (.A1(_08882_),
    .A2(_09016_),
    .A3(_09023_),
    .B1(_09024_),
    .C1(_07800_),
    .X(_00175_));
 sky130_fd_sc_hd__inv_2 _16969_ (.A(\top0.pid_q.curr_error[10] ),
    .Y(_09025_));
 sky130_fd_sc_hd__o21ba_1 _16970_ (.A1(_09025_),
    .A2(_09019_),
    .B1_N(\top0.pid_q.prev_error[10] ),
    .X(_09026_));
 sky130_fd_sc_hd__a21o_1 _16971_ (.A1(_09025_),
    .A2(_09019_),
    .B1(_09026_),
    .X(_09027_));
 sky130_fd_sc_hd__xor2_1 _16972_ (.A(\top0.pid_q.prev_error[11] ),
    .B(\top0.pid_q.curr_error[11] ),
    .X(_09028_));
 sky130_fd_sc_hd__xnor2_1 _16973_ (.A(_09027_),
    .B(_09028_),
    .Y(_09029_));
 sky130_fd_sc_hd__o21ai_1 _16974_ (.A1(\top0.currT_r[9] ),
    .A2(_08997_),
    .B1(\top0.currT_r[10] ),
    .Y(_09030_));
 sky130_fd_sc_hd__and2b_1 _16975_ (.A_N(net429),
    .B(\top0.currT_r[10] ),
    .X(_09031_));
 sky130_fd_sc_hd__o2bb2a_1 _16976_ (.A1_N(net429),
    .A2_N(_09030_),
    .B1(_09031_),
    .B2(_09011_),
    .X(_09032_));
 sky130_fd_sc_hd__o32a_2 _16977_ (.A1(\top0.currT_r[9] ),
    .A2(\top0.currT_r[10] ),
    .A3(_08997_),
    .B1(_09032_),
    .B2(_05601_),
    .X(_09033_));
 sky130_fd_sc_hd__nand2_1 _16978_ (.A(\top0.matmul0.beta_pass[11] ),
    .B(_05438_),
    .Y(_09034_));
 sky130_fd_sc_hd__xnor2_1 _16979_ (.A(\top0.currT_r[11] ),
    .B(_09034_),
    .Y(_09035_));
 sky130_fd_sc_hd__xnor2_2 _16980_ (.A(_09033_),
    .B(_09035_),
    .Y(_09036_));
 sky130_fd_sc_hd__a221o_1 _16981_ (.A1(net552),
    .A2(_09029_),
    .B1(_09036_),
    .B2(\top0.pid_q.state[3] ),
    .C1(_08881_),
    .X(_09037_));
 sky130_fd_sc_hd__o211a_1 _16982_ (.A1(net452),
    .A2(_08890_),
    .B1(_09037_),
    .C1(_08930_),
    .X(_00176_));
 sky130_fd_sc_hd__nand2_1 _16983_ (.A(\top0.currT_r[11] ),
    .B(_09033_),
    .Y(_09038_));
 sky130_fd_sc_hd__or2_1 _16984_ (.A(\top0.currT_r[11] ),
    .B(_09033_),
    .X(_09039_));
 sky130_fd_sc_hd__a21bo_1 _16985_ (.A1(\top0.matmul0.beta_pass[11] ),
    .A2(_09038_),
    .B1_N(_09039_),
    .X(_09040_));
 sky130_fd_sc_hd__xor2_1 _16986_ (.A(\top0.matmul0.beta_pass[12] ),
    .B(_09040_),
    .X(_09041_));
 sky130_fd_sc_hd__inv_2 _16987_ (.A(\top0.currT_r[12] ),
    .Y(_09042_));
 sky130_fd_sc_hd__a21oi_1 _16988_ (.A1(_05438_),
    .A2(_09041_),
    .B1(_09042_),
    .Y(_09043_));
 sky130_fd_sc_hd__and3_1 _16989_ (.A(_09042_),
    .B(_05438_),
    .C(_09041_),
    .X(_09044_));
 sky130_fd_sc_hd__o21a_1 _16990_ (.A1(_09043_),
    .A2(_09044_),
    .B1(net547),
    .X(_09045_));
 sky130_fd_sc_hd__xor2_1 _16991_ (.A(\top0.pid_q.prev_error[12] ),
    .B(\top0.pid_q.curr_error[12] ),
    .X(_09046_));
 sky130_fd_sc_hd__nor2_1 _16992_ (.A(\top0.pid_q.prev_error[11] ),
    .B(\top0.pid_q.curr_error[11] ),
    .Y(_09047_));
 sky130_fd_sc_hd__nand2_1 _16993_ (.A(\top0.pid_q.prev_error[11] ),
    .B(\top0.pid_q.curr_error[11] ),
    .Y(_09048_));
 sky130_fd_sc_hd__o21a_1 _16994_ (.A1(_09027_),
    .A2(_09047_),
    .B1(_09048_),
    .X(_09049_));
 sky130_fd_sc_hd__xnor2_1 _16995_ (.A(_09046_),
    .B(_09049_),
    .Y(_09050_));
 sky130_fd_sc_hd__a21o_1 _16996_ (.A1(net551),
    .A2(_09050_),
    .B1(_08881_),
    .X(_09051_));
 sky130_fd_sc_hd__o221a_1 _16997_ (.A1(net449),
    .A2(_08861_),
    .B1(_09045_),
    .B2(_09051_),
    .C1(_08889_),
    .X(_00177_));
 sky130_fd_sc_hd__o21ba_1 _16998_ (.A1(\top0.pid_q.prev_error[12] ),
    .A2(\top0.pid_q.curr_error[12] ),
    .B1_N(_09049_),
    .X(_09052_));
 sky130_fd_sc_hd__a21o_1 _16999_ (.A1(\top0.pid_q.prev_error[12] ),
    .A2(\top0.pid_q.curr_error[12] ),
    .B1(_09052_),
    .X(_09053_));
 sky130_fd_sc_hd__xnor2_1 _17000_ (.A(\top0.pid_q.prev_error[13] ),
    .B(\top0.pid_q.curr_error[13] ),
    .Y(_09054_));
 sky130_fd_sc_hd__xnor2_1 _17001_ (.A(_09053_),
    .B(_09054_),
    .Y(_09055_));
 sky130_fd_sc_hd__a21bo_1 _17002_ (.A1(\top0.currT_r[12] ),
    .A2(_09039_),
    .B1_N(\top0.matmul0.beta_pass[12] ),
    .X(_09056_));
 sky130_fd_sc_hd__o211a_1 _17003_ (.A1(\top0.matmul0.beta_pass[12] ),
    .A2(_09042_),
    .B1(_05436_),
    .C1(\top0.matmul0.beta_pass[11] ),
    .X(_09057_));
 sky130_fd_sc_hd__o2bb2a_1 _17004_ (.A1_N(_09057_),
    .A2_N(_09038_),
    .B1(\top0.currT_r[12] ),
    .B2(_09039_),
    .X(_09058_));
 sky130_fd_sc_hd__o21a_1 _17005_ (.A1(_08899_),
    .A2(_09056_),
    .B1(_09058_),
    .X(_09059_));
 sky130_fd_sc_hd__nand2_1 _17006_ (.A(\top0.matmul0.beta_pass[13] ),
    .B(_05437_),
    .Y(_09060_));
 sky130_fd_sc_hd__xnor2_1 _17007_ (.A(\top0.currT_r[13] ),
    .B(_09060_),
    .Y(_09061_));
 sky130_fd_sc_hd__xnor2_1 _17008_ (.A(_09059_),
    .B(_09061_),
    .Y(_09062_));
 sky130_fd_sc_hd__and2_1 _17009_ (.A(net547),
    .B(_09062_),
    .X(_09063_));
 sky130_fd_sc_hd__a211o_1 _17010_ (.A1(net551),
    .A2(_09055_),
    .B1(_09063_),
    .C1(_08882_),
    .X(_09064_));
 sky130_fd_sc_hd__o211a_1 _17011_ (.A1(net448),
    .A2(_08890_),
    .B1(_09064_),
    .C1(_08930_),
    .X(_00178_));
 sky130_fd_sc_hd__and4_1 _17012_ (.A(_05662_),
    .B(net428),
    .C(\top0.currT_r[13] ),
    .D(_05437_),
    .X(_09065_));
 sky130_fd_sc_hd__o2111a_1 _17013_ (.A1(_05662_),
    .A2(\top0.currT_r[13] ),
    .B1(_05437_),
    .C1(_09059_),
    .D1(net428),
    .X(_09066_));
 sky130_fd_sc_hd__a2111o_1 _17014_ (.A1(_05662_),
    .A2(\top0.currT_r[13] ),
    .B1(_08899_),
    .C1(_09059_),
    .D1(net428),
    .X(_09067_));
 sky130_fd_sc_hd__or4_1 _17015_ (.A(_05662_),
    .B(net428),
    .C(\top0.currT_r[13] ),
    .D(_08899_),
    .X(_09068_));
 sky130_fd_sc_hd__and4bb_1 _17016_ (.A_N(_09065_),
    .B_N(_09066_),
    .C(_09067_),
    .D(_09068_),
    .X(_09069_));
 sky130_fd_sc_hd__xnor2_2 _17017_ (.A(\top0.currT_r[14] ),
    .B(_09069_),
    .Y(_09070_));
 sky130_fd_sc_hd__or2_1 _17018_ (.A(\top0.pid_q.prev_error[13] ),
    .B(\top0.pid_q.curr_error[13] ),
    .X(_09071_));
 sky130_fd_sc_hd__and2_1 _17019_ (.A(\top0.pid_q.prev_error[13] ),
    .B(\top0.pid_q.curr_error[13] ),
    .X(_09072_));
 sky130_fd_sc_hd__a21o_1 _17020_ (.A1(_09053_),
    .A2(_09071_),
    .B1(_09072_),
    .X(_09073_));
 sky130_fd_sc_hd__and2_1 _17021_ (.A(\top0.pid_q.prev_error[14] ),
    .B(\top0.pid_q.curr_error[14] ),
    .X(_09074_));
 sky130_fd_sc_hd__or2_1 _17022_ (.A(\top0.pid_q.prev_error[14] ),
    .B(\top0.pid_q.curr_error[14] ),
    .X(_09075_));
 sky130_fd_sc_hd__or2b_1 _17023_ (.A(_09074_),
    .B_N(_09075_),
    .X(_09076_));
 sky130_fd_sc_hd__xnor2_1 _17024_ (.A(_09073_),
    .B(_09076_),
    .Y(_09077_));
 sky130_fd_sc_hd__a221o_1 _17025_ (.A1(\top0.pid_q.state[3] ),
    .A2(_09070_),
    .B1(_09077_),
    .B2(net551),
    .C1(_08881_),
    .X(_09078_));
 sky130_fd_sc_hd__o211a_1 _17026_ (.A1(net445),
    .A2(_08890_),
    .B1(_09078_),
    .C1(_08930_),
    .X(_00179_));
 sky130_fd_sc_hd__or2_1 _17027_ (.A(\top0.currT_r[13] ),
    .B(\top0.currT_r[14] ),
    .X(_09079_));
 sky130_fd_sc_hd__or3_1 _17028_ (.A(_05662_),
    .B(\top0.currT_r[14] ),
    .C(_08899_),
    .X(_09080_));
 sky130_fd_sc_hd__inv_2 _17029_ (.A(net428),
    .Y(_09081_));
 sky130_fd_sc_hd__or3_1 _17030_ (.A(_09081_),
    .B(\top0.currT_r[13] ),
    .C(_08899_),
    .X(_09082_));
 sky130_fd_sc_hd__or3_1 _17031_ (.A(_05662_),
    .B(_09081_),
    .C(_08899_),
    .X(_09083_));
 sky130_fd_sc_hd__a41o_1 _17032_ (.A1(_09079_),
    .A2(_09080_),
    .A3(_09082_),
    .A4(_09083_),
    .B1(_09059_),
    .X(_09084_));
 sky130_fd_sc_hd__a2111o_1 _17033_ (.A1(_09081_),
    .A2(\top0.currT_r[14] ),
    .B1(_08900_),
    .C1(\top0.currT_r[13] ),
    .D1(_05662_),
    .X(_09085_));
 sky130_fd_sc_hd__o31a_1 _17034_ (.A1(_09081_),
    .A2(\top0.currT_r[14] ),
    .A3(_08900_),
    .B1(_09085_),
    .X(_09086_));
 sky130_fd_sc_hd__nand2_1 _17035_ (.A(_09084_),
    .B(_09086_),
    .Y(_09087_));
 sky130_fd_sc_hd__nand2_1 _17036_ (.A(\top0.matmul0.beta_pass[15] ),
    .B(_05438_),
    .Y(_09088_));
 sky130_fd_sc_hd__xor2_1 _17037_ (.A(\top0.currT_r[15] ),
    .B(_09088_),
    .X(_09089_));
 sky130_fd_sc_hd__xnor2_2 _17038_ (.A(_09087_),
    .B(_09089_),
    .Y(_09090_));
 sky130_fd_sc_hd__o21a_1 _17039_ (.A1(_09073_),
    .A2(_09074_),
    .B1(_09075_),
    .X(_09091_));
 sky130_fd_sc_hd__xnor2_1 _17040_ (.A(\top0.pid_q.prev_error[15] ),
    .B(\top0.pid_q.curr_error[15] ),
    .Y(_09092_));
 sky130_fd_sc_hd__xnor2_1 _17041_ (.A(_09091_),
    .B(_09092_),
    .Y(_09093_));
 sky130_fd_sc_hd__and2_1 _17042_ (.A(net551),
    .B(_09093_),
    .X(_09094_));
 sky130_fd_sc_hd__a211o_1 _17043_ (.A1(net546),
    .A2(_09090_),
    .B1(_09094_),
    .C1(_08882_),
    .X(_09095_));
 sky130_fd_sc_hd__o211a_1 _17044_ (.A1(net443),
    .A2(_08861_),
    .B1(_09095_),
    .C1(_08930_),
    .X(_00180_));
 sky130_fd_sc_hd__or2_4 _17045_ (.A(net551),
    .B(_08881_),
    .X(_09096_));
 sky130_fd_sc_hd__mux2_1 _17046_ (.A0(_08885_),
    .A1(\top0.pid_q.curr_error[0] ),
    .S(_09096_),
    .X(_09097_));
 sky130_fd_sc_hd__and2_1 _17047_ (.A(net1018),
    .B(_09097_),
    .X(_09098_));
 sky130_fd_sc_hd__clkbuf_1 _17048_ (.A(_09098_),
    .X(_00181_));
 sky130_fd_sc_hd__or2_1 _17049_ (.A(_05448_),
    .B(_08855_),
    .X(_09099_));
 sky130_fd_sc_hd__clkbuf_4 _17050_ (.A(_09099_),
    .X(_09100_));
 sky130_fd_sc_hd__and3b_1 _17051_ (.A_N(net551),
    .B(_00008_),
    .C(_08854_),
    .X(_09101_));
 sky130_fd_sc_hd__clkbuf_4 _17052_ (.A(_09101_),
    .X(_09102_));
 sky130_fd_sc_hd__a22o_1 _17053_ (.A1(net983),
    .A2(_09100_),
    .B1(_09102_),
    .B2(_08894_),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _17054_ (.A0(_08907_),
    .A1(\top0.pid_q.curr_error[2] ),
    .S(_09096_),
    .X(_09103_));
 sky130_fd_sc_hd__and2_1 _17055_ (.A(net1018),
    .B(_09103_),
    .X(_09104_));
 sky130_fd_sc_hd__clkbuf_1 _17056_ (.A(_09104_),
    .X(_00183_));
 sky130_fd_sc_hd__a22o_1 _17057_ (.A1(\top0.pid_q.curr_error[3] ),
    .A2(_09100_),
    .B1(_09102_),
    .B2(_08920_),
    .X(_00184_));
 sky130_fd_sc_hd__a22o_1 _17058_ (.A1(net929),
    .A2(_09100_),
    .B1(_09102_),
    .B2(_08935_),
    .X(_00185_));
 sky130_fd_sc_hd__a22o_1 _17059_ (.A1(\top0.pid_q.curr_error[5] ),
    .A2(_09100_),
    .B1(_09102_),
    .B2(_08949_),
    .X(_00186_));
 sky130_fd_sc_hd__a22o_1 _17060_ (.A1(\top0.pid_q.curr_error[6] ),
    .A2(_09100_),
    .B1(_09102_),
    .B2(_08962_),
    .X(_00187_));
 sky130_fd_sc_hd__a22o_1 _17061_ (.A1(\top0.pid_q.curr_error[7] ),
    .A2(_09100_),
    .B1(_09102_),
    .B2(_08974_),
    .X(_00188_));
 sky130_fd_sc_hd__a22o_1 _17062_ (.A1(\top0.pid_q.curr_error[8] ),
    .A2(_09100_),
    .B1(_09102_),
    .B2(_08987_),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _17063_ (.A0(_09002_),
    .A1(\top0.pid_q.curr_error[9] ),
    .S(_09096_),
    .X(_09105_));
 sky130_fd_sc_hd__and2_1 _17064_ (.A(net1018),
    .B(_09105_),
    .X(_09106_));
 sky130_fd_sc_hd__clkbuf_1 _17065_ (.A(_09106_),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _17066_ (.A0(_09016_),
    .A1(\top0.pid_q.curr_error[10] ),
    .S(_09096_),
    .X(_09107_));
 sky130_fd_sc_hd__and2_1 _17067_ (.A(net1018),
    .B(_09107_),
    .X(_09108_));
 sky130_fd_sc_hd__clkbuf_1 _17068_ (.A(_09108_),
    .X(_00191_));
 sky130_fd_sc_hd__a22o_1 _17069_ (.A1(\top0.pid_q.curr_error[11] ),
    .A2(_09100_),
    .B1(_09102_),
    .B2(_09036_),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _17070_ (.A0(_09045_),
    .A1(\top0.pid_q.curr_error[12] ),
    .S(_09096_),
    .X(_09109_));
 sky130_fd_sc_hd__and2_1 _17071_ (.A(net1018),
    .B(_09109_),
    .X(_09110_));
 sky130_fd_sc_hd__clkbuf_1 _17072_ (.A(_09110_),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _17073_ (.A0(_09063_),
    .A1(\top0.pid_q.curr_error[13] ),
    .S(_09096_),
    .X(_09111_));
 sky130_fd_sc_hd__and2_1 _17074_ (.A(_08403_),
    .B(_09111_),
    .X(_09112_));
 sky130_fd_sc_hd__clkbuf_1 _17075_ (.A(_09112_),
    .X(_00194_));
 sky130_fd_sc_hd__a22o_1 _17076_ (.A1(net865),
    .A2(_09100_),
    .B1(_09102_),
    .B2(_09070_),
    .X(_00195_));
 sky130_fd_sc_hd__a22o_1 _17077_ (.A1(net885),
    .A2(_09100_),
    .B1(_09102_),
    .B2(_09090_),
    .X(_00196_));
 sky130_fd_sc_hd__or2_1 _17078_ (.A(_00008_),
    .B(_08855_),
    .X(_09113_));
 sky130_fd_sc_hd__buf_2 _17079_ (.A(_09113_),
    .X(_09114_));
 sky130_fd_sc_hd__clkbuf_4 _17080_ (.A(_09114_),
    .X(_09115_));
 sky130_fd_sc_hd__nor2_2 _17081_ (.A(_00008_),
    .B(_08855_),
    .Y(_09116_));
 sky130_fd_sc_hd__buf_2 _17082_ (.A(_09116_),
    .X(_09117_));
 sky130_fd_sc_hd__and3_1 _17083_ (.A(\top0.pid_q.curr_error[0] ),
    .B(_00011_),
    .C(_09117_),
    .X(_09118_));
 sky130_fd_sc_hd__a21o_1 _17084_ (.A1(net984),
    .A2(_09115_),
    .B1(_09118_),
    .X(_00197_));
 sky130_fd_sc_hd__and3_1 _17085_ (.A(\top0.pid_q.curr_error[1] ),
    .B(_00011_),
    .C(_09117_),
    .X(_09119_));
 sky130_fd_sc_hd__a21o_1 _17086_ (.A1(\top0.pid_q.prev_error[1] ),
    .A2(_09115_),
    .B1(_09119_),
    .X(_00198_));
 sky130_fd_sc_hd__and3_1 _17087_ (.A(\top0.pid_q.curr_error[2] ),
    .B(_00011_),
    .C(_09117_),
    .X(_09120_));
 sky130_fd_sc_hd__a21o_1 _17088_ (.A1(net897),
    .A2(_09115_),
    .B1(_09120_),
    .X(_00199_));
 sky130_fd_sc_hd__and3_1 _17089_ (.A(\top0.pid_q.curr_error[3] ),
    .B(_00011_),
    .C(_09117_),
    .X(_09121_));
 sky130_fd_sc_hd__a21o_1 _17090_ (.A1(net899),
    .A2(_09115_),
    .B1(_09121_),
    .X(_00200_));
 sky130_fd_sc_hd__and3_1 _17091_ (.A(\top0.pid_q.curr_error[4] ),
    .B(_00011_),
    .C(_09117_),
    .X(_09122_));
 sky130_fd_sc_hd__a21o_1 _17092_ (.A1(net860),
    .A2(_09115_),
    .B1(_09122_),
    .X(_00201_));
 sky130_fd_sc_hd__and3_1 _17093_ (.A(\top0.pid_q.curr_error[5] ),
    .B(_00011_),
    .C(_09117_),
    .X(_09123_));
 sky130_fd_sc_hd__a21o_1 _17094_ (.A1(net849),
    .A2(_09115_),
    .B1(_09123_),
    .X(_00202_));
 sky130_fd_sc_hd__and3_1 _17095_ (.A(\top0.pid_q.curr_error[6] ),
    .B(_00011_),
    .C(_09117_),
    .X(_09124_));
 sky130_fd_sc_hd__a21o_1 _17096_ (.A1(net842),
    .A2(_09115_),
    .B1(_09124_),
    .X(_00203_));
 sky130_fd_sc_hd__and3_1 _17097_ (.A(\top0.pid_q.curr_error[7] ),
    .B(_08860_),
    .C(_09117_),
    .X(_09125_));
 sky130_fd_sc_hd__a21o_1 _17098_ (.A1(net818),
    .A2(_09115_),
    .B1(_09125_),
    .X(_00204_));
 sky130_fd_sc_hd__and3_1 _17099_ (.A(\top0.pid_q.curr_error[8] ),
    .B(_08860_),
    .C(_09117_),
    .X(_09126_));
 sky130_fd_sc_hd__a21o_1 _17100_ (.A1(net812),
    .A2(_09115_),
    .B1(_09126_),
    .X(_00205_));
 sky130_fd_sc_hd__and3_1 _17101_ (.A(\top0.pid_q.curr_error[9] ),
    .B(_08860_),
    .C(_09117_),
    .X(_09127_));
 sky130_fd_sc_hd__a21o_1 _17102_ (.A1(net820),
    .A2(_09115_),
    .B1(_09127_),
    .X(_00206_));
 sky130_fd_sc_hd__and3_1 _17103_ (.A(\top0.pid_q.curr_error[10] ),
    .B(_08860_),
    .C(_09116_),
    .X(_09128_));
 sky130_fd_sc_hd__a21o_1 _17104_ (.A1(net826),
    .A2(_09114_),
    .B1(_09128_),
    .X(_00207_));
 sky130_fd_sc_hd__and3_1 _17105_ (.A(\top0.pid_q.curr_error[11] ),
    .B(_08860_),
    .C(_09116_),
    .X(_09129_));
 sky130_fd_sc_hd__a21o_1 _17106_ (.A1(net898),
    .A2(_09114_),
    .B1(_09129_),
    .X(_00208_));
 sky130_fd_sc_hd__and3_1 _17107_ (.A(\top0.pid_q.curr_error[12] ),
    .B(_08860_),
    .C(_09116_),
    .X(_09130_));
 sky130_fd_sc_hd__a21o_1 _17108_ (.A1(net909),
    .A2(_09114_),
    .B1(_09130_),
    .X(_00209_));
 sky130_fd_sc_hd__and3_1 _17109_ (.A(\top0.pid_q.curr_error[13] ),
    .B(_08860_),
    .C(_09116_),
    .X(_09131_));
 sky130_fd_sc_hd__a21o_1 _17110_ (.A1(net873),
    .A2(_09114_),
    .B1(_09131_),
    .X(_00210_));
 sky130_fd_sc_hd__and3_1 _17111_ (.A(\top0.pid_q.curr_error[14] ),
    .B(_08860_),
    .C(_09116_),
    .X(_09132_));
 sky130_fd_sc_hd__a21o_1 _17112_ (.A1(net728),
    .A2(_09114_),
    .B1(_09132_),
    .X(_00211_));
 sky130_fd_sc_hd__and3_1 _17113_ (.A(\top0.pid_q.curr_error[15] ),
    .B(_08860_),
    .C(_09116_),
    .X(_09133_));
 sky130_fd_sc_hd__a21o_1 _17114_ (.A1(net758),
    .A2(_09114_),
    .B1(_09133_),
    .X(_00212_));
 sky130_fd_sc_hd__nor2_2 _17115_ (.A(net546),
    .B(_08853_),
    .Y(_09134_));
 sky130_fd_sc_hd__o211a_2 _17116_ (.A1(net549),
    .A2(_07698_),
    .B1(_09134_),
    .C1(_05442_),
    .X(_09135_));
 sky130_fd_sc_hd__clkbuf_4 _17117_ (.A(_09135_),
    .X(_09136_));
 sky130_fd_sc_hd__xor2_1 _17118_ (.A(\top0.pid_q.curr_int[0] ),
    .B(\top0.pid_q.prev_int[0] ),
    .X(_09137_));
 sky130_fd_sc_hd__and2b_1 _17119_ (.A_N(_07697_),
    .B(net543),
    .X(_09138_));
 sky130_fd_sc_hd__a211o_1 _17120_ (.A1(net553),
    .A2(_09137_),
    .B1(_09138_),
    .C1(_08887_),
    .X(_09139_));
 sky130_fd_sc_hd__nor2_2 _17121_ (.A(net15),
    .B(_09134_),
    .Y(_09140_));
 sky130_fd_sc_hd__clkbuf_4 _17122_ (.A(_09140_),
    .X(_09141_));
 sky130_fd_sc_hd__a22o_1 _17123_ (.A1(_09136_),
    .A2(_09139_),
    .B1(_09141_),
    .B2(\top0.pid_q.curr_int[0] ),
    .X(_00213_));
 sky130_fd_sc_hd__xor2_1 _17124_ (.A(\top0.pid_q.curr_int[1] ),
    .B(\top0.pid_q.prev_int[1] ),
    .X(_09142_));
 sky130_fd_sc_hd__a21o_1 _17125_ (.A1(\top0.pid_q.curr_int[0] ),
    .A2(\top0.pid_q.prev_int[0] ),
    .B1(_09142_),
    .X(_09143_));
 sky130_fd_sc_hd__nand3_1 _17126_ (.A(\top0.pid_q.curr_int[0] ),
    .B(\top0.pid_q.prev_int[0] ),
    .C(_09142_),
    .Y(_09144_));
 sky130_fd_sc_hd__a32o_1 _17127_ (.A1(net553),
    .A2(_09143_),
    .A3(_09144_),
    .B1(net548),
    .B2(_08897_),
    .X(_09145_));
 sky130_fd_sc_hd__a21o_1 _17128_ (.A1(net543),
    .A2(_07795_),
    .B1(_09145_),
    .X(_09146_));
 sky130_fd_sc_hd__a22o_1 _17129_ (.A1(\top0.pid_q.curr_int[1] ),
    .A2(_09141_),
    .B1(_09146_),
    .B2(_09136_),
    .X(_00214_));
 sky130_fd_sc_hd__nand2_1 _17130_ (.A(\top0.pid_q.curr_int[1] ),
    .B(\top0.pid_q.prev_int[1] ),
    .Y(_09147_));
 sky130_fd_sc_hd__o211ai_2 _17131_ (.A1(\top0.pid_q.curr_int[1] ),
    .A2(\top0.pid_q.prev_int[1] ),
    .B1(\top0.pid_q.prev_int[0] ),
    .C1(\top0.pid_q.curr_int[0] ),
    .Y(_09148_));
 sky130_fd_sc_hd__nand2_1 _17132_ (.A(_09147_),
    .B(_09148_),
    .Y(_09149_));
 sky130_fd_sc_hd__xnor2_1 _17133_ (.A(\top0.pid_q.curr_int[2] ),
    .B(\top0.pid_q.prev_int[2] ),
    .Y(_09150_));
 sky130_fd_sc_hd__xnor2_1 _17134_ (.A(_09149_),
    .B(_09150_),
    .Y(_09151_));
 sky130_fd_sc_hd__a221o_1 _17135_ (.A1(net543),
    .A2(_07895_),
    .B1(_09151_),
    .B2(net553),
    .C1(_08913_),
    .X(_09152_));
 sky130_fd_sc_hd__a22o_1 _17136_ (.A1(\top0.pid_q.curr_int[2] ),
    .A2(_09141_),
    .B1(_09152_),
    .B2(_09136_),
    .X(_00215_));
 sky130_fd_sc_hd__inv_2 _17137_ (.A(\top0.pid_q.prev_int[2] ),
    .Y(_09153_));
 sky130_fd_sc_hd__a21o_1 _17138_ (.A1(_09147_),
    .A2(_09148_),
    .B1(_09153_),
    .X(_09154_));
 sky130_fd_sc_hd__inv_2 _17139_ (.A(\top0.pid_q.curr_int[2] ),
    .Y(_09155_));
 sky130_fd_sc_hd__a31o_1 _17140_ (.A1(_09153_),
    .A2(_09147_),
    .A3(_09148_),
    .B1(_09155_),
    .X(_09156_));
 sky130_fd_sc_hd__and2_1 _17141_ (.A(_09154_),
    .B(_09156_),
    .X(_09157_));
 sky130_fd_sc_hd__xnor2_1 _17142_ (.A(\top0.pid_q.curr_int[3] ),
    .B(\top0.pid_q.prev_int[3] ),
    .Y(_09158_));
 sky130_fd_sc_hd__nand2_1 _17143_ (.A(_09157_),
    .B(_09158_),
    .Y(_09159_));
 sky130_fd_sc_hd__or2_1 _17144_ (.A(_09157_),
    .B(_09158_),
    .X(_09160_));
 sky130_fd_sc_hd__a32o_1 _17145_ (.A1(net553),
    .A2(_09159_),
    .A3(_09160_),
    .B1(net548),
    .B2(_08928_),
    .X(_09161_));
 sky130_fd_sc_hd__a21o_1 _17146_ (.A1(net543),
    .A2(_07991_),
    .B1(_09161_),
    .X(_09162_));
 sky130_fd_sc_hd__a22o_1 _17147_ (.A1(\top0.pid_q.curr_int[3] ),
    .A2(_09141_),
    .B1(_09162_),
    .B2(_09136_),
    .X(_00216_));
 sky130_fd_sc_hd__inv_2 _17148_ (.A(\top0.pid_q.prev_int[3] ),
    .Y(_09163_));
 sky130_fd_sc_hd__a31o_1 _17149_ (.A1(_09163_),
    .A2(_09154_),
    .A3(_09156_),
    .B1(_08076_),
    .X(_09164_));
 sky130_fd_sc_hd__o21ai_2 _17150_ (.A1(_09163_),
    .A2(_09157_),
    .B1(_09164_),
    .Y(_09165_));
 sky130_fd_sc_hd__xor2_1 _17151_ (.A(\top0.pid_q.curr_int[4] ),
    .B(\top0.pid_q.prev_int[4] ),
    .X(_09166_));
 sky130_fd_sc_hd__or2_1 _17152_ (.A(_09165_),
    .B(_09166_),
    .X(_09167_));
 sky130_fd_sc_hd__nand2_1 _17153_ (.A(_09165_),
    .B(_09166_),
    .Y(_09168_));
 sky130_fd_sc_hd__a32o_1 _17154_ (.A1(net553),
    .A2(_09167_),
    .A3(_09168_),
    .B1(net548),
    .B2(_08942_),
    .X(_09169_));
 sky130_fd_sc_hd__a21o_1 _17155_ (.A1(net543),
    .A2(_08075_),
    .B1(_09169_),
    .X(_09170_));
 sky130_fd_sc_hd__a22o_1 _17156_ (.A1(\top0.pid_q.curr_int[4] ),
    .A2(_09141_),
    .B1(_09170_),
    .B2(_09136_),
    .X(_00217_));
 sky130_fd_sc_hd__a21o_1 _17157_ (.A1(\top0.pid_q.prev_int[4] ),
    .A2(_09165_),
    .B1(\top0.pid_q.curr_int[4] ),
    .X(_09171_));
 sky130_fd_sc_hd__o21a_2 _17158_ (.A1(\top0.pid_q.prev_int[4] ),
    .A2(_09165_),
    .B1(_09171_),
    .X(_09172_));
 sky130_fd_sc_hd__xnor2_1 _17159_ (.A(\top0.pid_q.curr_int[5] ),
    .B(\top0.pid_q.prev_int[5] ),
    .Y(_09173_));
 sky130_fd_sc_hd__xnor2_1 _17160_ (.A(_09172_),
    .B(_09173_),
    .Y(_09174_));
 sky130_fd_sc_hd__a221o_1 _17161_ (.A1(net543),
    .A2(_08157_),
    .B1(_09174_),
    .B2(net553),
    .C1(_08955_),
    .X(_09175_));
 sky130_fd_sc_hd__a22o_1 _17162_ (.A1(\top0.pid_q.curr_int[5] ),
    .A2(_09141_),
    .B1(_09175_),
    .B2(_09136_),
    .X(_00218_));
 sky130_fd_sc_hd__nand2_1 _17163_ (.A(_00007_),
    .B(_09134_),
    .Y(_09176_));
 sky130_fd_sc_hd__a21o_1 _17164_ (.A1(\top0.pid_q.prev_int[5] ),
    .A2(_09172_),
    .B1(\top0.pid_q.curr_int[5] ),
    .X(_09177_));
 sky130_fd_sc_hd__o21ai_1 _17165_ (.A1(\top0.pid_q.prev_int[5] ),
    .A2(_09172_),
    .B1(_09177_),
    .Y(_09178_));
 sky130_fd_sc_hd__xnor2_1 _17166_ (.A(\top0.pid_q.curr_int[6] ),
    .B(\top0.pid_q.prev_int[6] ),
    .Y(_09179_));
 sky130_fd_sc_hd__nand2_1 _17167_ (.A(_09178_),
    .B(_09179_),
    .Y(_09180_));
 sky130_fd_sc_hd__or2_1 _17168_ (.A(_09178_),
    .B(_09179_),
    .X(_09181_));
 sky130_fd_sc_hd__a31o_1 _17169_ (.A1(net553),
    .A2(_09180_),
    .A3(_09181_),
    .B1(_08968_),
    .X(_09182_));
 sky130_fd_sc_hd__a22oi_1 _17170_ (.A1(\top0.pid_q.curr_int[6] ),
    .A2(_09141_),
    .B1(_09182_),
    .B2(_09136_),
    .Y(_09183_));
 sky130_fd_sc_hd__o21ai_1 _17171_ (.A1(_08235_),
    .A2(_09176_),
    .B1(_09183_),
    .Y(_00219_));
 sky130_fd_sc_hd__o211a_1 _17172_ (.A1(\top0.pid_q.prev_int[5] ),
    .A2(_09172_),
    .B1(_09177_),
    .C1(\top0.pid_q.prev_int[6] ),
    .X(_09184_));
 sky130_fd_sc_hd__o21a_1 _17173_ (.A1(\top0.pid_q.prev_int[5] ),
    .A2(_09172_),
    .B1(\top0.pid_q.curr_int[5] ),
    .X(_09185_));
 sky130_fd_sc_hd__a211o_1 _17174_ (.A1(\top0.pid_q.prev_int[5] ),
    .A2(_09172_),
    .B1(_09185_),
    .C1(\top0.pid_q.prev_int[6] ),
    .X(_09186_));
 sky130_fd_sc_hd__o21ai_2 _17175_ (.A1(\top0.pid_q.curr_int[6] ),
    .A2(_09184_),
    .B1(_09186_),
    .Y(_09187_));
 sky130_fd_sc_hd__xor2_1 _17176_ (.A(\top0.pid_q.curr_int[7] ),
    .B(\top0.pid_q.prev_int[7] ),
    .X(_09188_));
 sky130_fd_sc_hd__xnor2_1 _17177_ (.A(_09187_),
    .B(_09188_),
    .Y(_09189_));
 sky130_fd_sc_hd__a221o_1 _17178_ (.A1(net543),
    .A2(_08320_),
    .B1(_09189_),
    .B2(net554),
    .C1(_08981_),
    .X(_09190_));
 sky130_fd_sc_hd__a22o_1 _17179_ (.A1(\top0.pid_q.curr_int[7] ),
    .A2(_09141_),
    .B1(_09190_),
    .B2(_09136_),
    .X(_00220_));
 sky130_fd_sc_hd__and3_1 _17180_ (.A(net543),
    .B(_05441_),
    .C(_09134_),
    .X(_09191_));
 sky130_fd_sc_hd__buf_2 _17181_ (.A(_09191_),
    .X(_09192_));
 sky130_fd_sc_hd__inv_2 _17182_ (.A(\top0.pid_q.prev_int[7] ),
    .Y(_09193_));
 sky130_fd_sc_hd__o21a_1 _17183_ (.A1(_09193_),
    .A2(_09187_),
    .B1(_08324_),
    .X(_09194_));
 sky130_fd_sc_hd__a21o_1 _17184_ (.A1(_09193_),
    .A2(_09187_),
    .B1(_09194_),
    .X(_09195_));
 sky130_fd_sc_hd__xnor2_1 _17185_ (.A(\top0.pid_q.curr_int[8] ),
    .B(\top0.pid_q.prev_int[8] ),
    .Y(_09196_));
 sky130_fd_sc_hd__nand2_1 _17186_ (.A(_09195_),
    .B(_09196_),
    .Y(_09197_));
 sky130_fd_sc_hd__or2_1 _17187_ (.A(_09195_),
    .B(_09196_),
    .X(_09198_));
 sky130_fd_sc_hd__a31o_1 _17188_ (.A1(net554),
    .A2(_09197_),
    .A3(_09198_),
    .B1(_08994_),
    .X(_09199_));
 sky130_fd_sc_hd__a22o_1 _17189_ (.A1(\top0.pid_q.curr_int[8] ),
    .A2(_09140_),
    .B1(_09199_),
    .B2(_09135_),
    .X(_09200_));
 sky130_fd_sc_hd__a21o_1 _17190_ (.A1(_08399_),
    .A2(_09192_),
    .B1(_09200_),
    .X(_00221_));
 sky130_fd_sc_hd__inv_2 _17191_ (.A(\top0.pid_q.prev_int[8] ),
    .Y(_09201_));
 sky130_fd_sc_hd__o21ai_1 _17192_ (.A1(_09201_),
    .A2(_09195_),
    .B1(_08404_),
    .Y(_09202_));
 sky130_fd_sc_hd__a21bo_1 _17193_ (.A1(_09201_),
    .A2(_09195_),
    .B1_N(_09202_),
    .X(_09203_));
 sky130_fd_sc_hd__xor2_1 _17194_ (.A(\top0.pid_q.curr_int[9] ),
    .B(\top0.pid_q.prev_int[9] ),
    .X(_09204_));
 sky130_fd_sc_hd__xnor2_1 _17195_ (.A(_09203_),
    .B(_09204_),
    .Y(_09205_));
 sky130_fd_sc_hd__a221o_1 _17196_ (.A1(\top0.pid_q.state[5] ),
    .A2(_08479_),
    .B1(_09205_),
    .B2(net554),
    .C1(_09009_),
    .X(_09206_));
 sky130_fd_sc_hd__a22o_1 _17197_ (.A1(\top0.pid_q.curr_int[9] ),
    .A2(_09141_),
    .B1(_09206_),
    .B2(_09136_),
    .X(_00222_));
 sky130_fd_sc_hd__inv_2 _17198_ (.A(\top0.pid_q.prev_int[9] ),
    .Y(_09207_));
 sky130_fd_sc_hd__a21bo_1 _17199_ (.A1(_09207_),
    .A2(_09203_),
    .B1_N(\top0.pid_q.curr_int[9] ),
    .X(_09208_));
 sky130_fd_sc_hd__o21a_1 _17200_ (.A1(_09207_),
    .A2(_09203_),
    .B1(_09208_),
    .X(_09209_));
 sky130_fd_sc_hd__xnor2_1 _17201_ (.A(\top0.pid_q.curr_int[10] ),
    .B(\top0.pid_q.prev_int[10] ),
    .Y(_09210_));
 sky130_fd_sc_hd__nand2_1 _17202_ (.A(_09209_),
    .B(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__or2_1 _17203_ (.A(_09209_),
    .B(_09210_),
    .X(_09212_));
 sky130_fd_sc_hd__a31o_1 _17204_ (.A1(net554),
    .A2(_09211_),
    .A3(_09212_),
    .B1(_09023_),
    .X(_09213_));
 sky130_fd_sc_hd__a22o_1 _17205_ (.A1(\top0.pid_q.curr_int[10] ),
    .A2(_09140_),
    .B1(_09213_),
    .B2(_09135_),
    .X(_09214_));
 sky130_fd_sc_hd__a21o_1 _17206_ (.A1(_08550_),
    .A2(_09192_),
    .B1(_09214_),
    .X(_00223_));
 sky130_fd_sc_hd__inv_2 _17207_ (.A(\top0.pid_q.prev_int[10] ),
    .Y(_09215_));
 sky130_fd_sc_hd__o21ba_1 _17208_ (.A1(_09215_),
    .A2(_09209_),
    .B1_N(\top0.pid_q.curr_int[10] ),
    .X(_09216_));
 sky130_fd_sc_hd__a21oi_1 _17209_ (.A1(_09215_),
    .A2(_09209_),
    .B1(_09216_),
    .Y(_09217_));
 sky130_fd_sc_hd__xnor2_1 _17210_ (.A(\top0.pid_q.curr_int[11] ),
    .B(\top0.pid_q.prev_int[11] ),
    .Y(_09218_));
 sky130_fd_sc_hd__xnor2_1 _17211_ (.A(_09217_),
    .B(_09218_),
    .Y(_09219_));
 sky130_fd_sc_hd__a22o_1 _17212_ (.A1(net548),
    .A2(_09029_),
    .B1(_09219_),
    .B2(net554),
    .X(_09220_));
 sky130_fd_sc_hd__nor2_1 _17213_ (.A(_08609_),
    .B(_09176_),
    .Y(_09221_));
 sky130_fd_sc_hd__a221o_1 _17214_ (.A1(\top0.pid_q.curr_int[11] ),
    .A2(_09141_),
    .B1(_09220_),
    .B2(_09136_),
    .C1(_09221_),
    .X(_00224_));
 sky130_fd_sc_hd__inv_2 _17215_ (.A(_08685_),
    .Y(_09222_));
 sky130_fd_sc_hd__or2_1 _17216_ (.A(\top0.pid_q.curr_int[11] ),
    .B(\top0.pid_q.prev_int[11] ),
    .X(_09223_));
 sky130_fd_sc_hd__and2_1 _17217_ (.A(\top0.pid_q.curr_int[11] ),
    .B(\top0.pid_q.prev_int[11] ),
    .X(_09224_));
 sky130_fd_sc_hd__a21o_1 _17218_ (.A1(_09217_),
    .A2(_09223_),
    .B1(_09224_),
    .X(_09225_));
 sky130_fd_sc_hd__xnor2_1 _17219_ (.A(\top0.pid_q.curr_int[12] ),
    .B(\top0.pid_q.prev_int[12] ),
    .Y(_09226_));
 sky130_fd_sc_hd__xnor2_1 _17220_ (.A(_09225_),
    .B(_09226_),
    .Y(_09227_));
 sky130_fd_sc_hd__a22o_1 _17221_ (.A1(net551),
    .A2(_09050_),
    .B1(_09227_),
    .B2(net553),
    .X(_09228_));
 sky130_fd_sc_hd__a22o_1 _17222_ (.A1(\top0.pid_q.curr_int[12] ),
    .A2(_09140_),
    .B1(_09192_),
    .B2(_08679_),
    .X(_09229_));
 sky130_fd_sc_hd__a221o_1 _17223_ (.A1(_09222_),
    .A2(_09192_),
    .B1(_09228_),
    .B2(_09135_),
    .C1(_09229_),
    .X(_00225_));
 sky130_fd_sc_hd__o21a_1 _17224_ (.A1(\top0.pid_q.curr_int[12] ),
    .A2(\top0.pid_q.prev_int[12] ),
    .B1(_09225_),
    .X(_09230_));
 sky130_fd_sc_hd__a21o_1 _17225_ (.A1(\top0.pid_q.curr_int[12] ),
    .A2(\top0.pid_q.prev_int[12] ),
    .B1(_09230_),
    .X(_09231_));
 sky130_fd_sc_hd__xnor2_1 _17226_ (.A(\top0.pid_q.curr_int[13] ),
    .B(\top0.pid_q.prev_int[13] ),
    .Y(_09232_));
 sky130_fd_sc_hd__xnor2_1 _17227_ (.A(_09231_),
    .B(_09232_),
    .Y(_09233_));
 sky130_fd_sc_hd__a22o_1 _17228_ (.A1(net551),
    .A2(_09055_),
    .B1(_09233_),
    .B2(net554),
    .X(_09234_));
 sky130_fd_sc_hd__a22o_1 _17229_ (.A1(\top0.pid_q.curr_int[13] ),
    .A2(_09140_),
    .B1(_09234_),
    .B2(_09135_),
    .X(_09235_));
 sky130_fd_sc_hd__a21o_1 _17230_ (.A1(_08738_),
    .A2(_09192_),
    .B1(_09235_),
    .X(_00226_));
 sky130_fd_sc_hd__or2_1 _17231_ (.A(net546),
    .B(_08853_),
    .X(_09236_));
 sky130_fd_sc_hd__nor2_1 _17232_ (.A(\top0.pid_q.curr_int[14] ),
    .B(_09236_),
    .Y(_09237_));
 sky130_fd_sc_hd__a21o_1 _17233_ (.A1(\top0.pid_q.prev_int[13] ),
    .A2(_09231_),
    .B1(\top0.pid_q.curr_int[13] ),
    .X(_09238_));
 sky130_fd_sc_hd__o21ai_1 _17234_ (.A1(\top0.pid_q.prev_int[13] ),
    .A2(_09231_),
    .B1(_09238_),
    .Y(_09239_));
 sky130_fd_sc_hd__xnor2_1 _17235_ (.A(\top0.pid_q.prev_int[14] ),
    .B(_09239_),
    .Y(_09240_));
 sky130_fd_sc_hd__mux2_1 _17236_ (.A0(\top0.pid_q.curr_int[14] ),
    .A1(_09237_),
    .S(_09240_),
    .X(_09241_));
 sky130_fd_sc_hd__a22o_1 _17237_ (.A1(\top0.pid_q.curr_int[14] ),
    .A2(_09236_),
    .B1(_09241_),
    .B2(net554),
    .X(_09242_));
 sky130_fd_sc_hd__and3_1 _17238_ (.A(net551),
    .B(_09077_),
    .C(_09135_),
    .X(_09243_));
 sky130_fd_sc_hd__a221o_1 _17239_ (.A1(_08791_),
    .A2(_09192_),
    .B1(_09242_),
    .B2(net1019),
    .C1(_09243_),
    .X(_00227_));
 sky130_fd_sc_hd__nand2_1 _17240_ (.A(\top0.pid_q.curr_int[14] ),
    .B(\top0.pid_q.prev_int[14] ),
    .Y(_09244_));
 sky130_fd_sc_hd__nor2_1 _17241_ (.A(\top0.pid_q.curr_int[14] ),
    .B(\top0.pid_q.prev_int[14] ),
    .Y(_09245_));
 sky130_fd_sc_hd__a21oi_1 _17242_ (.A1(_09239_),
    .A2(_09244_),
    .B1(_09245_),
    .Y(_09246_));
 sky130_fd_sc_hd__xnor2_1 _17243_ (.A(\top0.pid_q.curr_int[15] ),
    .B(\top0.pid_q.prev_int[15] ),
    .Y(_09247_));
 sky130_fd_sc_hd__xnor2_1 _17244_ (.A(_09246_),
    .B(_09247_),
    .Y(_09248_));
 sky130_fd_sc_hd__a22o_1 _17245_ (.A1(\top0.pid_q.curr_int[15] ),
    .A2(_09140_),
    .B1(_09192_),
    .B2(_08849_),
    .X(_09249_));
 sky130_fd_sc_hd__a41o_1 _17246_ (.A1(net554),
    .A2(_05443_),
    .A3(_09134_),
    .A4(_09248_),
    .B1(_09249_),
    .X(_09250_));
 sky130_fd_sc_hd__a221o_1 _17247_ (.A1(_09094_),
    .A2(_09135_),
    .B1(_09192_),
    .B2(_08842_),
    .C1(_09250_),
    .X(_00228_));
 sky130_fd_sc_hd__xor2_1 _17248_ (.A(\top0.matmul0.matmul_stage_inst.mult1[0] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[0] ),
    .X(_09251_));
 sky130_fd_sc_hd__mux2_1 _17249_ (.A0(\top0.matmul0.beta_pass[0] ),
    .A1(_09251_),
    .S(net563),
    .X(_09252_));
 sky130_fd_sc_hd__clkbuf_1 _17250_ (.A(_09252_),
    .X(_00229_));
 sky130_fd_sc_hd__nand2_1 _17251_ (.A(\top0.matmul0.matmul_stage_inst.mult1[0] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[0] ),
    .Y(_09253_));
 sky130_fd_sc_hd__xor2_1 _17252_ (.A(\top0.matmul0.matmul_stage_inst.mult1[1] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[1] ),
    .X(_09254_));
 sky130_fd_sc_hd__xnor2_1 _17253_ (.A(_09253_),
    .B(_09254_),
    .Y(_09255_));
 sky130_fd_sc_hd__mux2_1 _17254_ (.A0(\top0.matmul0.beta_pass[1] ),
    .A1(_09255_),
    .S(net563),
    .X(_09256_));
 sky130_fd_sc_hd__clkbuf_1 _17255_ (.A(_09256_),
    .X(_00230_));
 sky130_fd_sc_hd__a21o_1 _17256_ (.A1(\top0.matmul0.matmul_stage_inst.mult1[0] ),
    .A2(\top0.matmul0.matmul_stage_inst.mult2[0] ),
    .B1(\top0.matmul0.matmul_stage_inst.mult2[1] ),
    .X(_09257_));
 sky130_fd_sc_hd__a31o_1 _17257_ (.A1(\top0.matmul0.matmul_stage_inst.mult2[1] ),
    .A2(\top0.matmul0.matmul_stage_inst.mult1[0] ),
    .A3(\top0.matmul0.matmul_stage_inst.mult2[0] ),
    .B1(\top0.matmul0.matmul_stage_inst.mult1[1] ),
    .X(_09258_));
 sky130_fd_sc_hd__nand2_1 _17258_ (.A(_09257_),
    .B(_09258_),
    .Y(_09259_));
 sky130_fd_sc_hd__xor2_1 _17259_ (.A(\top0.matmul0.matmul_stage_inst.mult1[2] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[2] ),
    .X(_09260_));
 sky130_fd_sc_hd__xnor2_1 _17260_ (.A(_09259_),
    .B(_09260_),
    .Y(_09261_));
 sky130_fd_sc_hd__mux2_1 _17261_ (.A0(\top0.matmul0.beta_pass[2] ),
    .A1(_09261_),
    .S(net563),
    .X(_09262_));
 sky130_fd_sc_hd__clkbuf_1 _17262_ (.A(_09262_),
    .X(_00231_));
 sky130_fd_sc_hd__inv_2 _17263_ (.A(\top0.matmul0.matmul_stage_inst.mult2[2] ),
    .Y(_09263_));
 sky130_fd_sc_hd__a31o_1 _17264_ (.A1(\top0.matmul0.matmul_stage_inst.mult2[2] ),
    .A2(_09257_),
    .A3(_09258_),
    .B1(\top0.matmul0.matmul_stage_inst.mult1[2] ),
    .X(_09264_));
 sky130_fd_sc_hd__a21boi_2 _17265_ (.A1(_09263_),
    .A2(_09259_),
    .B1_N(_09264_),
    .Y(_09265_));
 sky130_fd_sc_hd__xnor2_1 _17266_ (.A(\top0.matmul0.matmul_stage_inst.mult1[3] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[3] ),
    .Y(_09266_));
 sky130_fd_sc_hd__xnor2_1 _17267_ (.A(_09265_),
    .B(_09266_),
    .Y(_09267_));
 sky130_fd_sc_hd__mux2_1 _17268_ (.A0(\top0.matmul0.beta_pass[3] ),
    .A1(_09267_),
    .S(net563),
    .X(_09268_));
 sky130_fd_sc_hd__clkbuf_1 _17269_ (.A(_09268_),
    .X(_00232_));
 sky130_fd_sc_hd__a21o_1 _17270_ (.A1(\top0.matmul0.matmul_stage_inst.mult2[3] ),
    .A2(_09265_),
    .B1(\top0.matmul0.matmul_stage_inst.mult1[3] ),
    .X(_09269_));
 sky130_fd_sc_hd__o21ai_2 _17271_ (.A1(\top0.matmul0.matmul_stage_inst.mult2[3] ),
    .A2(_09265_),
    .B1(_09269_),
    .Y(_09270_));
 sky130_fd_sc_hd__xor2_1 _17272_ (.A(\top0.matmul0.matmul_stage_inst.mult1[4] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[4] ),
    .X(_09271_));
 sky130_fd_sc_hd__xnor2_1 _17273_ (.A(_09270_),
    .B(_09271_),
    .Y(_09272_));
 sky130_fd_sc_hd__mux2_1 _17274_ (.A0(\top0.matmul0.beta_pass[4] ),
    .A1(_09272_),
    .S(net562),
    .X(_09273_));
 sky130_fd_sc_hd__clkbuf_1 _17275_ (.A(_09273_),
    .X(_00233_));
 sky130_fd_sc_hd__inv_2 _17276_ (.A(\top0.matmul0.matmul_stage_inst.mult2[4] ),
    .Y(_09274_));
 sky130_fd_sc_hd__o21ba_1 _17277_ (.A1(_09274_),
    .A2(_09270_),
    .B1_N(\top0.matmul0.matmul_stage_inst.mult1[4] ),
    .X(_09275_));
 sky130_fd_sc_hd__a21o_1 _17278_ (.A1(_09274_),
    .A2(_09270_),
    .B1(_09275_),
    .X(_09276_));
 sky130_fd_sc_hd__xor2_1 _17279_ (.A(\top0.matmul0.matmul_stage_inst.mult1[5] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[5] ),
    .X(_09277_));
 sky130_fd_sc_hd__xnor2_1 _17280_ (.A(_09276_),
    .B(_09277_),
    .Y(_09278_));
 sky130_fd_sc_hd__mux2_1 _17281_ (.A0(\top0.matmul0.beta_pass[5] ),
    .A1(_09278_),
    .S(net562),
    .X(_09279_));
 sky130_fd_sc_hd__clkbuf_1 _17282_ (.A(_09279_),
    .X(_00234_));
 sky130_fd_sc_hd__inv_2 _17283_ (.A(\top0.matmul0.matmul_stage_inst.mult2[5] ),
    .Y(_09280_));
 sky130_fd_sc_hd__o21ba_1 _17284_ (.A1(_09280_),
    .A2(_09276_),
    .B1_N(\top0.matmul0.matmul_stage_inst.mult1[5] ),
    .X(_09281_));
 sky130_fd_sc_hd__a21o_1 _17285_ (.A1(_09280_),
    .A2(_09276_),
    .B1(_09281_),
    .X(_09282_));
 sky130_fd_sc_hd__xor2_1 _17286_ (.A(\top0.matmul0.matmul_stage_inst.mult1[6] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[6] ),
    .X(_09283_));
 sky130_fd_sc_hd__xnor2_1 _17287_ (.A(_09282_),
    .B(_09283_),
    .Y(_09284_));
 sky130_fd_sc_hd__mux2_1 _17288_ (.A0(\top0.matmul0.beta_pass[6] ),
    .A1(_09284_),
    .S(net562),
    .X(_09285_));
 sky130_fd_sc_hd__clkbuf_1 _17289_ (.A(_09285_),
    .X(_00235_));
 sky130_fd_sc_hd__inv_2 _17290_ (.A(\top0.matmul0.matmul_stage_inst.mult2[6] ),
    .Y(_09286_));
 sky130_fd_sc_hd__a21bo_1 _17291_ (.A1(_09286_),
    .A2(_09282_),
    .B1_N(\top0.matmul0.matmul_stage_inst.mult1[6] ),
    .X(_09287_));
 sky130_fd_sc_hd__o21a_1 _17292_ (.A1(_09286_),
    .A2(_09282_),
    .B1(_09287_),
    .X(_09288_));
 sky130_fd_sc_hd__xor2_1 _17293_ (.A(\top0.matmul0.matmul_stage_inst.mult1[7] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[7] ),
    .X(_09289_));
 sky130_fd_sc_hd__xnor2_1 _17294_ (.A(_09288_),
    .B(_09289_),
    .Y(_09290_));
 sky130_fd_sc_hd__mux2_1 _17295_ (.A0(\top0.matmul0.beta_pass[7] ),
    .A1(_09290_),
    .S(net563),
    .X(_09291_));
 sky130_fd_sc_hd__clkbuf_1 _17296_ (.A(_09291_),
    .X(_00236_));
 sky130_fd_sc_hd__inv_2 _17297_ (.A(\top0.matmul0.matmul_stage_inst.mult2[7] ),
    .Y(_09292_));
 sky130_fd_sc_hd__o21ba_1 _17298_ (.A1(_09292_),
    .A2(_09288_),
    .B1_N(\top0.matmul0.matmul_stage_inst.mult1[7] ),
    .X(_09293_));
 sky130_fd_sc_hd__a21o_1 _17299_ (.A1(_09292_),
    .A2(_09288_),
    .B1(_09293_),
    .X(_09294_));
 sky130_fd_sc_hd__xor2_1 _17300_ (.A(\top0.matmul0.matmul_stage_inst.mult1[8] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[8] ),
    .X(_09295_));
 sky130_fd_sc_hd__xnor2_1 _17301_ (.A(_09294_),
    .B(_09295_),
    .Y(_09296_));
 sky130_fd_sc_hd__mux2_1 _17302_ (.A0(\top0.matmul0.beta_pass[8] ),
    .A1(_09296_),
    .S(net562),
    .X(_09297_));
 sky130_fd_sc_hd__clkbuf_1 _17303_ (.A(_09297_),
    .X(_00237_));
 sky130_fd_sc_hd__inv_2 _17304_ (.A(\top0.matmul0.matmul_stage_inst.mult2[8] ),
    .Y(_09298_));
 sky130_fd_sc_hd__o21ba_1 _17305_ (.A1(_09298_),
    .A2(_09294_),
    .B1_N(\top0.matmul0.matmul_stage_inst.mult1[8] ),
    .X(_09299_));
 sky130_fd_sc_hd__a21o_1 _17306_ (.A1(_09298_),
    .A2(_09294_),
    .B1(_09299_),
    .X(_09300_));
 sky130_fd_sc_hd__xor2_1 _17307_ (.A(\top0.matmul0.matmul_stage_inst.mult1[9] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[9] ),
    .X(_09301_));
 sky130_fd_sc_hd__xnor2_1 _17308_ (.A(_09300_),
    .B(_09301_),
    .Y(_09302_));
 sky130_fd_sc_hd__mux2_1 _17309_ (.A0(\top0.matmul0.beta_pass[9] ),
    .A1(_09302_),
    .S(net562),
    .X(_09303_));
 sky130_fd_sc_hd__clkbuf_1 _17310_ (.A(_09303_),
    .X(_00238_));
 sky130_fd_sc_hd__inv_2 _17311_ (.A(\top0.matmul0.matmul_stage_inst.mult2[9] ),
    .Y(_09304_));
 sky130_fd_sc_hd__o21ba_1 _17312_ (.A1(_09304_),
    .A2(_09300_),
    .B1_N(\top0.matmul0.matmul_stage_inst.mult1[9] ),
    .X(_09305_));
 sky130_fd_sc_hd__a21o_1 _17313_ (.A1(_09304_),
    .A2(_09300_),
    .B1(_09305_),
    .X(_09306_));
 sky130_fd_sc_hd__xor2_1 _17314_ (.A(\top0.matmul0.matmul_stage_inst.mult1[10] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[10] ),
    .X(_09307_));
 sky130_fd_sc_hd__xnor2_1 _17315_ (.A(_09306_),
    .B(_09307_),
    .Y(_09308_));
 sky130_fd_sc_hd__mux2_1 _17316_ (.A0(net430),
    .A1(_09308_),
    .S(net562),
    .X(_09309_));
 sky130_fd_sc_hd__clkbuf_1 _17317_ (.A(_09309_),
    .X(_00239_));
 sky130_fd_sc_hd__inv_2 _17318_ (.A(\top0.matmul0.matmul_stage_inst.mult2[10] ),
    .Y(_09310_));
 sky130_fd_sc_hd__o21ba_1 _17319_ (.A1(_09310_),
    .A2(_09306_),
    .B1_N(\top0.matmul0.matmul_stage_inst.mult1[10] ),
    .X(_09311_));
 sky130_fd_sc_hd__a21o_1 _17320_ (.A1(_09310_),
    .A2(_09306_),
    .B1(_09311_),
    .X(_09312_));
 sky130_fd_sc_hd__xor2_1 _17321_ (.A(\top0.matmul0.matmul_stage_inst.mult1[11] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[11] ),
    .X(_09313_));
 sky130_fd_sc_hd__xnor2_2 _17322_ (.A(_09312_),
    .B(_09313_),
    .Y(_09314_));
 sky130_fd_sc_hd__mux2_1 _17323_ (.A0(\top0.matmul0.beta_pass[11] ),
    .A1(_09314_),
    .S(net562),
    .X(_09315_));
 sky130_fd_sc_hd__clkbuf_1 _17324_ (.A(_09315_),
    .X(_00240_));
 sky130_fd_sc_hd__nand2_1 _17325_ (.A(\top0.matmul0.matmul_stage_inst.mult1[11] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[11] ),
    .Y(_09316_));
 sky130_fd_sc_hd__nor2_1 _17326_ (.A(\top0.matmul0.matmul_stage_inst.mult1[11] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[11] ),
    .Y(_09317_));
 sky130_fd_sc_hd__a21oi_2 _17327_ (.A1(_09312_),
    .A2(_09316_),
    .B1(_09317_),
    .Y(_09318_));
 sky130_fd_sc_hd__xnor2_1 _17328_ (.A(\top0.matmul0.matmul_stage_inst.mult1[12] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[12] ),
    .Y(_09319_));
 sky130_fd_sc_hd__xnor2_2 _17329_ (.A(_09318_),
    .B(_09319_),
    .Y(_09320_));
 sky130_fd_sc_hd__mux2_1 _17330_ (.A0(\top0.matmul0.beta_pass[12] ),
    .A1(_09320_),
    .S(net562),
    .X(_09321_));
 sky130_fd_sc_hd__clkbuf_1 _17331_ (.A(_09321_),
    .X(_00241_));
 sky130_fd_sc_hd__a21o_1 _17332_ (.A1(\top0.matmul0.matmul_stage_inst.mult2[12] ),
    .A2(_09318_),
    .B1(\top0.matmul0.matmul_stage_inst.mult1[12] ),
    .X(_09322_));
 sky130_fd_sc_hd__o21ai_2 _17333_ (.A1(\top0.matmul0.matmul_stage_inst.mult2[12] ),
    .A2(_09318_),
    .B1(_09322_),
    .Y(_09323_));
 sky130_fd_sc_hd__xor2_1 _17334_ (.A(\top0.matmul0.matmul_stage_inst.mult1[13] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[13] ),
    .X(_09324_));
 sky130_fd_sc_hd__xnor2_2 _17335_ (.A(_09323_),
    .B(_09324_),
    .Y(_09325_));
 sky130_fd_sc_hd__mux2_1 _17336_ (.A0(\top0.matmul0.beta_pass[13] ),
    .A1(_09325_),
    .S(net563),
    .X(_09326_));
 sky130_fd_sc_hd__clkbuf_1 _17337_ (.A(_09326_),
    .X(_00242_));
 sky130_fd_sc_hd__nand2_1 _17338_ (.A(\top0.matmul0.matmul_stage_inst.mult1[13] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[13] ),
    .Y(_09327_));
 sky130_fd_sc_hd__nor2_1 _17339_ (.A(\top0.matmul0.matmul_stage_inst.mult1[13] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[13] ),
    .Y(_09328_));
 sky130_fd_sc_hd__a21o_1 _17340_ (.A1(_09323_),
    .A2(_09327_),
    .B1(_09328_),
    .X(_09329_));
 sky130_fd_sc_hd__xor2_1 _17341_ (.A(\top0.matmul0.matmul_stage_inst.mult1[14] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[14] ),
    .X(_09330_));
 sky130_fd_sc_hd__xnor2_2 _17342_ (.A(_09329_),
    .B(_09330_),
    .Y(_09331_));
 sky130_fd_sc_hd__mux2_1 _17343_ (.A0(\top0.matmul0.beta_pass[14] ),
    .A1(_09331_),
    .S(net562),
    .X(_09332_));
 sky130_fd_sc_hd__clkbuf_1 _17344_ (.A(_09332_),
    .X(_00243_));
 sky130_fd_sc_hd__xor2_1 _17345_ (.A(\top0.matmul0.matmul_stage_inst.mult1[15] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[15] ),
    .X(_09333_));
 sky130_fd_sc_hd__nor2_1 _17346_ (.A(\top0.matmul0.matmul_stage_inst.mult1[14] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[14] ),
    .Y(_09334_));
 sky130_fd_sc_hd__nand2_1 _17347_ (.A(\top0.matmul0.matmul_stage_inst.mult1[14] ),
    .B(\top0.matmul0.matmul_stage_inst.mult2[14] ),
    .Y(_09335_));
 sky130_fd_sc_hd__o21a_1 _17348_ (.A1(_09329_),
    .A2(_09334_),
    .B1(_09335_),
    .X(_09336_));
 sky130_fd_sc_hd__xnor2_2 _17349_ (.A(_09333_),
    .B(_09336_),
    .Y(_09337_));
 sky130_fd_sc_hd__mux2_1 _17350_ (.A0(\top0.matmul0.beta_pass[15] ),
    .A1(_09337_),
    .S(net562),
    .X(_09338_));
 sky130_fd_sc_hd__clkbuf_1 _17351_ (.A(_09338_),
    .X(_00244_));
 sky130_fd_sc_hd__clkbuf_4 _17352_ (.A(_07141_),
    .X(_09339_));
 sky130_fd_sc_hd__nand2_1 _17353_ (.A(net418),
    .B(net344),
    .Y(_09340_));
 sky130_fd_sc_hd__nand2_1 _17354_ (.A(net423),
    .B(net340),
    .Y(_09341_));
 sky130_fd_sc_hd__nand2_1 _17355_ (.A(net415),
    .B(net348),
    .Y(_09342_));
 sky130_fd_sc_hd__o21ai_1 _17356_ (.A1(_09340_),
    .A2(_09341_),
    .B1(_09342_),
    .Y(_09343_));
 sky130_fd_sc_hd__a21bo_1 _17357_ (.A1(_09340_),
    .A2(_09341_),
    .B1_N(_09343_),
    .X(_09344_));
 sky130_fd_sc_hd__nand2_1 _17358_ (.A(net417),
    .B(net343),
    .Y(_09345_));
 sky130_fd_sc_hd__nand2_1 _17359_ (.A(net412),
    .B(net347),
    .Y(_09346_));
 sky130_fd_sc_hd__nand2_1 _17360_ (.A(net418),
    .B(net340),
    .Y(_09347_));
 sky130_fd_sc_hd__xnor2_1 _17361_ (.A(_09346_),
    .B(_09347_),
    .Y(_09348_));
 sky130_fd_sc_hd__xnor2_2 _17362_ (.A(_09345_),
    .B(_09348_),
    .Y(_09349_));
 sky130_fd_sc_hd__nor2_1 _17363_ (.A(_09344_),
    .B(_09349_),
    .Y(_09350_));
 sky130_fd_sc_hd__inv_2 _17364_ (.A(net396),
    .Y(_09351_));
 sky130_fd_sc_hd__inv_2 _17365_ (.A(net400),
    .Y(_09352_));
 sky130_fd_sc_hd__clkbuf_4 _17366_ (.A(_09352_),
    .X(_09353_));
 sky130_fd_sc_hd__nor2_1 _17367_ (.A(net407),
    .B(_09353_),
    .Y(_09354_));
 sky130_fd_sc_hd__inv_2 _17368_ (.A(net353),
    .Y(_09355_));
 sky130_fd_sc_hd__buf_4 _17369_ (.A(_09355_),
    .X(_09356_));
 sky130_fd_sc_hd__nor2_1 _17370_ (.A(_09351_),
    .B(_09356_),
    .Y(_09357_));
 sky130_fd_sc_hd__a22o_1 _17371_ (.A1(net405),
    .A2(_09351_),
    .B1(_09354_),
    .B2(_09357_),
    .X(_09358_));
 sky130_fd_sc_hd__nand2_1 _17372_ (.A(net400),
    .B(net353),
    .Y(_09359_));
 sky130_fd_sc_hd__nand2_2 _17373_ (.A(net395),
    .B(net357),
    .Y(_09360_));
 sky130_fd_sc_hd__a22oi_2 _17374_ (.A1(net357),
    .A2(_09358_),
    .B1(_09359_),
    .B2(_09360_),
    .Y(_09361_));
 sky130_fd_sc_hd__nand2_1 _17375_ (.A(net354),
    .B(net358),
    .Y(_09362_));
 sky130_fd_sc_hd__buf_2 _17376_ (.A(_09362_),
    .X(_09363_));
 sky130_fd_sc_hd__clkbuf_4 _17377_ (.A(_09363_),
    .X(_09364_));
 sky130_fd_sc_hd__nand2_1 _17378_ (.A(net410),
    .B(net405),
    .Y(_09365_));
 sky130_fd_sc_hd__nor2_1 _17379_ (.A(_09364_),
    .B(_09365_),
    .Y(_09366_));
 sky130_fd_sc_hd__a22o_1 _17380_ (.A1(_09350_),
    .A2(_09361_),
    .B1(_09366_),
    .B2(_09353_),
    .X(_09367_));
 sky130_fd_sc_hd__o21ai_2 _17381_ (.A1(_09350_),
    .A2(_09361_),
    .B1(_09367_),
    .Y(_09368_));
 sky130_fd_sc_hd__nand2_1 _17382_ (.A(net417),
    .B(net340),
    .Y(_09369_));
 sky130_fd_sc_hd__nand2_1 _17383_ (.A(net412),
    .B(net343),
    .Y(_09370_));
 sky130_fd_sc_hd__nand2_1 _17384_ (.A(net408),
    .B(net347),
    .Y(_09371_));
 sky130_fd_sc_hd__xnor2_1 _17385_ (.A(_09370_),
    .B(_09371_),
    .Y(_09372_));
 sky130_fd_sc_hd__xnor2_2 _17386_ (.A(_09369_),
    .B(_09372_),
    .Y(_09373_));
 sky130_fd_sc_hd__o21a_1 _17387_ (.A1(_09346_),
    .A2(_09347_),
    .B1(_09345_),
    .X(_09374_));
 sky130_fd_sc_hd__a21oi_2 _17388_ (.A1(_09346_),
    .A2(_09347_),
    .B1(_09374_),
    .Y(_09375_));
 sky130_fd_sc_hd__xnor2_1 _17389_ (.A(_09373_),
    .B(_09375_),
    .Y(_09376_));
 sky130_fd_sc_hd__and2_1 _17390_ (.A(net334),
    .B(net338),
    .X(_09377_));
 sky130_fd_sc_hd__and3_1 _17391_ (.A(net423),
    .B(\top0.pid_d.mult0.a[0] ),
    .C(_09377_),
    .X(_09378_));
 sky130_fd_sc_hd__buf_2 _17392_ (.A(_09378_),
    .X(_09379_));
 sky130_fd_sc_hd__nand2_1 _17393_ (.A(net419),
    .B(net337),
    .Y(_09380_));
 sky130_fd_sc_hd__nand2_1 _17394_ (.A(net330),
    .B(net427),
    .Y(_09381_));
 sky130_fd_sc_hd__nand2_1 _17395_ (.A(net333),
    .B(net422),
    .Y(_09382_));
 sky130_fd_sc_hd__xor2_1 _17396_ (.A(_09381_),
    .B(_09382_),
    .X(_09383_));
 sky130_fd_sc_hd__xnor2_2 _17397_ (.A(_09380_),
    .B(_09383_),
    .Y(_09384_));
 sky130_fd_sc_hd__xnor2_1 _17398_ (.A(_09379_),
    .B(_09384_),
    .Y(_09385_));
 sky130_fd_sc_hd__xnor2_1 _17399_ (.A(_09376_),
    .B(_09385_),
    .Y(_09386_));
 sky130_fd_sc_hd__nand2_1 _17400_ (.A(net334),
    .B(\top0.pid_d.mult0.a[0] ),
    .Y(_09387_));
 sky130_fd_sc_hd__nand2_1 _17401_ (.A(net338),
    .B(net423),
    .Y(_09388_));
 sky130_fd_sc_hd__xnor2_1 _17402_ (.A(_09387_),
    .B(_09388_),
    .Y(_09389_));
 sky130_fd_sc_hd__a21oi_1 _17403_ (.A1(_09344_),
    .A2(_09349_),
    .B1(_09389_),
    .Y(_09390_));
 sky130_fd_sc_hd__nor2_1 _17404_ (.A(_09386_),
    .B(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__nor2_1 _17405_ (.A(_09350_),
    .B(_09390_),
    .Y(_09392_));
 sky130_fd_sc_hd__or2b_1 _17406_ (.A(_09392_),
    .B_N(_09386_),
    .X(_09393_));
 sky130_fd_sc_hd__inv_2 _17407_ (.A(net357),
    .Y(_09394_));
 sky130_fd_sc_hd__buf_4 _17408_ (.A(_09394_),
    .X(_09395_));
 sky130_fd_sc_hd__and4_1 _17409_ (.A(net410),
    .B(_09352_),
    .C(_09351_),
    .D(net357),
    .X(_09396_));
 sky130_fd_sc_hd__a21o_1 _17410_ (.A1(net400),
    .A2(net395),
    .B1(_09396_),
    .X(_09397_));
 sky130_fd_sc_hd__a22o_1 _17411_ (.A1(net400),
    .A2(_09395_),
    .B1(_09397_),
    .B2(net405),
    .X(_09398_));
 sky130_fd_sc_hd__nor2_1 _17412_ (.A(_09353_),
    .B(net396),
    .Y(_09399_));
 sky130_fd_sc_hd__a2bb2o_1 _17413_ (.A1_N(net400),
    .A2_N(_09360_),
    .B1(_09399_),
    .B2(net352),
    .X(_09400_));
 sky130_fd_sc_hd__inv_2 _17414_ (.A(net407),
    .Y(_09401_));
 sky130_fd_sc_hd__o21a_1 _17415_ (.A1(net410),
    .A2(_09401_),
    .B1(net352),
    .X(_09402_));
 sky130_fd_sc_hd__nor2_1 _17416_ (.A(_09360_),
    .B(_09402_),
    .Y(_09403_));
 sky130_fd_sc_hd__a221o_1 _17417_ (.A1(net353),
    .A2(_09398_),
    .B1(_09400_),
    .B2(_09401_),
    .C1(_09403_),
    .X(_09404_));
 sky130_fd_sc_hd__mux2_1 _17418_ (.A0(_09393_),
    .A1(_09350_),
    .S(_09404_),
    .X(_09405_));
 sky130_fd_sc_hd__or2_1 _17419_ (.A(_09391_),
    .B(_09405_),
    .X(_09406_));
 sky130_fd_sc_hd__and2_2 _17420_ (.A(net417),
    .B(net337),
    .X(_09407_));
 sky130_fd_sc_hd__nand2_1 _17421_ (.A(net419),
    .B(net333),
    .Y(_09408_));
 sky130_fd_sc_hd__nand2_1 _17422_ (.A(net330),
    .B(net422),
    .Y(_09409_));
 sky130_fd_sc_hd__xor2_2 _17423_ (.A(_09408_),
    .B(_09409_),
    .X(_09410_));
 sky130_fd_sc_hd__xnor2_4 _17424_ (.A(_09407_),
    .B(_09410_),
    .Y(_09411_));
 sky130_fd_sc_hd__nand2_2 _17425_ (.A(net329),
    .B(net425),
    .Y(_09412_));
 sky130_fd_sc_hd__xor2_4 _17426_ (.A(_09411_),
    .B(_09412_),
    .X(_09413_));
 sky130_fd_sc_hd__and2_2 _17427_ (.A(net413),
    .B(net340),
    .X(_09414_));
 sky130_fd_sc_hd__nand2_1 _17428_ (.A(net407),
    .B(net343),
    .Y(_09415_));
 sky130_fd_sc_hd__nand2_1 _17429_ (.A(net403),
    .B(net347),
    .Y(_09416_));
 sky130_fd_sc_hd__xor2_2 _17430_ (.A(_09415_),
    .B(_09416_),
    .X(_09417_));
 sky130_fd_sc_hd__xnor2_4 _17431_ (.A(_09414_),
    .B(_09417_),
    .Y(_09418_));
 sky130_fd_sc_hd__nand4_1 _17432_ (.A(net413),
    .B(net407),
    .C(net343),
    .D(net347),
    .Y(_09419_));
 sky130_fd_sc_hd__a22o_1 _17433_ (.A1(net413),
    .A2(net343),
    .B1(net347),
    .B2(net407),
    .X(_09420_));
 sky130_fd_sc_hd__a21bo_2 _17434_ (.A1(_09369_),
    .A2(_09419_),
    .B1_N(_09420_),
    .X(_09421_));
 sky130_fd_sc_hd__nand4_1 _17435_ (.A(net330),
    .B(net333),
    .C(net422),
    .D(net425),
    .Y(_09422_));
 sky130_fd_sc_hd__a22oi_1 _17436_ (.A1(net333),
    .A2(net422),
    .B1(net427),
    .B2(net330),
    .Y(_09423_));
 sky130_fd_sc_hd__a21oi_2 _17437_ (.A1(_09380_),
    .A2(_09422_),
    .B1(_09423_),
    .Y(_09424_));
 sky130_fd_sc_hd__xnor2_1 _17438_ (.A(_09421_),
    .B(_09424_),
    .Y(_09425_));
 sky130_fd_sc_hd__xnor2_2 _17439_ (.A(_09418_),
    .B(_09425_),
    .Y(_09426_));
 sky130_fd_sc_hd__xnor2_4 _17440_ (.A(_09413_),
    .B(_09426_),
    .Y(_09427_));
 sky130_fd_sc_hd__nand2_1 _17441_ (.A(net392),
    .B(net357),
    .Y(_09428_));
 sky130_fd_sc_hd__nor2_1 _17442_ (.A(_09351_),
    .B(net392),
    .Y(_09429_));
 sky130_fd_sc_hd__a2bb2o_1 _17443_ (.A1_N(net395),
    .A2_N(_09428_),
    .B1(_09429_),
    .B2(net352),
    .X(_09430_));
 sky130_fd_sc_hd__nand2_2 _17444_ (.A(net407),
    .B(net357),
    .Y(_09431_));
 sky130_fd_sc_hd__or2_1 _17445_ (.A(net395),
    .B(net392),
    .X(_09432_));
 sky130_fd_sc_hd__nand2_1 _17446_ (.A(net396),
    .B(net391),
    .Y(_09433_));
 sky130_fd_sc_hd__o21ai_1 _17447_ (.A1(_09431_),
    .A2(_09432_),
    .B1(_09433_),
    .Y(_09434_));
 sky130_fd_sc_hd__a22o_1 _17448_ (.A1(net398),
    .A2(_09395_),
    .B1(_09434_),
    .B2(net400),
    .X(_09435_));
 sky130_fd_sc_hd__o21ba_1 _17449_ (.A1(_09356_),
    .A2(_09354_),
    .B1_N(_09428_),
    .X(_09436_));
 sky130_fd_sc_hd__a221o_2 _17450_ (.A1(_09353_),
    .A2(_09430_),
    .B1(_09435_),
    .B2(net355),
    .C1(_09436_),
    .X(_09437_));
 sky130_fd_sc_hd__nand2_1 _17451_ (.A(_09379_),
    .B(_09384_),
    .Y(_09438_));
 sky130_fd_sc_hd__or2b_1 _17452_ (.A(_09373_),
    .B_N(_09375_),
    .X(_09439_));
 sky130_fd_sc_hd__nor2_1 _17453_ (.A(_09379_),
    .B(_09384_),
    .Y(_09440_));
 sky130_fd_sc_hd__inv_2 _17454_ (.A(_09440_),
    .Y(_09441_));
 sky130_fd_sc_hd__a21oi_1 _17455_ (.A1(_09379_),
    .A2(_09384_),
    .B1(_09375_),
    .Y(_09442_));
 sky130_fd_sc_hd__o21ai_1 _17456_ (.A1(_09442_),
    .A2(_09440_),
    .B1(_09373_),
    .Y(_09443_));
 sky130_fd_sc_hd__o221a_1 _17457_ (.A1(_09438_),
    .A2(_09439_),
    .B1(_09441_),
    .B2(_09375_),
    .C1(_09443_),
    .X(_09444_));
 sky130_fd_sc_hd__xor2_1 _17458_ (.A(_09437_),
    .B(_09444_),
    .X(_09445_));
 sky130_fd_sc_hd__xnor2_2 _17459_ (.A(_09427_),
    .B(_09445_),
    .Y(_09446_));
 sky130_fd_sc_hd__xnor2_1 _17460_ (.A(_09406_),
    .B(_09446_),
    .Y(_09447_));
 sky130_fd_sc_hd__nand2_1 _17461_ (.A(_09368_),
    .B(_09447_),
    .Y(_09448_));
 sky130_fd_sc_hd__or3b_1 _17462_ (.A(_09368_),
    .B(_09446_),
    .C_N(_09406_),
    .X(_09449_));
 sky130_fd_sc_hd__o21ai_1 _17463_ (.A1(_09376_),
    .A2(_09379_),
    .B1(_09384_),
    .Y(_09450_));
 sky130_fd_sc_hd__o21a_1 _17464_ (.A1(_09427_),
    .A2(_09440_),
    .B1(_09439_),
    .X(_09451_));
 sky130_fd_sc_hd__a211oi_1 _17465_ (.A1(_09373_),
    .A2(_09442_),
    .B1(_09451_),
    .C1(_09437_),
    .Y(_09452_));
 sky130_fd_sc_hd__nor2_1 _17466_ (.A(_09427_),
    .B(_09438_),
    .Y(_09453_));
 sky130_fd_sc_hd__nand2_1 _17467_ (.A(_09376_),
    .B(_09379_),
    .Y(_09454_));
 sky130_fd_sc_hd__o211a_1 _17468_ (.A1(_09439_),
    .A2(_09453_),
    .B1(_09454_),
    .C1(_09437_),
    .X(_09455_));
 sky130_fd_sc_hd__o2bb2a_1 _17469_ (.A1_N(_09427_),
    .A2_N(_09450_),
    .B1(_09452_),
    .B2(_09455_),
    .X(_09456_));
 sky130_fd_sc_hd__a21bo_1 _17470_ (.A1(_09375_),
    .A2(_09379_),
    .B1_N(_09373_),
    .X(_09457_));
 sky130_fd_sc_hd__o21ai_1 _17471_ (.A1(_09375_),
    .A2(_09379_),
    .B1(_09457_),
    .Y(_09458_));
 sky130_fd_sc_hd__nand2_1 _17472_ (.A(_09351_),
    .B(net390),
    .Y(_09459_));
 sky130_fd_sc_hd__nand2_1 _17473_ (.A(net407),
    .B(net400),
    .Y(_09460_));
 sky130_fd_sc_hd__or3_1 _17474_ (.A(_09363_),
    .B(_09459_),
    .C(_09460_),
    .X(_09461_));
 sky130_fd_sc_hd__o21ai_1 _17475_ (.A1(net400),
    .A2(net394),
    .B1(net359),
    .Y(_09462_));
 sky130_fd_sc_hd__o21ai_1 _17476_ (.A1(net395),
    .A2(_09431_),
    .B1(_09433_),
    .Y(_09463_));
 sky130_fd_sc_hd__a22o_1 _17477_ (.A1(net398),
    .A2(_09462_),
    .B1(_09463_),
    .B2(net400),
    .X(_09464_));
 sky130_fd_sc_hd__nand2_1 _17478_ (.A(net354),
    .B(_09464_),
    .Y(_09465_));
 sky130_fd_sc_hd__or2_1 _17479_ (.A(_09357_),
    .B(_09428_),
    .X(_09466_));
 sky130_fd_sc_hd__a22o_1 _17480_ (.A1(_09458_),
    .A2(_09461_),
    .B1(_09465_),
    .B2(_09466_),
    .X(_09467_));
 sky130_fd_sc_hd__and2_1 _17481_ (.A(net408),
    .B(net340),
    .X(_09468_));
 sky130_fd_sc_hd__nand2_1 _17482_ (.A(net403),
    .B(net343),
    .Y(_09469_));
 sky130_fd_sc_hd__nand2_1 _17483_ (.A(net398),
    .B(net350),
    .Y(_09470_));
 sky130_fd_sc_hd__xor2_1 _17484_ (.A(_09469_),
    .B(_09470_),
    .X(_09471_));
 sky130_fd_sc_hd__xnor2_2 _17485_ (.A(_09468_),
    .B(_09471_),
    .Y(_09472_));
 sky130_fd_sc_hd__and4_1 _17486_ (.A(net408),
    .B(net403),
    .C(net343),
    .D(net347),
    .X(_09473_));
 sky130_fd_sc_hd__a22o_1 _17487_ (.A1(net408),
    .A2(net343),
    .B1(net347),
    .B2(net403),
    .X(_09474_));
 sky130_fd_sc_hd__o21a_1 _17488_ (.A1(_09414_),
    .A2(_09473_),
    .B1(_09474_),
    .X(_09475_));
 sky130_fd_sc_hd__and4_1 _17489_ (.A(net419),
    .B(net330),
    .C(net333),
    .D(net422),
    .X(_09476_));
 sky130_fd_sc_hd__a22o_1 _17490_ (.A1(net419),
    .A2(net333),
    .B1(net422),
    .B2(net330),
    .X(_09477_));
 sky130_fd_sc_hd__o21a_1 _17491_ (.A1(_09407_),
    .A2(_09476_),
    .B1(_09477_),
    .X(_09478_));
 sky130_fd_sc_hd__xor2_1 _17492_ (.A(_09475_),
    .B(_09478_),
    .X(_09479_));
 sky130_fd_sc_hd__xnor2_2 _17493_ (.A(_09472_),
    .B(_09479_),
    .Y(_09480_));
 sky130_fd_sc_hd__nor2_1 _17494_ (.A(_09411_),
    .B(_09412_),
    .Y(_09481_));
 sky130_fd_sc_hd__nand2_1 _17495_ (.A(net413),
    .B(net337),
    .Y(_09482_));
 sky130_fd_sc_hd__and2_1 _17496_ (.A(net417),
    .B(net333),
    .X(_09483_));
 sky130_fd_sc_hd__nand2_1 _17497_ (.A(net419),
    .B(net330),
    .Y(_09484_));
 sky130_fd_sc_hd__xor2_1 _17498_ (.A(_09483_),
    .B(_09484_),
    .X(_09485_));
 sky130_fd_sc_hd__xnor2_1 _17499_ (.A(_09482_),
    .B(_09485_),
    .Y(_09486_));
 sky130_fd_sc_hd__nand2_1 _17500_ (.A(net325),
    .B(net427),
    .Y(_09487_));
 sky130_fd_sc_hd__nand2_1 _17501_ (.A(net329),
    .B(net422),
    .Y(_09488_));
 sky130_fd_sc_hd__xor2_1 _17502_ (.A(_09487_),
    .B(_09488_),
    .X(_09489_));
 sky130_fd_sc_hd__xnor2_1 _17503_ (.A(_09486_),
    .B(_09489_),
    .Y(_09490_));
 sky130_fd_sc_hd__xnor2_1 _17504_ (.A(_09481_),
    .B(_09490_),
    .Y(_09491_));
 sky130_fd_sc_hd__xor2_1 _17505_ (.A(_09480_),
    .B(_09491_),
    .X(_09492_));
 sky130_fd_sc_hd__inv_2 _17506_ (.A(net390),
    .Y(_09493_));
 sky130_fd_sc_hd__nor2_1 _17507_ (.A(_09493_),
    .B(net385),
    .Y(_09494_));
 sky130_fd_sc_hd__nand2_1 _17508_ (.A(net388),
    .B(net357),
    .Y(_09495_));
 sky130_fd_sc_hd__o2bb2a_1 _17509_ (.A1_N(net353),
    .A2_N(_09494_),
    .B1(_09495_),
    .B2(net390),
    .X(_09496_));
 sky130_fd_sc_hd__a21oi_1 _17510_ (.A1(_09352_),
    .A2(net395),
    .B1(_09355_),
    .Y(_09497_));
 sky130_fd_sc_hd__nand2_1 _17511_ (.A(net391),
    .B(net385),
    .Y(_09498_));
 sky130_fd_sc_hd__or4bb_1 _17512_ (.A(net390),
    .B(net386),
    .C_N(net358),
    .D_N(net401),
    .X(_09499_));
 sky130_fd_sc_hd__nand2_1 _17513_ (.A(_09498_),
    .B(_09499_),
    .Y(_09500_));
 sky130_fd_sc_hd__a22o_1 _17514_ (.A1(net391),
    .A2(_09395_),
    .B1(_09500_),
    .B2(net395),
    .X(_09501_));
 sky130_fd_sc_hd__nand2_1 _17515_ (.A(net352),
    .B(_09501_),
    .Y(_09502_));
 sky130_fd_sc_hd__o221a_2 _17516_ (.A1(net395),
    .A2(_09496_),
    .B1(_09497_),
    .B2(_09495_),
    .C1(_09502_),
    .X(_09503_));
 sky130_fd_sc_hd__xnor2_1 _17517_ (.A(_09492_),
    .B(_09503_),
    .Y(_09504_));
 sky130_fd_sc_hd__nand2_1 _17518_ (.A(_09418_),
    .B(_09421_),
    .Y(_09505_));
 sky130_fd_sc_hd__inv_2 _17519_ (.A(_09424_),
    .Y(_09506_));
 sky130_fd_sc_hd__o21ai_1 _17520_ (.A1(_09418_),
    .A2(_09421_),
    .B1(_09506_),
    .Y(_09507_));
 sky130_fd_sc_hd__a21o_1 _17521_ (.A1(_09505_),
    .A2(_09507_),
    .B1(_09413_),
    .X(_09508_));
 sky130_fd_sc_hd__or2_1 _17522_ (.A(_09424_),
    .B(_09505_),
    .X(_09509_));
 sky130_fd_sc_hd__nand2_1 _17523_ (.A(_09413_),
    .B(_09424_),
    .Y(_09510_));
 sky130_fd_sc_hd__or3_1 _17524_ (.A(_09418_),
    .B(_09421_),
    .C(_09510_),
    .X(_09511_));
 sky130_fd_sc_hd__and3_1 _17525_ (.A(_09508_),
    .B(_09509_),
    .C(_09511_),
    .X(_09512_));
 sky130_fd_sc_hd__xnor2_2 _17526_ (.A(_09504_),
    .B(_09512_),
    .Y(_09513_));
 sky130_fd_sc_hd__xnor2_1 _17527_ (.A(_09467_),
    .B(_09513_),
    .Y(_09514_));
 sky130_fd_sc_hd__xnor2_1 _17528_ (.A(_09456_),
    .B(_09514_),
    .Y(_09515_));
 sky130_fd_sc_hd__a21o_1 _17529_ (.A1(_09448_),
    .A2(_09449_),
    .B1(_09515_),
    .X(_09516_));
 sky130_fd_sc_hd__or4b_1 _17530_ (.A(_09391_),
    .B(_09368_),
    .C(_09405_),
    .D_N(_09446_),
    .X(_09517_));
 sky130_fd_sc_hd__nor2_4 _17531_ (.A(_09355_),
    .B(_09395_),
    .Y(_09518_));
 sky130_fd_sc_hd__and3_1 _17532_ (.A(net415),
    .B(net412),
    .C(_09354_),
    .X(_09519_));
 sky130_fd_sc_hd__xnor2_1 _17533_ (.A(_09340_),
    .B(_09341_),
    .Y(_09520_));
 sky130_fd_sc_hd__xnor2_2 _17534_ (.A(_09342_),
    .B(_09520_),
    .Y(_09521_));
 sky130_fd_sc_hd__nand2_1 _17535_ (.A(net422),
    .B(net343),
    .Y(_09522_));
 sky130_fd_sc_hd__nand2_1 _17536_ (.A(net340),
    .B(net425),
    .Y(_09523_));
 sky130_fd_sc_hd__and3_1 _17537_ (.A(net423),
    .B(net343),
    .C(net425),
    .X(_09524_));
 sky130_fd_sc_hd__and2_1 _17538_ (.A(net418),
    .B(net349),
    .X(_09525_));
 sky130_fd_sc_hd__a21oi_1 _17539_ (.A1(net340),
    .A2(_09524_),
    .B1(_09525_),
    .Y(_09526_));
 sky130_fd_sc_hd__a21o_1 _17540_ (.A1(_09522_),
    .A2(_09523_),
    .B1(_09526_),
    .X(_09527_));
 sky130_fd_sc_hd__nor2_1 _17541_ (.A(_09521_),
    .B(_09527_),
    .Y(_09528_));
 sky130_fd_sc_hd__nand2_1 _17542_ (.A(net407),
    .B(net354),
    .Y(_09529_));
 sky130_fd_sc_hd__o21ai_1 _17543_ (.A1(net412),
    .A2(net403),
    .B1(net358),
    .Y(_09530_));
 sky130_fd_sc_hd__nand2_1 _17544_ (.A(net417),
    .B(net358),
    .Y(_09531_));
 sky130_fd_sc_hd__o21ai_1 _17545_ (.A1(net407),
    .A2(_09531_),
    .B1(_09460_),
    .Y(_09532_));
 sky130_fd_sc_hd__a22o_1 _17546_ (.A1(net407),
    .A2(_09530_),
    .B1(_09532_),
    .B2(net412),
    .X(_09533_));
 sky130_fd_sc_hd__a32o_1 _17547_ (.A1(net403),
    .A2(net358),
    .A3(_09529_),
    .B1(_09533_),
    .B2(net354),
    .X(_09534_));
 sky130_fd_sc_hd__a22o_1 _17548_ (.A1(_09518_),
    .A2(_09519_),
    .B1(_09528_),
    .B2(_09534_),
    .X(_09535_));
 sky130_fd_sc_hd__a21boi_1 _17549_ (.A1(_09518_),
    .A2(_09519_),
    .B1_N(_09534_),
    .Y(_09536_));
 sky130_fd_sc_hd__xor2_2 _17550_ (.A(_09528_),
    .B(_09536_),
    .X(_09537_));
 sky130_fd_sc_hd__xor2_1 _17551_ (.A(_09344_),
    .B(_09389_),
    .X(_09538_));
 sky130_fd_sc_hd__xnor2_2 _17552_ (.A(_09349_),
    .B(_09538_),
    .Y(_09539_));
 sky130_fd_sc_hd__nand2_1 _17553_ (.A(net337),
    .B(net425),
    .Y(_09540_));
 sky130_fd_sc_hd__xnor2_2 _17554_ (.A(_09521_),
    .B(_09527_),
    .Y(_09541_));
 sky130_fd_sc_hd__nor2_1 _17555_ (.A(_09540_),
    .B(_09541_),
    .Y(_09542_));
 sky130_fd_sc_hd__a21o_1 _17556_ (.A1(_09537_),
    .A2(_09539_),
    .B1(_09542_),
    .X(_09543_));
 sky130_fd_sc_hd__o21a_1 _17557_ (.A1(_09537_),
    .A2(_09539_),
    .B1(_09543_),
    .X(_09544_));
 sky130_fd_sc_hd__xor2_1 _17558_ (.A(_09404_),
    .B(_09392_),
    .X(_09545_));
 sky130_fd_sc_hd__xnor2_1 _17559_ (.A(_09386_),
    .B(_09545_),
    .Y(_09546_));
 sky130_fd_sc_hd__or2_1 _17560_ (.A(_09544_),
    .B(_09546_),
    .X(_09547_));
 sky130_fd_sc_hd__a21o_1 _17561_ (.A1(_09544_),
    .A2(_09546_),
    .B1(_09535_),
    .X(_09548_));
 sky130_fd_sc_hd__and2_1 _17562_ (.A(net418),
    .B(net340),
    .X(_09549_));
 sky130_fd_sc_hd__nor2_1 _17563_ (.A(net418),
    .B(net340),
    .Y(_09550_));
 sky130_fd_sc_hd__o211ai_2 _17564_ (.A1(_09549_),
    .A2(_09550_),
    .B1(net347),
    .C1(_09524_),
    .Y(_09551_));
 sky130_fd_sc_hd__nand2_1 _17565_ (.A(net418),
    .B(net354),
    .Y(_09552_));
 sky130_fd_sc_hd__or3_1 _17566_ (.A(net412),
    .B(_09531_),
    .C(_09552_),
    .X(_09553_));
 sky130_fd_sc_hd__nand2_1 _17567_ (.A(_09551_),
    .B(_09553_),
    .Y(_09554_));
 sky130_fd_sc_hd__xor2_2 _17568_ (.A(_09540_),
    .B(_09541_),
    .X(_09555_));
 sky130_fd_sc_hd__nor2_1 _17569_ (.A(_09551_),
    .B(_09553_),
    .Y(_09556_));
 sky130_fd_sc_hd__or2_1 _17570_ (.A(_09555_),
    .B(_09556_),
    .X(_09557_));
 sky130_fd_sc_hd__or2_1 _17571_ (.A(_09555_),
    .B(_09554_),
    .X(_09558_));
 sky130_fd_sc_hd__or2b_1 _17572_ (.A(net415),
    .B_N(net410),
    .X(_09559_));
 sky130_fd_sc_hd__a2bb2o_1 _17573_ (.A1_N(_09529_),
    .A2_N(_09559_),
    .B1(net415),
    .B2(_09401_),
    .X(_09560_));
 sky130_fd_sc_hd__nand2_1 _17574_ (.A(net410),
    .B(net352),
    .Y(_09561_));
 sky130_fd_sc_hd__a22oi_4 _17575_ (.A1(net359),
    .A2(_09560_),
    .B1(_09431_),
    .B2(_09561_),
    .Y(_09562_));
 sky130_fd_sc_hd__a22o_1 _17576_ (.A1(_09554_),
    .A2(_09557_),
    .B1(_09558_),
    .B2(_09562_),
    .X(_09563_));
 sky130_fd_sc_hd__xnor2_1 _17577_ (.A(_09539_),
    .B(_09542_),
    .Y(_09564_));
 sky130_fd_sc_hd__xnor2_1 _17578_ (.A(_09537_),
    .B(_09564_),
    .Y(_09565_));
 sky130_fd_sc_hd__a31o_1 _17579_ (.A1(_09555_),
    .A2(_09562_),
    .A3(_09556_),
    .B1(_09565_),
    .X(_09566_));
 sky130_fd_sc_hd__inv_2 _17580_ (.A(net420),
    .Y(_09567_));
 sky130_fd_sc_hd__and4b_1 _17581_ (.A_N(net415),
    .B(net418),
    .C(net423),
    .D(net358),
    .X(_09568_));
 sky130_fd_sc_hd__a21oi_1 _17582_ (.A1(net415),
    .A2(_09567_),
    .B1(_09568_),
    .Y(_09569_));
 sky130_fd_sc_hd__a21o_1 _17583_ (.A1(net412),
    .A2(net418),
    .B1(_09395_),
    .X(_09570_));
 sky130_fd_sc_hd__a2bb2o_1 _17584_ (.A1_N(net412),
    .A2_N(_09569_),
    .B1(_09570_),
    .B2(net415),
    .X(_09571_));
 sky130_fd_sc_hd__a21oi_1 _17585_ (.A1(net418),
    .A2(net423),
    .B1(net415),
    .Y(_09572_));
 sky130_fd_sc_hd__o211a_1 _17586_ (.A1(_09356_),
    .A2(_09572_),
    .B1(net360),
    .C1(net410),
    .X(_09573_));
 sky130_fd_sc_hd__a21oi_1 _17587_ (.A1(net354),
    .A2(_09571_),
    .B1(_09573_),
    .Y(_09574_));
 sky130_fd_sc_hd__o22ai_1 _17588_ (.A1(net342),
    .A2(net349),
    .B1(net425),
    .B2(_09525_),
    .Y(_09575_));
 sky130_fd_sc_hd__o21ai_1 _17589_ (.A1(net425),
    .A2(_09522_),
    .B1(_09523_),
    .Y(_09576_));
 sky130_fd_sc_hd__a22o_1 _17590_ (.A1(net425),
    .A2(_09550_),
    .B1(_09576_),
    .B2(net418),
    .X(_09577_));
 sky130_fd_sc_hd__and3b_1 _17591_ (.A_N(net347),
    .B(_09524_),
    .C(net340),
    .X(_09578_));
 sky130_fd_sc_hd__a221o_1 _17592_ (.A1(_09522_),
    .A2(_09575_),
    .B1(_09577_),
    .B2(net347),
    .C1(_09578_),
    .X(_09579_));
 sky130_fd_sc_hd__a21o_1 _17593_ (.A1(net422),
    .A2(net358),
    .B1(_09552_),
    .X(_09580_));
 sky130_fd_sc_hd__nand2_1 _17594_ (.A(_09531_),
    .B(_09580_),
    .Y(_09581_));
 sky130_fd_sc_hd__o31a_1 _17595_ (.A1(net423),
    .A2(_09531_),
    .A3(_09552_),
    .B1(_09581_),
    .X(_09582_));
 sky130_fd_sc_hd__a21o_1 _17596_ (.A1(_09567_),
    .A2(net359),
    .B1(net349),
    .X(_09583_));
 sky130_fd_sc_hd__a32o_1 _17597_ (.A1(net423),
    .A2(net354),
    .A3(_09583_),
    .B1(_09525_),
    .B2(net359),
    .X(_09584_));
 sky130_fd_sc_hd__nand2_1 _17598_ (.A(net422),
    .B(net349),
    .Y(_09585_));
 sky130_fd_sc_hd__and3_1 _17599_ (.A(net345),
    .B(net426),
    .C(_09585_),
    .X(_09586_));
 sky130_fd_sc_hd__a21oi_1 _17600_ (.A1(net345),
    .A2(net426),
    .B1(_09585_),
    .Y(_09587_));
 sky130_fd_sc_hd__a311o_1 _17601_ (.A1(net425),
    .A2(_09582_),
    .A3(_09584_),
    .B1(_09586_),
    .C1(_09587_),
    .X(_09588_));
 sky130_fd_sc_hd__a21o_1 _17602_ (.A1(net425),
    .A2(_09584_),
    .B1(_09582_),
    .X(_09589_));
 sky130_fd_sc_hd__nor2_1 _17603_ (.A(_09574_),
    .B(_09579_),
    .Y(_09590_));
 sky130_fd_sc_hd__a21oi_1 _17604_ (.A1(_09588_),
    .A2(_09589_),
    .B1(_09590_),
    .Y(_09591_));
 sky130_fd_sc_hd__a21oi_1 _17605_ (.A1(_09574_),
    .A2(_09579_),
    .B1(_09591_),
    .Y(_09592_));
 sky130_fd_sc_hd__inv_2 _17606_ (.A(net423),
    .Y(_09593_));
 sky130_fd_sc_hd__or4_1 _17607_ (.A(_09567_),
    .B(_09593_),
    .C(_09364_),
    .D(_09559_),
    .X(_09594_));
 sky130_fd_sc_hd__xnor2_1 _17608_ (.A(_09551_),
    .B(_09553_),
    .Y(_09595_));
 sky130_fd_sc_hd__xnor2_1 _17609_ (.A(_09562_),
    .B(_09595_),
    .Y(_09596_));
 sky130_fd_sc_hd__xnor2_1 _17610_ (.A(_09555_),
    .B(_09596_),
    .Y(_09597_));
 sky130_fd_sc_hd__nor2_1 _17611_ (.A(_09594_),
    .B(_09597_),
    .Y(_09598_));
 sky130_fd_sc_hd__nand2_1 _17612_ (.A(_09594_),
    .B(_09597_),
    .Y(_09599_));
 sky130_fd_sc_hd__o221a_1 _17613_ (.A1(_09565_),
    .A2(_09563_),
    .B1(_09592_),
    .B2(_09598_),
    .C1(_09599_),
    .X(_09600_));
 sky130_fd_sc_hd__a21o_1 _17614_ (.A1(_09563_),
    .A2(_09566_),
    .B1(_09600_),
    .X(_09601_));
 sky130_fd_sc_hd__a21o_1 _17615_ (.A1(_09547_),
    .A2(_09548_),
    .B1(_09601_),
    .X(_09602_));
 sky130_fd_sc_hd__o21ai_1 _17616_ (.A1(_09535_),
    .A2(_09547_),
    .B1(_09602_),
    .Y(_09603_));
 sky130_fd_sc_hd__nand2_1 _17617_ (.A(net408),
    .B(net337),
    .Y(_09604_));
 sky130_fd_sc_hd__nand2_1 _17618_ (.A(net413),
    .B(net335),
    .Y(_09605_));
 sky130_fd_sc_hd__nand2_1 _17619_ (.A(net417),
    .B(net331),
    .Y(_09606_));
 sky130_fd_sc_hd__xor2_1 _17620_ (.A(_09605_),
    .B(_09606_),
    .X(_09607_));
 sky130_fd_sc_hd__xnor2_2 _17621_ (.A(_09604_),
    .B(_09607_),
    .Y(_09608_));
 sky130_fd_sc_hd__nand2_2 _17622_ (.A(net325),
    .B(net424),
    .Y(_09609_));
 sky130_fd_sc_hd__and2_1 _17623_ (.A(net1023),
    .B(net427),
    .X(_09610_));
 sky130_fd_sc_hd__o22a_1 _17624_ (.A1(net420),
    .A2(net426),
    .B1(_09610_),
    .B2(net1022),
    .X(_09611_));
 sky130_fd_sc_hd__nand2_2 _17625_ (.A(net1022),
    .B(net420),
    .Y(_09612_));
 sky130_fd_sc_hd__o21a_1 _17626_ (.A1(net1022),
    .A2(_09609_),
    .B1(_09612_),
    .X(_09613_));
 sky130_fd_sc_hd__nor2_1 _17627_ (.A(net1023),
    .B(_09612_),
    .Y(_09614_));
 sky130_fd_sc_hd__a21oi_1 _17628_ (.A1(net1023),
    .A2(_09613_),
    .B1(_09614_),
    .Y(_09615_));
 sky130_fd_sc_hd__inv_2 _17629_ (.A(net427),
    .Y(_09616_));
 sky130_fd_sc_hd__or3b_1 _17630_ (.A(net426),
    .B(_09612_),
    .C_N(_09609_),
    .X(_09617_));
 sky130_fd_sc_hd__o221a_1 _17631_ (.A1(_09609_),
    .A2(_09611_),
    .B1(_09615_),
    .B2(_09616_),
    .C1(_09617_),
    .X(_09618_));
 sky130_fd_sc_hd__xor2_2 _17632_ (.A(_09608_),
    .B(_09618_),
    .X(_09619_));
 sky130_fd_sc_hd__nand2_1 _17633_ (.A(net392),
    .B(net349),
    .Y(_09620_));
 sky130_fd_sc_hd__nand2_1 _17634_ (.A(net403),
    .B(net342),
    .Y(_09621_));
 sky130_fd_sc_hd__nand2_1 _17635_ (.A(net398),
    .B(net345),
    .Y(_09622_));
 sky130_fd_sc_hd__xnor2_1 _17636_ (.A(_09621_),
    .B(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__xnor2_2 _17637_ (.A(_09620_),
    .B(_09623_),
    .Y(_09624_));
 sky130_fd_sc_hd__and4_1 _17638_ (.A(net403),
    .B(net398),
    .C(net344),
    .D(net348),
    .X(_09625_));
 sky130_fd_sc_hd__a22o_1 _17639_ (.A1(net403),
    .A2(net344),
    .B1(net348),
    .B2(net398),
    .X(_09626_));
 sky130_fd_sc_hd__o21a_1 _17640_ (.A1(_09468_),
    .A2(_09625_),
    .B1(_09626_),
    .X(_09627_));
 sky130_fd_sc_hd__and4_1 _17641_ (.A(net412),
    .B(net419),
    .C(net330),
    .D(net337),
    .X(_09628_));
 sky130_fd_sc_hd__a22o_1 _17642_ (.A1(net419),
    .A2(net330),
    .B1(net337),
    .B2(net412),
    .X(_09629_));
 sky130_fd_sc_hd__o21a_1 _17643_ (.A1(_09483_),
    .A2(_09628_),
    .B1(_09629_),
    .X(_09630_));
 sky130_fd_sc_hd__xnor2_1 _17644_ (.A(_09627_),
    .B(_09630_),
    .Y(_09631_));
 sky130_fd_sc_hd__xnor2_2 _17645_ (.A(_09624_),
    .B(_09631_),
    .Y(_09632_));
 sky130_fd_sc_hd__or2b_1 _17646_ (.A(_09486_),
    .B_N(_09489_),
    .X(_09633_));
 sky130_fd_sc_hd__o21a_1 _17647_ (.A1(_09619_),
    .A2(_09632_),
    .B1(_09633_),
    .X(_09634_));
 sky130_fd_sc_hd__a21o_1 _17648_ (.A1(_09619_),
    .A2(_09632_),
    .B1(_09634_),
    .X(_09635_));
 sky130_fd_sc_hd__nand2_2 _17649_ (.A(net426),
    .B(net319),
    .Y(_09636_));
 sky130_fd_sc_hd__nand2_1 _17650_ (.A(net382),
    .B(net355),
    .Y(_09637_));
 sky130_fd_sc_hd__o21a_1 _17651_ (.A1(net388),
    .A2(net378),
    .B1(net359),
    .X(_09638_));
 sky130_fd_sc_hd__mux2_1 _17652_ (.A0(net388),
    .A1(net359),
    .S(_09637_),
    .X(_09639_));
 sky130_fd_sc_hd__a2bb2o_1 _17653_ (.A1_N(_09637_),
    .A2_N(_09638_),
    .B1(_09639_),
    .B2(net378),
    .X(_09640_));
 sky130_fd_sc_hd__xnor2_1 _17654_ (.A(_09636_),
    .B(_09640_),
    .Y(_09641_));
 sky130_fd_sc_hd__nand2_1 _17655_ (.A(_09627_),
    .B(_09630_),
    .Y(_09642_));
 sky130_fd_sc_hd__nor2_1 _17656_ (.A(_09627_),
    .B(_09630_),
    .Y(_09643_));
 sky130_fd_sc_hd__a21o_1 _17657_ (.A1(_09642_),
    .A2(_09624_),
    .B1(_09643_),
    .X(_09644_));
 sky130_fd_sc_hd__or3_2 _17658_ (.A(net382),
    .B(_09362_),
    .C(_09498_),
    .X(_09645_));
 sky130_fd_sc_hd__xor2_1 _17659_ (.A(_09644_),
    .B(_09645_),
    .X(_09646_));
 sky130_fd_sc_hd__xnor2_1 _17660_ (.A(_09641_),
    .B(_09646_),
    .Y(_09647_));
 sky130_fd_sc_hd__nand2_1 _17661_ (.A(net322),
    .B(net424),
    .Y(_09648_));
 sky130_fd_sc_hd__nand2_1 _17662_ (.A(\top0.pid_d.mult0.a[3] ),
    .B(net329),
    .Y(_09649_));
 sky130_fd_sc_hd__nand2_1 _17663_ (.A(net326),
    .B(net420),
    .Y(_09650_));
 sky130_fd_sc_hd__xnor2_1 _17664_ (.A(_09649_),
    .B(_09650_),
    .Y(_09651_));
 sky130_fd_sc_hd__xnor2_2 _17665_ (.A(_09648_),
    .B(_09651_),
    .Y(_09652_));
 sky130_fd_sc_hd__nor2_1 _17666_ (.A(_09609_),
    .B(_09612_),
    .Y(_09653_));
 sky130_fd_sc_hd__nand2_1 _17667_ (.A(_09609_),
    .B(_09612_),
    .Y(_09654_));
 sky130_fd_sc_hd__o21ai_1 _17668_ (.A1(_09610_),
    .A2(_09653_),
    .B1(_09654_),
    .Y(_09655_));
 sky130_fd_sc_hd__nand2_1 _17669_ (.A(net404),
    .B(net337),
    .Y(_09656_));
 sky130_fd_sc_hd__nand2_1 _17670_ (.A(net409),
    .B(net333),
    .Y(_09657_));
 sky130_fd_sc_hd__nand2_1 _17671_ (.A(net414),
    .B(net330),
    .Y(_09658_));
 sky130_fd_sc_hd__xnor2_1 _17672_ (.A(_09657_),
    .B(_09658_),
    .Y(_09659_));
 sky130_fd_sc_hd__xnor2_2 _17673_ (.A(_09656_),
    .B(_09659_),
    .Y(_09660_));
 sky130_fd_sc_hd__xnor2_1 _17674_ (.A(_09655_),
    .B(_09660_),
    .Y(_09661_));
 sky130_fd_sc_hd__xnor2_2 _17675_ (.A(_09652_),
    .B(_09661_),
    .Y(_09662_));
 sky130_fd_sc_hd__or3_1 _17676_ (.A(net426),
    .B(_09609_),
    .C(_09612_),
    .X(_09663_));
 sky130_fd_sc_hd__mux2_1 _17677_ (.A0(_09654_),
    .A1(_09613_),
    .S(_09610_),
    .X(_09664_));
 sky130_fd_sc_hd__nor2_1 _17678_ (.A(net322),
    .B(net420),
    .Y(_09665_));
 sky130_fd_sc_hd__and2_1 _17679_ (.A(net322),
    .B(net420),
    .X(_09666_));
 sky130_fd_sc_hd__and4_1 _17680_ (.A(net326),
    .B(net329),
    .C(net424),
    .D(net427),
    .X(_09667_));
 sky130_fd_sc_hd__o21a_1 _17681_ (.A1(_09665_),
    .A2(_09666_),
    .B1(_09667_),
    .X(_09668_));
 sky130_fd_sc_hd__a31o_1 _17682_ (.A1(_09608_),
    .A2(_09663_),
    .A3(_09664_),
    .B1(_09668_),
    .X(_09669_));
 sky130_fd_sc_hd__nand2_1 _17683_ (.A(net388),
    .B(net349),
    .Y(_09670_));
 sky130_fd_sc_hd__nand2_1 _17684_ (.A(net399),
    .B(net342),
    .Y(_09671_));
 sky130_fd_sc_hd__nand2_1 _17685_ (.A(net393),
    .B(net345),
    .Y(_09672_));
 sky130_fd_sc_hd__xnor2_1 _17686_ (.A(_09671_),
    .B(_09672_),
    .Y(_09673_));
 sky130_fd_sc_hd__xnor2_1 _17687_ (.A(_09670_),
    .B(_09673_),
    .Y(_09674_));
 sky130_fd_sc_hd__a22o_1 _17688_ (.A1(net413),
    .A2(net333),
    .B1(net339),
    .B2(net408),
    .X(_09675_));
 sky130_fd_sc_hd__and4_1 _17689_ (.A(net413),
    .B(net408),
    .C(net333),
    .D(net339),
    .X(_09676_));
 sky130_fd_sc_hd__a31o_1 _17690_ (.A1(net417),
    .A2(net332),
    .A3(_09675_),
    .B1(_09676_),
    .X(_09677_));
 sky130_fd_sc_hd__nand4_1 _17691_ (.A(net398),
    .B(net392),
    .C(net345),
    .D(net349),
    .Y(_09678_));
 sky130_fd_sc_hd__a22oi_1 _17692_ (.A1(net398),
    .A2(net345),
    .B1(net349),
    .B2(net392),
    .Y(_09679_));
 sky130_fd_sc_hd__a21oi_2 _17693_ (.A1(_09621_),
    .A2(_09678_),
    .B1(_09679_),
    .Y(_09680_));
 sky130_fd_sc_hd__xnor2_1 _17694_ (.A(_09677_),
    .B(_09680_),
    .Y(_09681_));
 sky130_fd_sc_hd__xnor2_1 _17695_ (.A(_09674_),
    .B(_09681_),
    .Y(_09682_));
 sky130_fd_sc_hd__xnor2_1 _17696_ (.A(_09669_),
    .B(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__xnor2_2 _17697_ (.A(_09662_),
    .B(_09683_),
    .Y(_09684_));
 sky130_fd_sc_hd__xnor2_1 _17698_ (.A(_09647_),
    .B(_09684_),
    .Y(_09685_));
 sky130_fd_sc_hd__xnor2_1 _17699_ (.A(_09635_),
    .B(_09685_),
    .Y(_09686_));
 sky130_fd_sc_hd__nand2_1 _17700_ (.A(net381),
    .B(net358),
    .Y(_09687_));
 sky130_fd_sc_hd__inv_2 _17701_ (.A(net387),
    .Y(_09688_));
 sky130_fd_sc_hd__nor2_1 _17702_ (.A(_09688_),
    .B(net381),
    .Y(_09689_));
 sky130_fd_sc_hd__a2bb2o_1 _17703_ (.A1_N(net385),
    .A2_N(_09687_),
    .B1(_09689_),
    .B2(net352),
    .X(_09690_));
 sky130_fd_sc_hd__or2_1 _17704_ (.A(net386),
    .B(net381),
    .X(_09691_));
 sky130_fd_sc_hd__nand2_1 _17705_ (.A(net385),
    .B(net381),
    .Y(_09692_));
 sky130_fd_sc_hd__o21ai_1 _17706_ (.A1(_09360_),
    .A2(_09691_),
    .B1(_09692_),
    .Y(_09693_));
 sky130_fd_sc_hd__a22o_1 _17707_ (.A1(net386),
    .A2(_09394_),
    .B1(_09693_),
    .B2(net391),
    .X(_09694_));
 sky130_fd_sc_hd__a21oi_1 _17708_ (.A1(net352),
    .A2(_09459_),
    .B1(_09687_),
    .Y(_09695_));
 sky130_fd_sc_hd__a221o_2 _17709_ (.A1(_09493_),
    .A2(_09690_),
    .B1(_09694_),
    .B2(net352),
    .C1(_09695_),
    .X(_09696_));
 sky130_fd_sc_hd__a21bo_1 _17710_ (.A1(_09475_),
    .A2(_09478_),
    .B1_N(_09472_),
    .X(_09697_));
 sky130_fd_sc_hd__o21ai_2 _17711_ (.A1(_09475_),
    .A2(_09478_),
    .B1(_09697_),
    .Y(_09698_));
 sky130_fd_sc_hd__xnor2_2 _17712_ (.A(_09696_),
    .B(_09698_),
    .Y(_09699_));
 sky130_fd_sc_hd__xor2_1 _17713_ (.A(_09632_),
    .B(_09633_),
    .X(_09700_));
 sky130_fd_sc_hd__xnor2_2 _17714_ (.A(_09619_),
    .B(_09700_),
    .Y(_09701_));
 sky130_fd_sc_hd__or2_1 _17715_ (.A(_09699_),
    .B(_09701_),
    .X(_09702_));
 sky130_fd_sc_hd__o21a_1 _17716_ (.A1(_09481_),
    .A2(_09480_),
    .B1(_09490_),
    .X(_09703_));
 sky130_fd_sc_hd__a21o_1 _17717_ (.A1(_09481_),
    .A2(_09480_),
    .B1(_09703_),
    .X(_09704_));
 sky130_fd_sc_hd__a21o_1 _17718_ (.A1(_09699_),
    .A2(_09701_),
    .B1(_09704_),
    .X(_09705_));
 sky130_fd_sc_hd__inv_2 _17719_ (.A(net383),
    .Y(_09706_));
 sky130_fd_sc_hd__or4_1 _17720_ (.A(net385),
    .B(_09706_),
    .C(_09362_),
    .D(_09433_),
    .X(_09707_));
 sky130_fd_sc_hd__nand2_1 _17721_ (.A(net385),
    .B(net352),
    .Y(_09708_));
 sky130_fd_sc_hd__o21ai_1 _17722_ (.A1(net391),
    .A2(net381),
    .B1(net357),
    .Y(_09709_));
 sky130_fd_sc_hd__o21ai_1 _17723_ (.A1(net386),
    .A2(_09360_),
    .B1(_09692_),
    .Y(_09710_));
 sky130_fd_sc_hd__a22o_1 _17724_ (.A1(net385),
    .A2(_09709_),
    .B1(_09710_),
    .B2(net391),
    .X(_09711_));
 sky130_fd_sc_hd__a32o_1 _17725_ (.A1(net382),
    .A2(net357),
    .A3(_09708_),
    .B1(_09711_),
    .B2(net352),
    .X(_09712_));
 sky130_fd_sc_hd__a21boi_1 _17726_ (.A1(_09698_),
    .A2(_09707_),
    .B1_N(_09712_),
    .Y(_09713_));
 sky130_fd_sc_hd__and3_1 _17727_ (.A(_09702_),
    .B(_09705_),
    .C(_09713_),
    .X(_09714_));
 sky130_fd_sc_hd__a21oi_1 _17728_ (.A1(_09702_),
    .A2(_09705_),
    .B1(_09713_),
    .Y(_09715_));
 sky130_fd_sc_hd__or3_1 _17729_ (.A(_09686_),
    .B(_09714_),
    .C(_09715_),
    .X(_09716_));
 sky130_fd_sc_hd__o21ai_1 _17730_ (.A1(_09714_),
    .A2(_09715_),
    .B1(_09686_),
    .Y(_09717_));
 sky130_fd_sc_hd__and2_1 _17731_ (.A(_09716_),
    .B(_09717_),
    .X(_09718_));
 sky130_fd_sc_hd__or4_1 _17732_ (.A(_09353_),
    .B(_09351_),
    .C(net392),
    .D(_09363_),
    .X(_09719_));
 sky130_fd_sc_hd__a2bb2o_1 _17733_ (.A1_N(_09459_),
    .A2_N(_09708_),
    .B1(net395),
    .B2(_09688_),
    .X(_09720_));
 sky130_fd_sc_hd__nand2_1 _17734_ (.A(net392),
    .B(net353),
    .Y(_09721_));
 sky130_fd_sc_hd__a22o_1 _17735_ (.A1(net357),
    .A2(_09720_),
    .B1(_09721_),
    .B2(_09495_),
    .X(_09722_));
 sky130_fd_sc_hd__o2bb2a_1 _17736_ (.A1_N(_09505_),
    .A2_N(_09507_),
    .B1(_09719_),
    .B2(_09722_),
    .X(_09723_));
 sky130_fd_sc_hd__a21o_1 _17737_ (.A1(_09719_),
    .A2(_09722_),
    .B1(_09723_),
    .X(_09724_));
 sky130_fd_sc_hd__xor2_1 _17738_ (.A(_09699_),
    .B(_09704_),
    .X(_09725_));
 sky130_fd_sc_hd__xnor2_2 _17739_ (.A(_09701_),
    .B(_09725_),
    .Y(_09726_));
 sky130_fd_sc_hd__inv_2 _17740_ (.A(_09413_),
    .Y(_09727_));
 sky130_fd_sc_hd__xnor2_1 _17741_ (.A(_09418_),
    .B(_09421_),
    .Y(_09728_));
 sky130_fd_sc_hd__mux2_1 _17742_ (.A0(_09505_),
    .A1(_09728_),
    .S(_09506_),
    .X(_09729_));
 sky130_fd_sc_hd__nor2_1 _17743_ (.A(_09418_),
    .B(_09421_),
    .Y(_09730_));
 sky130_fd_sc_hd__nand2_1 _17744_ (.A(_09424_),
    .B(_09730_),
    .Y(_09731_));
 sky130_fd_sc_hd__mux2_1 _17745_ (.A0(_09729_),
    .A1(_09731_),
    .S(_09503_),
    .X(_09732_));
 sky130_fd_sc_hd__o21a_1 _17746_ (.A1(_09727_),
    .A2(_09732_),
    .B1(_09492_),
    .X(_09733_));
 sky130_fd_sc_hd__a2bb2o_1 _17747_ (.A1_N(_09506_),
    .A2_N(_09728_),
    .B1(_09730_),
    .B2(_09510_),
    .X(_09734_));
 sky130_fd_sc_hd__nand2_1 _17748_ (.A(_09508_),
    .B(_09509_),
    .Y(_09735_));
 sky130_fd_sc_hd__mux2_1 _17749_ (.A0(_09734_),
    .A1(_09735_),
    .S(_09503_),
    .X(_09736_));
 sky130_fd_sc_hd__or2_1 _17750_ (.A(_09733_),
    .B(_09736_),
    .X(_09737_));
 sky130_fd_sc_hd__or2_1 _17751_ (.A(_09726_),
    .B(_09737_),
    .X(_09738_));
 sky130_fd_sc_hd__and2_1 _17752_ (.A(_09726_),
    .B(_09737_),
    .X(_09739_));
 sky130_fd_sc_hd__a21o_1 _17753_ (.A1(_09724_),
    .A2(_09738_),
    .B1(_09739_),
    .X(_09740_));
 sky130_fd_sc_hd__a21bo_1 _17754_ (.A1(_09513_),
    .A2(_09456_),
    .B1_N(_09467_),
    .X(_09741_));
 sky130_fd_sc_hd__o21ai_1 _17755_ (.A1(_09513_),
    .A2(_09456_),
    .B1(_09741_),
    .Y(_09742_));
 sky130_fd_sc_hd__xnor2_2 _17756_ (.A(_09726_),
    .B(_09737_),
    .Y(_09743_));
 sky130_fd_sc_hd__xnor2_1 _17757_ (.A(_09724_),
    .B(_09743_),
    .Y(_09744_));
 sky130_fd_sc_hd__a22o_1 _17758_ (.A1(_09718_),
    .A2(_09740_),
    .B1(_09742_),
    .B2(_09744_),
    .X(_09745_));
 sky130_fd_sc_hd__a211o_1 _17759_ (.A1(_09516_),
    .A2(_09517_),
    .B1(_09603_),
    .C1(_09745_),
    .X(_09746_));
 sky130_fd_sc_hd__and3_1 _17760_ (.A(_09718_),
    .B(_09726_),
    .C(_09737_),
    .X(_09747_));
 sky130_fd_sc_hd__a21bo_1 _17761_ (.A1(_09406_),
    .A2(_09368_),
    .B1_N(_09446_),
    .X(_09748_));
 sky130_fd_sc_hd__o21a_1 _17762_ (.A1(_09406_),
    .A2(_09368_),
    .B1(_09748_),
    .X(_09749_));
 sky130_fd_sc_hd__o21a_1 _17763_ (.A1(_09515_),
    .A2(_09749_),
    .B1(_09742_),
    .X(_09750_));
 sky130_fd_sc_hd__inv_2 _17764_ (.A(_09743_),
    .Y(_09751_));
 sky130_fd_sc_hd__a31o_1 _17765_ (.A1(_09716_),
    .A2(_09717_),
    .A3(_09738_),
    .B1(_09743_),
    .X(_09752_));
 sky130_fd_sc_hd__mux2_1 _17766_ (.A0(_09751_),
    .A1(_09752_),
    .S(_09724_),
    .X(_09753_));
 sky130_fd_sc_hd__nand2_1 _17767_ (.A(_09662_),
    .B(_09682_),
    .Y(_09754_));
 sky130_fd_sc_hd__o21bai_1 _17768_ (.A1(_09662_),
    .A2(_09682_),
    .B1_N(_09669_),
    .Y(_09755_));
 sky130_fd_sc_hd__nand2_1 _17769_ (.A(_09754_),
    .B(_09755_),
    .Y(_09756_));
 sky130_fd_sc_hd__nand2_1 _17770_ (.A(net424),
    .B(net319),
    .Y(_09757_));
 sky130_fd_sc_hd__nand2_1 _17771_ (.A(net375),
    .B(net361),
    .Y(_09758_));
 sky130_fd_sc_hd__nand2_1 _17772_ (.A(net379),
    .B(net355),
    .Y(_09759_));
 sky130_fd_sc_hd__xnor2_1 _17773_ (.A(_09758_),
    .B(_09759_),
    .Y(_09760_));
 sky130_fd_sc_hd__xnor2_2 _17774_ (.A(_09757_),
    .B(_09760_),
    .Y(_09761_));
 sky130_fd_sc_hd__nand2_1 _17775_ (.A(net378),
    .B(net359),
    .Y(_09762_));
 sky130_fd_sc_hd__o21a_1 _17776_ (.A1(_09636_),
    .A2(_09762_),
    .B1(_09637_),
    .X(_09763_));
 sky130_fd_sc_hd__a21o_1 _17777_ (.A1(_09636_),
    .A2(_09762_),
    .B1(_09763_),
    .X(_09764_));
 sky130_fd_sc_hd__nand2_1 _17778_ (.A(net426),
    .B(net315),
    .Y(_09765_));
 sky130_fd_sc_hd__xor2_1 _17779_ (.A(_09764_),
    .B(_09765_),
    .X(_09766_));
 sky130_fd_sc_hd__xnor2_2 _17780_ (.A(_09761_),
    .B(_09766_),
    .Y(_09767_));
 sky130_fd_sc_hd__nor2_1 _17781_ (.A(_09677_),
    .B(_09680_),
    .Y(_09768_));
 sky130_fd_sc_hd__nand2_1 _17782_ (.A(_09677_),
    .B(_09680_),
    .Y(_09769_));
 sky130_fd_sc_hd__o21ai_1 _17783_ (.A1(_09674_),
    .A2(_09768_),
    .B1(_09769_),
    .Y(_09770_));
 sky130_fd_sc_hd__nor2_2 _17784_ (.A(_09688_),
    .B(_09706_),
    .Y(_09771_));
 sky130_fd_sc_hd__xor2_1 _17785_ (.A(net378),
    .B(_09636_),
    .X(_09772_));
 sky130_fd_sc_hd__and3_1 _17786_ (.A(_09518_),
    .B(_09771_),
    .C(_09772_),
    .X(_09773_));
 sky130_fd_sc_hd__xnor2_1 _17787_ (.A(_09770_),
    .B(_09773_),
    .Y(_09774_));
 sky130_fd_sc_hd__xnor2_2 _17788_ (.A(_09767_),
    .B(_09774_),
    .Y(_09775_));
 sky130_fd_sc_hd__nand2_1 _17789_ (.A(net399),
    .B(net339),
    .Y(_09776_));
 sky130_fd_sc_hd__nand2_1 _17790_ (.A(net404),
    .B(net336),
    .Y(_09777_));
 sky130_fd_sc_hd__nand2_1 _17791_ (.A(net409),
    .B(net332),
    .Y(_09778_));
 sky130_fd_sc_hd__xor2_1 _17792_ (.A(_09777_),
    .B(_09778_),
    .X(_09779_));
 sky130_fd_sc_hd__xnor2_1 _17793_ (.A(_09776_),
    .B(_09779_),
    .Y(_09780_));
 sky130_fd_sc_hd__o21ai_1 _17794_ (.A1(_09649_),
    .A2(_09650_),
    .B1(_09648_),
    .Y(_09781_));
 sky130_fd_sc_hd__a21bo_1 _17795_ (.A1(_09649_),
    .A2(_09650_),
    .B1_N(_09781_),
    .X(_09782_));
 sky130_fd_sc_hd__nand2_1 _17796_ (.A(net413),
    .B(net329),
    .Y(_09783_));
 sky130_fd_sc_hd__nand2_1 _17797_ (.A(\top0.pid_d.mult0.a[3] ),
    .B(net326),
    .Y(_09784_));
 sky130_fd_sc_hd__xor2_1 _17798_ (.A(_09783_),
    .B(_09784_),
    .X(_09785_));
 sky130_fd_sc_hd__xnor2_2 _17799_ (.A(_09666_),
    .B(_09785_),
    .Y(_09786_));
 sky130_fd_sc_hd__xor2_1 _17800_ (.A(_09782_),
    .B(_09786_),
    .X(_09787_));
 sky130_fd_sc_hd__xnor2_1 _17801_ (.A(_09780_),
    .B(_09787_),
    .Y(_09788_));
 sky130_fd_sc_hd__or2_1 _17802_ (.A(_09652_),
    .B(_09660_),
    .X(_09789_));
 sky130_fd_sc_hd__a21o_1 _17803_ (.A1(_09652_),
    .A2(_09660_),
    .B1(_09655_),
    .X(_09790_));
 sky130_fd_sc_hd__nand2_1 _17804_ (.A(net384),
    .B(net350),
    .Y(_09791_));
 sky130_fd_sc_hd__nand2_1 _17805_ (.A(net388),
    .B(net346),
    .Y(_09792_));
 sky130_fd_sc_hd__nand2_1 _17806_ (.A(net393),
    .B(\top0.pid_d.mult0.b[4] ),
    .Y(_09793_));
 sky130_fd_sc_hd__xnor2_1 _17807_ (.A(_09792_),
    .B(_09793_),
    .Y(_09794_));
 sky130_fd_sc_hd__xnor2_2 _17808_ (.A(_09791_),
    .B(_09794_),
    .Y(_09795_));
 sky130_fd_sc_hd__nand4_1 _17809_ (.A(net409),
    .B(net404),
    .C(net335),
    .D(net337),
    .Y(_09796_));
 sky130_fd_sc_hd__a22oi_1 _17810_ (.A1(net409),
    .A2(net335),
    .B1(net337),
    .B2(net404),
    .Y(_09797_));
 sky130_fd_sc_hd__a21oi_2 _17811_ (.A1(_09658_),
    .A2(_09796_),
    .B1(_09797_),
    .Y(_09798_));
 sky130_fd_sc_hd__nand4_1 _17812_ (.A(net393),
    .B(net388),
    .C(net345),
    .D(net349),
    .Y(_09799_));
 sky130_fd_sc_hd__a22oi_1 _17813_ (.A1(net393),
    .A2(net345),
    .B1(net349),
    .B2(net388),
    .Y(_09800_));
 sky130_fd_sc_hd__a21oi_2 _17814_ (.A1(_09671_),
    .A2(_09799_),
    .B1(_09800_),
    .Y(_09801_));
 sky130_fd_sc_hd__xnor2_1 _17815_ (.A(_09798_),
    .B(_09801_),
    .Y(_09802_));
 sky130_fd_sc_hd__xnor2_1 _17816_ (.A(_09795_),
    .B(_09802_),
    .Y(_09803_));
 sky130_fd_sc_hd__and3_1 _17817_ (.A(_09789_),
    .B(_09790_),
    .C(_09803_),
    .X(_09804_));
 sky130_fd_sc_hd__a21o_1 _17818_ (.A1(_09789_),
    .A2(_09790_),
    .B1(_09803_),
    .X(_09805_));
 sky130_fd_sc_hd__and2b_1 _17819_ (.A_N(_09804_),
    .B(_09805_),
    .X(_09806_));
 sky130_fd_sc_hd__xnor2_1 _17820_ (.A(_09788_),
    .B(_09806_),
    .Y(_09807_));
 sky130_fd_sc_hd__xor2_1 _17821_ (.A(_09775_),
    .B(_09807_),
    .X(_09808_));
 sky130_fd_sc_hd__xnor2_2 _17822_ (.A(_09756_),
    .B(_09808_),
    .Y(_09809_));
 sky130_fd_sc_hd__and2b_1 _17823_ (.A_N(_09684_),
    .B(_09647_),
    .X(_09810_));
 sky130_fd_sc_hd__or2b_1 _17824_ (.A(_09647_),
    .B_N(_09684_),
    .X(_09811_));
 sky130_fd_sc_hd__o21a_1 _17825_ (.A1(_09810_),
    .A2(_09635_),
    .B1(_09811_),
    .X(_09812_));
 sky130_fd_sc_hd__or2b_1 _17826_ (.A(_09645_),
    .B_N(_09641_),
    .X(_09813_));
 sky130_fd_sc_hd__and2b_1 _17827_ (.A_N(_09641_),
    .B(_09645_),
    .X(_09814_));
 sky130_fd_sc_hd__a21o_1 _17828_ (.A1(_09644_),
    .A2(_09813_),
    .B1(_09814_),
    .X(_09815_));
 sky130_fd_sc_hd__xor2_1 _17829_ (.A(_09812_),
    .B(_09815_),
    .X(_09816_));
 sky130_fd_sc_hd__xnor2_1 _17830_ (.A(_09809_),
    .B(_09816_),
    .Y(_09817_));
 sky130_fd_sc_hd__a21o_1 _17831_ (.A1(_09702_),
    .A2(_09705_),
    .B1(_09713_),
    .X(_09818_));
 sky130_fd_sc_hd__a21oi_1 _17832_ (.A1(_09686_),
    .A2(_09818_),
    .B1(_09714_),
    .Y(_09819_));
 sky130_fd_sc_hd__o22a_1 _17833_ (.A1(_09817_),
    .A2(_09819_),
    .B1(_09718_),
    .B2(_09740_),
    .X(_09820_));
 sky130_fd_sc_hd__o31a_1 _17834_ (.A1(_09747_),
    .A2(_09750_),
    .A3(_09753_),
    .B1(_09820_),
    .X(_09821_));
 sky130_fd_sc_hd__and2_1 _17835_ (.A(_09817_),
    .B(_09819_),
    .X(_09822_));
 sky130_fd_sc_hd__a21o_1 _17836_ (.A1(_09746_),
    .A2(_09821_),
    .B1(_09822_),
    .X(_09823_));
 sky130_fd_sc_hd__nor2_1 _17837_ (.A(_09812_),
    .B(_09815_),
    .Y(_09824_));
 sky130_fd_sc_hd__nand2_1 _17838_ (.A(_09812_),
    .B(_09815_),
    .Y(_09825_));
 sky130_fd_sc_hd__o21ai_2 _17839_ (.A1(_09809_),
    .A2(_09824_),
    .B1(_09825_),
    .Y(_09826_));
 sky130_fd_sc_hd__nand2_2 _17840_ (.A(net329),
    .B(net408),
    .Y(_09827_));
 sky130_fd_sc_hd__nand2_1 _17841_ (.A(net326),
    .B(net414),
    .Y(_09828_));
 sky130_fd_sc_hd__nand2_1 _17842_ (.A(net322),
    .B(net417),
    .Y(_09829_));
 sky130_fd_sc_hd__xor2_1 _17843_ (.A(_09828_),
    .B(_09829_),
    .X(_09830_));
 sky130_fd_sc_hd__xnor2_2 _17844_ (.A(_09827_),
    .B(_09830_),
    .Y(_09831_));
 sky130_fd_sc_hd__o21bai_1 _17845_ (.A1(_09783_),
    .A2(_09784_),
    .B1_N(_09666_),
    .Y(_09832_));
 sky130_fd_sc_hd__a21bo_1 _17846_ (.A1(_09783_),
    .A2(_09784_),
    .B1_N(_09832_),
    .X(_09833_));
 sky130_fd_sc_hd__nand2_1 _17847_ (.A(net339),
    .B(net393),
    .Y(_09834_));
 sky130_fd_sc_hd__nand2_1 _17848_ (.A(net336),
    .B(net399),
    .Y(_09835_));
 sky130_fd_sc_hd__nand2_1 _17849_ (.A(net332),
    .B(net404),
    .Y(_09836_));
 sky130_fd_sc_hd__xnor2_1 _17850_ (.A(_09835_),
    .B(_09836_),
    .Y(_09837_));
 sky130_fd_sc_hd__xnor2_1 _17851_ (.A(_09834_),
    .B(_09837_),
    .Y(_09838_));
 sky130_fd_sc_hd__xnor2_1 _17852_ (.A(_09833_),
    .B(_09838_),
    .Y(_09839_));
 sky130_fd_sc_hd__xnor2_2 _17853_ (.A(_09831_),
    .B(_09839_),
    .Y(_09840_));
 sky130_fd_sc_hd__nand2_1 _17854_ (.A(_09782_),
    .B(_09786_),
    .Y(_09841_));
 sky130_fd_sc_hd__o21bai_1 _17855_ (.A1(_09782_),
    .A2(_09786_),
    .B1_N(_09780_),
    .Y(_09842_));
 sky130_fd_sc_hd__nand2_1 _17856_ (.A(_09841_),
    .B(_09842_),
    .Y(_09843_));
 sky130_fd_sc_hd__nand2_2 _17857_ (.A(net351),
    .B(net380),
    .Y(_09844_));
 sky130_fd_sc_hd__nand2_1 _17858_ (.A(net346),
    .B(net383),
    .Y(_09845_));
 sky130_fd_sc_hd__nand2_1 _17859_ (.A(net342),
    .B(net388),
    .Y(_09846_));
 sky130_fd_sc_hd__xnor2_1 _17860_ (.A(_09845_),
    .B(_09846_),
    .Y(_09847_));
 sky130_fd_sc_hd__xnor2_2 _17861_ (.A(_09844_),
    .B(_09847_),
    .Y(_09848_));
 sky130_fd_sc_hd__nand4_1 _17862_ (.A(net389),
    .B(net346),
    .C(net384),
    .D(net351),
    .Y(_09849_));
 sky130_fd_sc_hd__a22oi_1 _17863_ (.A1(net389),
    .A2(net346),
    .B1(net384),
    .B2(net351),
    .Y(_09850_));
 sky130_fd_sc_hd__a21oi_2 _17864_ (.A1(_09793_),
    .A2(_09849_),
    .B1(_09850_),
    .Y(_09851_));
 sky130_fd_sc_hd__nand4_1 _17865_ (.A(net404),
    .B(net336),
    .C(net399),
    .D(net339),
    .Y(_09852_));
 sky130_fd_sc_hd__a22oi_1 _17866_ (.A1(net404),
    .A2(net336),
    .B1(net399),
    .B2(net339),
    .Y(_09853_));
 sky130_fd_sc_hd__a21oi_2 _17867_ (.A1(_09778_),
    .A2(_09852_),
    .B1(_09853_),
    .Y(_09854_));
 sky130_fd_sc_hd__xor2_1 _17868_ (.A(_09851_),
    .B(_09854_),
    .X(_09855_));
 sky130_fd_sc_hd__xnor2_2 _17869_ (.A(_09848_),
    .B(_09855_),
    .Y(_09856_));
 sky130_fd_sc_hd__xnor2_1 _17870_ (.A(_09843_),
    .B(_09856_),
    .Y(_09857_));
 sky130_fd_sc_hd__xnor2_2 _17871_ (.A(_09840_),
    .B(_09857_),
    .Y(_09858_));
 sky130_fd_sc_hd__a21oi_1 _17872_ (.A1(_09788_),
    .A2(_09805_),
    .B1(_09804_),
    .Y(_09859_));
 sky130_fd_sc_hd__o21a_1 _17873_ (.A1(_09764_),
    .A2(_09761_),
    .B1(_09765_),
    .X(_09860_));
 sky130_fd_sc_hd__a21o_1 _17874_ (.A1(_09764_),
    .A2(_09761_),
    .B1(_09860_),
    .X(_09861_));
 sky130_fd_sc_hd__nand2_1 _17875_ (.A(net420),
    .B(net319),
    .Y(_09862_));
 sky130_fd_sc_hd__nand2_2 _17876_ (.A(net361),
    .B(net372),
    .Y(_09863_));
 sky130_fd_sc_hd__nand2_1 _17877_ (.A(net355),
    .B(net374),
    .Y(_09864_));
 sky130_fd_sc_hd__xnor2_1 _17878_ (.A(_09863_),
    .B(_09864_),
    .Y(_09865_));
 sky130_fd_sc_hd__xnor2_2 _17879_ (.A(_09862_),
    .B(_09865_),
    .Y(_09866_));
 sky130_fd_sc_hd__nand4_1 _17880_ (.A(net378),
    .B(net355),
    .C(net375),
    .D(net359),
    .Y(_09867_));
 sky130_fd_sc_hd__a22oi_1 _17881_ (.A1(net378),
    .A2(net355),
    .B1(net375),
    .B2(net359),
    .Y(_09868_));
 sky130_fd_sc_hd__a21oi_2 _17882_ (.A1(_09757_),
    .A2(_09867_),
    .B1(_09868_),
    .Y(_09869_));
 sky130_fd_sc_hd__nand2_1 _17883_ (.A(net426),
    .B(net313),
    .Y(_09870_));
 sky130_fd_sc_hd__nand2_1 _17884_ (.A(net424),
    .B(net315),
    .Y(_09871_));
 sky130_fd_sc_hd__xor2_2 _17885_ (.A(_09870_),
    .B(_09871_),
    .X(_09872_));
 sky130_fd_sc_hd__xor2_1 _17886_ (.A(_09869_),
    .B(_09872_),
    .X(_09873_));
 sky130_fd_sc_hd__xnor2_2 _17887_ (.A(_09866_),
    .B(_09873_),
    .Y(_09874_));
 sky130_fd_sc_hd__nand2_1 _17888_ (.A(_09798_),
    .B(_09801_),
    .Y(_09875_));
 sky130_fd_sc_hd__nor2_1 _17889_ (.A(_09798_),
    .B(_09801_),
    .Y(_09876_));
 sky130_fd_sc_hd__a21oi_2 _17890_ (.A1(_09795_),
    .A2(_09875_),
    .B1(_09876_),
    .Y(_09877_));
 sky130_fd_sc_hd__xor2_1 _17891_ (.A(_09874_),
    .B(_09877_),
    .X(_09878_));
 sky130_fd_sc_hd__xnor2_1 _17892_ (.A(_09861_),
    .B(_09878_),
    .Y(_09879_));
 sky130_fd_sc_hd__nor2_1 _17893_ (.A(_09859_),
    .B(_09879_),
    .Y(_09880_));
 sky130_fd_sc_hd__nand2_1 _17894_ (.A(_09859_),
    .B(_09879_),
    .Y(_09881_));
 sky130_fd_sc_hd__and2b_1 _17895_ (.A_N(_09880_),
    .B(_09881_),
    .X(_09882_));
 sky130_fd_sc_hd__xnor2_2 _17896_ (.A(_09858_),
    .B(_09882_),
    .Y(_09883_));
 sky130_fd_sc_hd__a21o_1 _17897_ (.A1(_09767_),
    .A2(_09773_),
    .B1(_09770_),
    .X(_09884_));
 sky130_fd_sc_hd__o21a_2 _17898_ (.A1(_09767_),
    .A2(_09773_),
    .B1(_09884_),
    .X(_09885_));
 sky130_fd_sc_hd__and3_1 _17899_ (.A(_09754_),
    .B(_09755_),
    .C(_09775_),
    .X(_09886_));
 sky130_fd_sc_hd__a21o_1 _17900_ (.A1(_09754_),
    .A2(_09755_),
    .B1(_09775_),
    .X(_09887_));
 sky130_fd_sc_hd__o21a_1 _17901_ (.A1(_09807_),
    .A2(_09886_),
    .B1(_09887_),
    .X(_09888_));
 sky130_fd_sc_hd__xor2_1 _17902_ (.A(_09885_),
    .B(_09888_),
    .X(_09889_));
 sky130_fd_sc_hd__xnor2_1 _17903_ (.A(_09883_),
    .B(_09889_),
    .Y(_09890_));
 sky130_fd_sc_hd__xnor2_1 _17904_ (.A(_09826_),
    .B(_09890_),
    .Y(_09891_));
 sky130_fd_sc_hd__nand2_1 _17905_ (.A(_09823_),
    .B(_09891_),
    .Y(_09892_));
 sky130_fd_sc_hd__or2_2 _17906_ (.A(_09823_),
    .B(_09891_),
    .X(_09893_));
 sky130_fd_sc_hd__and4_1 _17907_ (.A(net439),
    .B(_09339_),
    .C(_09892_),
    .D(_09893_),
    .X(_09894_));
 sky130_fd_sc_hd__inv_2 _17908_ (.A(\top0.pid_d.curr_int[0] ),
    .Y(_09895_));
 sky130_fd_sc_hd__nor2_1 _17909_ (.A(_09895_),
    .B(_07138_),
    .Y(_09896_));
 sky130_fd_sc_hd__mux2_1 _17910_ (.A0(_09896_),
    .A1(_09895_),
    .S(\top0.pid_d.out[0] ),
    .X(_09897_));
 sky130_fd_sc_hd__a22o_1 _17911_ (.A1(\top0.pid_d.out[0] ),
    .A2(_07138_),
    .B1(_09897_),
    .B2(net434),
    .X(_09898_));
 sky130_fd_sc_hd__o21a_1 _17912_ (.A1(_09894_),
    .A2(_09898_),
    .B1(_07710_),
    .X(_00245_));
 sky130_fd_sc_hd__xor2_1 _17913_ (.A(\top0.pid_d.out[1] ),
    .B(\top0.pid_d.curr_int[1] ),
    .X(_09899_));
 sky130_fd_sc_hd__a21o_1 _17914_ (.A1(\top0.pid_d.out[0] ),
    .A2(\top0.pid_d.curr_int[0] ),
    .B1(_09899_),
    .X(_09900_));
 sky130_fd_sc_hd__nand3_1 _17915_ (.A(\top0.pid_d.out[0] ),
    .B(\top0.pid_d.curr_int[0] ),
    .C(_09899_),
    .Y(_09901_));
 sky130_fd_sc_hd__or2_1 _17916_ (.A(_09826_),
    .B(_09890_),
    .X(_09902_));
 sky130_fd_sc_hd__nand2_2 _17917_ (.A(net339),
    .B(net388),
    .Y(_09903_));
 sky130_fd_sc_hd__nand2_1 _17918_ (.A(net336),
    .B(net393),
    .Y(_09904_));
 sky130_fd_sc_hd__nand2_1 _17919_ (.A(net332),
    .B(net399),
    .Y(_09905_));
 sky130_fd_sc_hd__xnor2_1 _17920_ (.A(_09904_),
    .B(_09905_),
    .Y(_09906_));
 sky130_fd_sc_hd__xnor2_2 _17921_ (.A(_09903_),
    .B(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__o21ai_1 _17922_ (.A1(_09827_),
    .A2(_09828_),
    .B1(_09829_),
    .Y(_09908_));
 sky130_fd_sc_hd__a21bo_1 _17923_ (.A1(_09827_),
    .A2(_09828_),
    .B1_N(_09908_),
    .X(_09909_));
 sky130_fd_sc_hd__nand2_2 _17924_ (.A(net1022),
    .B(net404),
    .Y(_09910_));
 sky130_fd_sc_hd__nand2_1 _17925_ (.A(net325),
    .B(net408),
    .Y(_09911_));
 sky130_fd_sc_hd__nand2_1 _17926_ (.A(net1023),
    .B(net413),
    .Y(_09912_));
 sky130_fd_sc_hd__xnor2_1 _17927_ (.A(_09911_),
    .B(_09912_),
    .Y(_09913_));
 sky130_fd_sc_hd__xnor2_2 _17928_ (.A(_09910_),
    .B(_09913_),
    .Y(_09914_));
 sky130_fd_sc_hd__xnor2_1 _17929_ (.A(_09909_),
    .B(_09914_),
    .Y(_09915_));
 sky130_fd_sc_hd__xnor2_2 _17930_ (.A(_09907_),
    .B(_09915_),
    .Y(_09916_));
 sky130_fd_sc_hd__o21ba_1 _17931_ (.A1(_09833_),
    .A2(_09838_),
    .B1_N(_09831_),
    .X(_09917_));
 sky130_fd_sc_hd__a21o_1 _17932_ (.A1(_09833_),
    .A2(_09838_),
    .B1(_09917_),
    .X(_09918_));
 sky130_fd_sc_hd__nand2_2 _17933_ (.A(net351),
    .B(net375),
    .Y(_09919_));
 sky130_fd_sc_hd__nand2_1 _17934_ (.A(net346),
    .B(net380),
    .Y(_09920_));
 sky130_fd_sc_hd__nand2_1 _17935_ (.A(net342),
    .B(net383),
    .Y(_09921_));
 sky130_fd_sc_hd__xnor2_1 _17936_ (.A(_09920_),
    .B(_09921_),
    .Y(_09922_));
 sky130_fd_sc_hd__xnor2_2 _17937_ (.A(_09919_),
    .B(_09922_),
    .Y(_09923_));
 sky130_fd_sc_hd__o21a_1 _17938_ (.A1(_09844_),
    .A2(_09845_),
    .B1(_09846_),
    .X(_09924_));
 sky130_fd_sc_hd__a21oi_2 _17939_ (.A1(_09844_),
    .A2(_09845_),
    .B1(_09924_),
    .Y(_09925_));
 sky130_fd_sc_hd__o21a_1 _17940_ (.A1(_09834_),
    .A2(_09835_),
    .B1(_09836_),
    .X(_09926_));
 sky130_fd_sc_hd__a21oi_2 _17941_ (.A1(_09834_),
    .A2(_09835_),
    .B1(_09926_),
    .Y(_09927_));
 sky130_fd_sc_hd__xnor2_1 _17942_ (.A(_09925_),
    .B(_09927_),
    .Y(_09928_));
 sky130_fd_sc_hd__xnor2_2 _17943_ (.A(_09923_),
    .B(_09928_),
    .Y(_09929_));
 sky130_fd_sc_hd__xor2_1 _17944_ (.A(_09918_),
    .B(_09929_),
    .X(_09930_));
 sky130_fd_sc_hd__xnor2_2 _17945_ (.A(_09916_),
    .B(_09930_),
    .Y(_09931_));
 sky130_fd_sc_hd__a21o_1 _17946_ (.A1(_09841_),
    .A2(_09842_),
    .B1(_09856_),
    .X(_09932_));
 sky130_fd_sc_hd__and3_1 _17947_ (.A(_09841_),
    .B(_09842_),
    .C(_09856_),
    .X(_09933_));
 sky130_fd_sc_hd__a21oi_1 _17948_ (.A1(_09840_),
    .A2(_09932_),
    .B1(_09933_),
    .Y(_09934_));
 sky130_fd_sc_hd__nand2_1 _17949_ (.A(net361),
    .B(net370),
    .Y(_09935_));
 sky130_fd_sc_hd__nand2_1 _17950_ (.A(net355),
    .B(net372),
    .Y(_09936_));
 sky130_fd_sc_hd__nand2_1 _17951_ (.A(net416),
    .B(net319),
    .Y(_09937_));
 sky130_fd_sc_hd__xnor2_1 _17952_ (.A(_09936_),
    .B(_09937_),
    .Y(_09938_));
 sky130_fd_sc_hd__xnor2_1 _17953_ (.A(_09935_),
    .B(_09938_),
    .Y(_09939_));
 sky130_fd_sc_hd__o21a_1 _17954_ (.A1(_09863_),
    .A2(_09864_),
    .B1(_09862_),
    .X(_09940_));
 sky130_fd_sc_hd__a21o_1 _17955_ (.A1(_09863_),
    .A2(_09864_),
    .B1(_09940_),
    .X(_09941_));
 sky130_fd_sc_hd__nand2_2 _17956_ (.A(net426),
    .B(net310),
    .Y(_09942_));
 sky130_fd_sc_hd__nand2_1 _17957_ (.A(net420),
    .B(net315),
    .Y(_09943_));
 sky130_fd_sc_hd__nand2_1 _17958_ (.A(net424),
    .B(net313),
    .Y(_09944_));
 sky130_fd_sc_hd__xnor2_1 _17959_ (.A(_09943_),
    .B(_09944_),
    .Y(_09945_));
 sky130_fd_sc_hd__xnor2_2 _17960_ (.A(_09942_),
    .B(_09945_),
    .Y(_09946_));
 sky130_fd_sc_hd__xnor2_1 _17961_ (.A(_09941_),
    .B(_09946_),
    .Y(_09947_));
 sky130_fd_sc_hd__xnor2_1 _17962_ (.A(_09939_),
    .B(_09947_),
    .Y(_09948_));
 sky130_fd_sc_hd__nand2_1 _17963_ (.A(_09869_),
    .B(_09872_),
    .Y(_09949_));
 sky130_fd_sc_hd__nor2_1 _17964_ (.A(_09869_),
    .B(_09872_),
    .Y(_09950_));
 sky130_fd_sc_hd__a21oi_2 _17965_ (.A1(_09866_),
    .A2(_09949_),
    .B1(_09950_),
    .Y(_09951_));
 sky130_fd_sc_hd__nand2_1 _17966_ (.A(_09851_),
    .B(_09854_),
    .Y(_09952_));
 sky130_fd_sc_hd__nor2_1 _17967_ (.A(_09851_),
    .B(_09854_),
    .Y(_09953_));
 sky130_fd_sc_hd__a21oi_2 _17968_ (.A1(_09848_),
    .A2(_09952_),
    .B1(_09953_),
    .Y(_09954_));
 sky130_fd_sc_hd__xnor2_1 _17969_ (.A(_09951_),
    .B(_09954_),
    .Y(_09955_));
 sky130_fd_sc_hd__xnor2_1 _17970_ (.A(_09948_),
    .B(_09955_),
    .Y(_09956_));
 sky130_fd_sc_hd__nor2_1 _17971_ (.A(_09934_),
    .B(_09956_),
    .Y(_09957_));
 sky130_fd_sc_hd__nand2_1 _17972_ (.A(_09934_),
    .B(_09956_),
    .Y(_09958_));
 sky130_fd_sc_hd__or2b_1 _17973_ (.A(_09957_),
    .B_N(_09958_),
    .X(_09959_));
 sky130_fd_sc_hd__xnor2_2 _17974_ (.A(_09931_),
    .B(_09959_),
    .Y(_09960_));
 sky130_fd_sc_hd__a21o_1 _17975_ (.A1(_09858_),
    .A2(_09881_),
    .B1(_09880_),
    .X(_09961_));
 sky130_fd_sc_hd__nand2_1 _17976_ (.A(_09874_),
    .B(_09877_),
    .Y(_09962_));
 sky130_fd_sc_hd__nor2_1 _17977_ (.A(_09874_),
    .B(_09877_),
    .Y(_09963_));
 sky130_fd_sc_hd__a21o_1 _17978_ (.A1(_09861_),
    .A2(_09962_),
    .B1(_09963_),
    .X(_09964_));
 sky130_fd_sc_hd__inv_2 _17979_ (.A(net314),
    .Y(_09965_));
 sky130_fd_sc_hd__inv_2 _17980_ (.A(net311),
    .Y(_09966_));
 sky130_fd_sc_hd__nor2_4 _17981_ (.A(_09965_),
    .B(_09966_),
    .Y(_09967_));
 sky130_fd_sc_hd__and3_1 _17982_ (.A(net424),
    .B(net426),
    .C(_09967_),
    .X(_09968_));
 sky130_fd_sc_hd__xnor2_2 _17983_ (.A(_09964_),
    .B(_09968_),
    .Y(_09969_));
 sky130_fd_sc_hd__xor2_1 _17984_ (.A(_09961_),
    .B(_09969_),
    .X(_09970_));
 sky130_fd_sc_hd__xnor2_1 _17985_ (.A(_09960_),
    .B(_09970_),
    .Y(_09971_));
 sky130_fd_sc_hd__inv_2 _17986_ (.A(_09971_),
    .Y(_09972_));
 sky130_fd_sc_hd__a21o_1 _17987_ (.A1(_09885_),
    .A2(_09883_),
    .B1(_09888_),
    .X(_09973_));
 sky130_fd_sc_hd__o21ai_2 _17988_ (.A1(_09885_),
    .A2(_09883_),
    .B1(_09973_),
    .Y(_09974_));
 sky130_fd_sc_hd__xnor2_1 _17989_ (.A(_09972_),
    .B(_09974_),
    .Y(_09975_));
 sky130_fd_sc_hd__xnor2_2 _17990_ (.A(_09902_),
    .B(_09975_),
    .Y(_09976_));
 sky130_fd_sc_hd__xor2_2 _17991_ (.A(_09893_),
    .B(_09976_),
    .X(_09977_));
 sky130_fd_sc_hd__a32o_1 _17992_ (.A1(net434),
    .A2(_09900_),
    .A3(_09901_),
    .B1(_09977_),
    .B2(net439),
    .X(_09978_));
 sky130_fd_sc_hd__mux2_1 _17993_ (.A0(\top0.pid_d.out[1] ),
    .A1(_09978_),
    .S(net14),
    .X(_09979_));
 sky130_fd_sc_hd__and2_1 _17994_ (.A(net1018),
    .B(_09979_),
    .X(_09980_));
 sky130_fd_sc_hd__clkbuf_1 _17995_ (.A(_09980_),
    .X(_00246_));
 sky130_fd_sc_hd__a22o_1 _17996_ (.A1(\top0.pid_d.out[0] ),
    .A2(\top0.pid_d.curr_int[0] ),
    .B1(\top0.pid_d.curr_int[1] ),
    .B2(\top0.pid_d.out[1] ),
    .X(_09981_));
 sky130_fd_sc_hd__or2_1 _17997_ (.A(\top0.pid_d.out[1] ),
    .B(\top0.pid_d.curr_int[1] ),
    .X(_09982_));
 sky130_fd_sc_hd__and2_1 _17998_ (.A(_09981_),
    .B(_09982_),
    .X(_09983_));
 sky130_fd_sc_hd__xnor2_1 _17999_ (.A(\top0.pid_d.out[2] ),
    .B(\top0.pid_d.curr_int[2] ),
    .Y(_09984_));
 sky130_fd_sc_hd__xnor2_1 _18000_ (.A(_09983_),
    .B(_09984_),
    .Y(_09985_));
 sky130_fd_sc_hd__nand2_2 _18001_ (.A(net361),
    .B(net366),
    .Y(_09986_));
 sky130_fd_sc_hd__nand2_1 _18002_ (.A(net351),
    .B(net372),
    .Y(_09987_));
 sky130_fd_sc_hd__nand2_1 _18003_ (.A(net355),
    .B(net370),
    .Y(_09988_));
 sky130_fd_sc_hd__xor2_1 _18004_ (.A(_09987_),
    .B(_09988_),
    .X(_09989_));
 sky130_fd_sc_hd__xnor2_2 _18005_ (.A(_09986_),
    .B(_09989_),
    .Y(_09990_));
 sky130_fd_sc_hd__o21ai_1 _18006_ (.A1(_09935_),
    .A2(_09936_),
    .B1(_09937_),
    .Y(_09991_));
 sky130_fd_sc_hd__a21bo_1 _18007_ (.A1(_09935_),
    .A2(_09936_),
    .B1_N(_09991_),
    .X(_09992_));
 sky130_fd_sc_hd__nand2_1 _18008_ (.A(net421),
    .B(net313),
    .Y(_09993_));
 sky130_fd_sc_hd__nand2_1 _18009_ (.A(net411),
    .B(net319),
    .Y(_09994_));
 sky130_fd_sc_hd__nand2_1 _18010_ (.A(net416),
    .B(net315),
    .Y(_09995_));
 sky130_fd_sc_hd__xnor2_1 _18011_ (.A(_09994_),
    .B(_09995_),
    .Y(_09996_));
 sky130_fd_sc_hd__xnor2_1 _18012_ (.A(_09993_),
    .B(_09996_),
    .Y(_09997_));
 sky130_fd_sc_hd__nor2_1 _18013_ (.A(_09992_),
    .B(_09997_),
    .Y(_09998_));
 sky130_fd_sc_hd__nand2_1 _18014_ (.A(_09992_),
    .B(_09997_),
    .Y(_09999_));
 sky130_fd_sc_hd__and2b_1 _18015_ (.A_N(_09998_),
    .B(_09999_),
    .X(_10000_));
 sky130_fd_sc_hd__xnor2_2 _18016_ (.A(_09990_),
    .B(_10000_),
    .Y(_10001_));
 sky130_fd_sc_hd__a21bo_1 _18017_ (.A1(_09925_),
    .A2(_09927_),
    .B1_N(_09923_),
    .X(_10002_));
 sky130_fd_sc_hd__o21ai_1 _18018_ (.A1(_09925_),
    .A2(_09927_),
    .B1(_10002_),
    .Y(_10003_));
 sky130_fd_sc_hd__o21a_1 _18019_ (.A1(_09941_),
    .A2(_09946_),
    .B1(_09939_),
    .X(_10004_));
 sky130_fd_sc_hd__a21o_1 _18020_ (.A1(_09941_),
    .A2(_09946_),
    .B1(_10004_),
    .X(_10005_));
 sky130_fd_sc_hd__xnor2_1 _18021_ (.A(_10003_),
    .B(_10005_),
    .Y(_10006_));
 sky130_fd_sc_hd__xnor2_2 _18022_ (.A(_10001_),
    .B(_10006_),
    .Y(_10007_));
 sky130_fd_sc_hd__a21o_1 _18023_ (.A1(_09918_),
    .A2(_09929_),
    .B1(_09916_),
    .X(_10008_));
 sky130_fd_sc_hd__o21ai_2 _18024_ (.A1(_09918_),
    .A2(_09929_),
    .B1(_10008_),
    .Y(_10009_));
 sky130_fd_sc_hd__nand2_1 _18025_ (.A(net325),
    .B(net404),
    .Y(_10010_));
 sky130_fd_sc_hd__nand2_1 _18026_ (.A(net321),
    .B(net409),
    .Y(_10011_));
 sky130_fd_sc_hd__xnor2_1 _18027_ (.A(_10010_),
    .B(_10011_),
    .Y(_10012_));
 sky130_fd_sc_hd__xnor2_2 _18028_ (.A(net307),
    .B(_10012_),
    .Y(_10013_));
 sky130_fd_sc_hd__o21ai_1 _18029_ (.A1(_09910_),
    .A2(_09911_),
    .B1(_09912_),
    .Y(_10014_));
 sky130_fd_sc_hd__a21bo_1 _18030_ (.A1(_09910_),
    .A2(_09911_),
    .B1_N(_10014_),
    .X(_10015_));
 sky130_fd_sc_hd__nand2_2 _18031_ (.A(net335),
    .B(net389),
    .Y(_10016_));
 sky130_fd_sc_hd__nand2_1 _18032_ (.A(net1022),
    .B(net398),
    .Y(_10017_));
 sky130_fd_sc_hd__nand2_1 _18033_ (.A(net332),
    .B(net393),
    .Y(_10018_));
 sky130_fd_sc_hd__xnor2_1 _18034_ (.A(_10017_),
    .B(_10018_),
    .Y(_10019_));
 sky130_fd_sc_hd__xnor2_2 _18035_ (.A(_10016_),
    .B(_10019_),
    .Y(_10020_));
 sky130_fd_sc_hd__xnor2_1 _18036_ (.A(_10015_),
    .B(_10020_),
    .Y(_10021_));
 sky130_fd_sc_hd__xnor2_2 _18037_ (.A(_10013_),
    .B(_10021_),
    .Y(_10022_));
 sky130_fd_sc_hd__o21a_1 _18038_ (.A1(_09909_),
    .A2(_09914_),
    .B1(_09907_),
    .X(_10023_));
 sky130_fd_sc_hd__a21o_1 _18039_ (.A1(_09909_),
    .A2(_09914_),
    .B1(_10023_),
    .X(_10024_));
 sky130_fd_sc_hd__nand2_2 _18040_ (.A(net346),
    .B(net375),
    .Y(_10025_));
 sky130_fd_sc_hd__nand2_1 _18041_ (.A(\top0.pid_d.mult0.b[5] ),
    .B(net383),
    .Y(_10026_));
 sky130_fd_sc_hd__nand2_1 _18042_ (.A(net342),
    .B(net380),
    .Y(_10027_));
 sky130_fd_sc_hd__xnor2_1 _18043_ (.A(_10026_),
    .B(_10027_),
    .Y(_10028_));
 sky130_fd_sc_hd__xnor2_2 _18044_ (.A(_10025_),
    .B(_10028_),
    .Y(_10029_));
 sky130_fd_sc_hd__o21a_1 _18045_ (.A1(_09919_),
    .A2(_09920_),
    .B1(_09921_),
    .X(_10030_));
 sky130_fd_sc_hd__a21oi_2 _18046_ (.A1(_09919_),
    .A2(_09920_),
    .B1(_10030_),
    .Y(_10031_));
 sky130_fd_sc_hd__o21a_1 _18047_ (.A1(_09903_),
    .A2(_09904_),
    .B1(_09905_),
    .X(_10032_));
 sky130_fd_sc_hd__a21oi_2 _18048_ (.A1(_09903_),
    .A2(_09904_),
    .B1(_10032_),
    .Y(_10033_));
 sky130_fd_sc_hd__xnor2_1 _18049_ (.A(_10031_),
    .B(_10033_),
    .Y(_10034_));
 sky130_fd_sc_hd__xnor2_2 _18050_ (.A(_10029_),
    .B(_10034_),
    .Y(_10035_));
 sky130_fd_sc_hd__xnor2_1 _18051_ (.A(_10024_),
    .B(_10035_),
    .Y(_10036_));
 sky130_fd_sc_hd__xnor2_2 _18052_ (.A(_10022_),
    .B(_10036_),
    .Y(_10037_));
 sky130_fd_sc_hd__xor2_1 _18053_ (.A(_10009_),
    .B(_10037_),
    .X(_10038_));
 sky130_fd_sc_hd__xnor2_2 _18054_ (.A(_10007_),
    .B(_10038_),
    .Y(_10039_));
 sky130_fd_sc_hd__o21ai_1 _18055_ (.A1(_09931_),
    .A2(_09957_),
    .B1(_09958_),
    .Y(_10040_));
 sky130_fd_sc_hd__a21bo_1 _18056_ (.A1(_09951_),
    .A2(_09954_),
    .B1_N(_09948_),
    .X(_10041_));
 sky130_fd_sc_hd__o21ai_1 _18057_ (.A1(_09951_),
    .A2(_09954_),
    .B1(_10041_),
    .Y(_10042_));
 sky130_fd_sc_hd__o21a_1 _18058_ (.A1(_09942_),
    .A2(_09944_),
    .B1(_09943_),
    .X(_10043_));
 sky130_fd_sc_hd__a21o_1 _18059_ (.A1(_09942_),
    .A2(_09944_),
    .B1(_10043_),
    .X(_10044_));
 sky130_fd_sc_hd__nand2_1 _18060_ (.A(_09616_),
    .B(net307),
    .Y(_10045_));
 sky130_fd_sc_hd__nand2_1 _18061_ (.A(net424),
    .B(net310),
    .Y(_10046_));
 sky130_fd_sc_hd__xnor2_1 _18062_ (.A(_10045_),
    .B(_10046_),
    .Y(_10047_));
 sky130_fd_sc_hd__xnor2_1 _18063_ (.A(_10044_),
    .B(_10047_),
    .Y(_10048_));
 sky130_fd_sc_hd__xnor2_1 _18064_ (.A(_10042_),
    .B(_10048_),
    .Y(_10049_));
 sky130_fd_sc_hd__nand2_1 _18065_ (.A(_10040_),
    .B(_10049_),
    .Y(_10050_));
 sky130_fd_sc_hd__or2_1 _18066_ (.A(_10040_),
    .B(_10049_),
    .X(_10051_));
 sky130_fd_sc_hd__nand2_1 _18067_ (.A(_10050_),
    .B(_10051_),
    .Y(_10052_));
 sky130_fd_sc_hd__xnor2_2 _18068_ (.A(_10039_),
    .B(_10052_),
    .Y(_10053_));
 sky130_fd_sc_hd__and2b_1 _18069_ (.A_N(_09964_),
    .B(_09968_),
    .X(_10054_));
 sky130_fd_sc_hd__a21bo_1 _18070_ (.A1(_09960_),
    .A2(_09969_),
    .B1_N(_09961_),
    .X(_10055_));
 sky130_fd_sc_hd__o21a_1 _18071_ (.A1(_09960_),
    .A2(_09969_),
    .B1(_10055_),
    .X(_10056_));
 sky130_fd_sc_hd__xor2_1 _18072_ (.A(_10054_),
    .B(_10056_),
    .X(_10057_));
 sky130_fd_sc_hd__xnor2_1 _18073_ (.A(_10053_),
    .B(_10057_),
    .Y(_10058_));
 sky130_fd_sc_hd__a21o_1 _18074_ (.A1(_09972_),
    .A2(_09974_),
    .B1(_09902_),
    .X(_10059_));
 sky130_fd_sc_hd__a211o_1 _18075_ (.A1(_09972_),
    .A2(_09974_),
    .B1(_09822_),
    .C1(_09891_),
    .X(_10060_));
 sky130_fd_sc_hd__a21o_1 _18076_ (.A1(_09746_),
    .A2(_09821_),
    .B1(_10060_),
    .X(_10061_));
 sky130_fd_sc_hd__or2_1 _18077_ (.A(_09972_),
    .B(_09974_),
    .X(_10062_));
 sky130_fd_sc_hd__and4_1 _18078_ (.A(_10058_),
    .B(_10059_),
    .C(_10061_),
    .D(_10062_),
    .X(_10063_));
 sky130_fd_sc_hd__a31o_1 _18079_ (.A1(_10059_),
    .A2(_10061_),
    .A3(_10062_),
    .B1(_10058_),
    .X(_10064_));
 sky130_fd_sc_hd__and2b_1 _18080_ (.A_N(_10063_),
    .B(_10064_),
    .X(_10065_));
 sky130_fd_sc_hd__a221o_1 _18081_ (.A1(net434),
    .A2(_09985_),
    .B1(_10065_),
    .B2(net439),
    .C1(_07138_),
    .X(_10066_));
 sky130_fd_sc_hd__clkbuf_4 _18082_ (.A(net1019),
    .X(_10067_));
 sky130_fd_sc_hd__o211a_1 _18083_ (.A1(\top0.pid_d.out[2] ),
    .A2(_09339_),
    .B1(_10066_),
    .C1(_10067_),
    .X(_00247_));
 sky130_fd_sc_hd__a31o_1 _18084_ (.A1(\top0.pid_d.curr_int[2] ),
    .A2(_09981_),
    .A3(_09982_),
    .B1(\top0.pid_d.out[2] ),
    .X(_10068_));
 sky130_fd_sc_hd__o21a_1 _18085_ (.A1(\top0.pid_d.curr_int[2] ),
    .A2(_09983_),
    .B1(_10068_),
    .X(_10069_));
 sky130_fd_sc_hd__xnor2_1 _18086_ (.A(\top0.pid_d.out[3] ),
    .B(\top0.pid_d.curr_int[3] ),
    .Y(_10070_));
 sky130_fd_sc_hd__xnor2_1 _18087_ (.A(_10069_),
    .B(_10070_),
    .Y(_10071_));
 sky130_fd_sc_hd__a21o_1 _18088_ (.A1(_10053_),
    .A2(_10056_),
    .B1(_10054_),
    .X(_10072_));
 sky130_fd_sc_hd__o21a_1 _18089_ (.A1(_10053_),
    .A2(_10056_),
    .B1(_10072_),
    .X(_10073_));
 sky130_fd_sc_hd__xor2_4 _18090_ (.A(net356),
    .B(net361),
    .X(_10074_));
 sky130_fd_sc_hd__nand2_2 _18091_ (.A(net365),
    .B(_10074_),
    .Y(_10075_));
 sky130_fd_sc_hd__nand2_1 _18092_ (.A(net405),
    .B(net318),
    .Y(_10076_));
 sky130_fd_sc_hd__xor2_2 _18093_ (.A(_10075_),
    .B(_10076_),
    .X(_10077_));
 sky130_fd_sc_hd__o21ai_1 _18094_ (.A1(_09986_),
    .A2(_09988_),
    .B1(_09987_),
    .Y(_10078_));
 sky130_fd_sc_hd__a21bo_1 _18095_ (.A1(_09986_),
    .A2(_09988_),
    .B1_N(_10078_),
    .X(_10079_));
 sky130_fd_sc_hd__nand2_1 _18096_ (.A(net416),
    .B(net313),
    .Y(_10080_));
 sky130_fd_sc_hd__nand2_1 _18097_ (.A(net411),
    .B(net315),
    .Y(_10081_));
 sky130_fd_sc_hd__xor2_1 _18098_ (.A(_10080_),
    .B(_10081_),
    .X(_10082_));
 sky130_fd_sc_hd__nand2_1 _18099_ (.A(net421),
    .B(net310),
    .Y(_10083_));
 sky130_fd_sc_hd__xor2_1 _18100_ (.A(_10082_),
    .B(_10083_),
    .X(_10084_));
 sky130_fd_sc_hd__nor2_1 _18101_ (.A(_10079_),
    .B(_10084_),
    .Y(_10085_));
 sky130_fd_sc_hd__nand2_1 _18102_ (.A(_10079_),
    .B(_10084_),
    .Y(_10086_));
 sky130_fd_sc_hd__and2b_1 _18103_ (.A_N(_10085_),
    .B(_10086_),
    .X(_10087_));
 sky130_fd_sc_hd__xnor2_2 _18104_ (.A(_10077_),
    .B(_10087_),
    .Y(_10088_));
 sky130_fd_sc_hd__a21bo_1 _18105_ (.A1(_10031_),
    .A2(_10033_),
    .B1_N(_10029_),
    .X(_10089_));
 sky130_fd_sc_hd__o21ai_1 _18106_ (.A1(_10031_),
    .A2(_10033_),
    .B1(_10089_),
    .Y(_10090_));
 sky130_fd_sc_hd__a21oi_1 _18107_ (.A1(_09990_),
    .A2(_09999_),
    .B1(_09998_),
    .Y(_10091_));
 sky130_fd_sc_hd__nand2_1 _18108_ (.A(_10090_),
    .B(_10091_),
    .Y(_10092_));
 sky130_fd_sc_hd__or2_1 _18109_ (.A(_10090_),
    .B(_10091_),
    .X(_10093_));
 sky130_fd_sc_hd__nand2_1 _18110_ (.A(_10092_),
    .B(_10093_),
    .Y(_10094_));
 sky130_fd_sc_hd__xnor2_2 _18111_ (.A(_10088_),
    .B(_10094_),
    .Y(_10095_));
 sky130_fd_sc_hd__a21bo_1 _18112_ (.A1(_10024_),
    .A2(_10035_),
    .B1_N(_10022_),
    .X(_10096_));
 sky130_fd_sc_hd__o21a_1 _18113_ (.A1(_10024_),
    .A2(_10035_),
    .B1(_10096_),
    .X(_10097_));
 sky130_fd_sc_hd__nand2_1 _18114_ (.A(net338),
    .B(net378),
    .Y(_10098_));
 sky130_fd_sc_hd__nand2_1 _18115_ (.A(net332),
    .B(net389),
    .Y(_10099_));
 sky130_fd_sc_hd__nand2_1 _18116_ (.A(net334),
    .B(net383),
    .Y(_10100_));
 sky130_fd_sc_hd__xnor2_1 _18117_ (.A(_10099_),
    .B(_10100_),
    .Y(_10101_));
 sky130_fd_sc_hd__xnor2_1 _18118_ (.A(_10098_),
    .B(_10101_),
    .Y(_10102_));
 sky130_fd_sc_hd__inv_2 _18119_ (.A(net307),
    .Y(_10103_));
 sky130_fd_sc_hd__o21ai_1 _18120_ (.A1(_10103_),
    .A2(_10010_),
    .B1(_10011_),
    .Y(_10104_));
 sky130_fd_sc_hd__a21bo_1 _18121_ (.A1(_10103_),
    .A2(_10010_),
    .B1_N(_10104_),
    .X(_10105_));
 sky130_fd_sc_hd__nand2_1 _18122_ (.A(net328),
    .B(net394),
    .Y(_10106_));
 sky130_fd_sc_hd__nand2_1 _18123_ (.A(net1023),
    .B(net403),
    .Y(_10107_));
 sky130_fd_sc_hd__nand2_1 _18124_ (.A(net325),
    .B(net398),
    .Y(_10108_));
 sky130_fd_sc_hd__xnor2_1 _18125_ (.A(_10107_),
    .B(_10108_),
    .Y(_10109_));
 sky130_fd_sc_hd__xnor2_2 _18126_ (.A(_10106_),
    .B(_10109_),
    .Y(_10110_));
 sky130_fd_sc_hd__xnor2_1 _18127_ (.A(_10105_),
    .B(_10110_),
    .Y(_10111_));
 sky130_fd_sc_hd__xnor2_1 _18128_ (.A(_10102_),
    .B(_10111_),
    .Y(_10112_));
 sky130_fd_sc_hd__o21ba_1 _18129_ (.A1(_10015_),
    .A2(_10020_),
    .B1_N(_10013_),
    .X(_10113_));
 sky130_fd_sc_hd__a21o_1 _18130_ (.A1(_10015_),
    .A2(_10020_),
    .B1(_10113_),
    .X(_10114_));
 sky130_fd_sc_hd__nand2_2 _18131_ (.A(net350),
    .B(\top0.pid_d.mult0.a[14] ),
    .Y(_10115_));
 sky130_fd_sc_hd__nand2_1 _18132_ (.A(net342),
    .B(net375),
    .Y(_10116_));
 sky130_fd_sc_hd__nand2_1 _18133_ (.A(net346),
    .B(net372),
    .Y(_10117_));
 sky130_fd_sc_hd__xnor2_1 _18134_ (.A(_10116_),
    .B(_10117_),
    .Y(_10118_));
 sky130_fd_sc_hd__xnor2_2 _18135_ (.A(_10115_),
    .B(_10118_),
    .Y(_10119_));
 sky130_fd_sc_hd__o21a_1 _18136_ (.A1(_10025_),
    .A2(_10027_),
    .B1(_10026_),
    .X(_10120_));
 sky130_fd_sc_hd__a21oi_2 _18137_ (.A1(_10025_),
    .A2(_10027_),
    .B1(_10120_),
    .Y(_10121_));
 sky130_fd_sc_hd__o21a_1 _18138_ (.A1(_10016_),
    .A2(_10018_),
    .B1(_10017_),
    .X(_10122_));
 sky130_fd_sc_hd__a21oi_2 _18139_ (.A1(_10016_),
    .A2(_10018_),
    .B1(_10122_),
    .Y(_10123_));
 sky130_fd_sc_hd__xnor2_1 _18140_ (.A(_10121_),
    .B(_10123_),
    .Y(_10124_));
 sky130_fd_sc_hd__xnor2_2 _18141_ (.A(_10119_),
    .B(_10124_),
    .Y(_10125_));
 sky130_fd_sc_hd__xnor2_1 _18142_ (.A(_10114_),
    .B(_10125_),
    .Y(_10126_));
 sky130_fd_sc_hd__xnor2_1 _18143_ (.A(_10112_),
    .B(_10126_),
    .Y(_10127_));
 sky130_fd_sc_hd__nor2_1 _18144_ (.A(_10097_),
    .B(_10127_),
    .Y(_10128_));
 sky130_fd_sc_hd__and2_1 _18145_ (.A(_10097_),
    .B(_10127_),
    .X(_10129_));
 sky130_fd_sc_hd__nor2_1 _18146_ (.A(_10128_),
    .B(_10129_),
    .Y(_10130_));
 sky130_fd_sc_hd__xnor2_2 _18147_ (.A(_10095_),
    .B(_10130_),
    .Y(_10131_));
 sky130_fd_sc_hd__a21bo_1 _18148_ (.A1(_10009_),
    .A2(_10037_),
    .B1_N(_10007_),
    .X(_10132_));
 sky130_fd_sc_hd__o21a_1 _18149_ (.A1(_10009_),
    .A2(_10037_),
    .B1(_10132_),
    .X(_10133_));
 sky130_fd_sc_hd__o21a_1 _18150_ (.A1(_10001_),
    .A2(_10005_),
    .B1(_10003_),
    .X(_10134_));
 sky130_fd_sc_hd__a21o_1 _18151_ (.A1(_10001_),
    .A2(_10005_),
    .B1(_10134_),
    .X(_10135_));
 sky130_fd_sc_hd__a21o_1 _18152_ (.A1(_10044_),
    .A2(_10045_),
    .B1(_10046_),
    .X(_10136_));
 sky130_fd_sc_hd__o21ai_1 _18153_ (.A1(_10044_),
    .A2(_10045_),
    .B1(_10136_),
    .Y(_10137_));
 sky130_fd_sc_hd__nand2_1 _18154_ (.A(_09993_),
    .B(_09994_),
    .Y(_10138_));
 sky130_fd_sc_hd__nor2_1 _18155_ (.A(_09993_),
    .B(_09994_),
    .Y(_10139_));
 sky130_fd_sc_hd__a31o_1 _18156_ (.A1(net416),
    .A2(net315),
    .A3(_10138_),
    .B1(_10139_),
    .X(_10140_));
 sky130_fd_sc_hd__and3_1 _18157_ (.A(_09593_),
    .B(net307),
    .C(_10140_),
    .X(_10141_));
 sky130_fd_sc_hd__a21oi_1 _18158_ (.A1(_09593_),
    .A2(net307),
    .B1(_10140_),
    .Y(_10142_));
 sky130_fd_sc_hd__nor2_1 _18159_ (.A(_10141_),
    .B(_10142_),
    .Y(_10143_));
 sky130_fd_sc_hd__nor2_1 _18160_ (.A(_10137_),
    .B(_10143_),
    .Y(_10144_));
 sky130_fd_sc_hd__nand2_1 _18161_ (.A(_10137_),
    .B(_10143_),
    .Y(_10145_));
 sky130_fd_sc_hd__and2b_1 _18162_ (.A_N(_10144_),
    .B(_10145_),
    .X(_10146_));
 sky130_fd_sc_hd__xnor2_2 _18163_ (.A(_10135_),
    .B(_10146_),
    .Y(_10147_));
 sky130_fd_sc_hd__xor2_1 _18164_ (.A(_10133_),
    .B(_10147_),
    .X(_10148_));
 sky130_fd_sc_hd__xnor2_1 _18165_ (.A(_10131_),
    .B(_10148_),
    .Y(_10149_));
 sky130_fd_sc_hd__nor2_1 _18166_ (.A(_10040_),
    .B(_10049_),
    .Y(_10150_));
 sky130_fd_sc_hd__a21oi_2 _18167_ (.A1(_10039_),
    .A2(_10050_),
    .B1(_10150_),
    .Y(_10151_));
 sky130_fd_sc_hd__or2_1 _18168_ (.A(_10042_),
    .B(_10048_),
    .X(_10152_));
 sky130_fd_sc_hd__xnor2_1 _18169_ (.A(_10151_),
    .B(_10152_),
    .Y(_10153_));
 sky130_fd_sc_hd__xnor2_1 _18170_ (.A(_10149_),
    .B(_10153_),
    .Y(_10154_));
 sky130_fd_sc_hd__xnor2_1 _18171_ (.A(_10073_),
    .B(_10154_),
    .Y(_10155_));
 sky130_fd_sc_hd__xnor2_1 _18172_ (.A(_10064_),
    .B(_10155_),
    .Y(_10156_));
 sky130_fd_sc_hd__a221o_1 _18173_ (.A1(net434),
    .A2(_10071_),
    .B1(_10156_),
    .B2(net439),
    .C1(_07138_),
    .X(_10157_));
 sky130_fd_sc_hd__o211a_1 _18174_ (.A1(\top0.pid_d.out[3] ),
    .A2(_09339_),
    .B1(_10157_),
    .C1(_10067_),
    .X(_00248_));
 sky130_fd_sc_hd__a21o_1 _18175_ (.A1(\top0.pid_d.curr_int[3] ),
    .A2(_10069_),
    .B1(\top0.pid_d.out[3] ),
    .X(_10158_));
 sky130_fd_sc_hd__o21a_1 _18176_ (.A1(\top0.pid_d.curr_int[3] ),
    .A2(_10069_),
    .B1(_10158_),
    .X(_10159_));
 sky130_fd_sc_hd__xnor2_1 _18177_ (.A(\top0.pid_d.out[4] ),
    .B(\top0.pid_d.curr_int[4] ),
    .Y(_10160_));
 sky130_fd_sc_hd__xnor2_1 _18178_ (.A(_10159_),
    .B(_10160_),
    .Y(_10161_));
 sky130_fd_sc_hd__inv_2 _18179_ (.A(_10154_),
    .Y(_10162_));
 sky130_fd_sc_hd__nand2_1 _18180_ (.A(_10073_),
    .B(_10162_),
    .Y(_10163_));
 sky130_fd_sc_hd__nor2_1 _18181_ (.A(_10073_),
    .B(_10162_),
    .Y(_10164_));
 sky130_fd_sc_hd__a21oi_2 _18182_ (.A1(_10064_),
    .A2(_10163_),
    .B1(_10164_),
    .Y(_10165_));
 sky130_fd_sc_hd__o21a_1 _18183_ (.A1(_10151_),
    .A2(_10152_),
    .B1(_10149_),
    .X(_10166_));
 sky130_fd_sc_hd__a21o_1 _18184_ (.A1(_10151_),
    .A2(_10152_),
    .B1(_10166_),
    .X(_10167_));
 sky130_fd_sc_hd__nand2_2 _18185_ (.A(net338),
    .B(net376),
    .Y(_10168_));
 sky130_fd_sc_hd__nand2_1 _18186_ (.A(net331),
    .B(net382),
    .Y(_10169_));
 sky130_fd_sc_hd__nand2_1 _18187_ (.A(net334),
    .B(net378),
    .Y(_10170_));
 sky130_fd_sc_hd__xor2_1 _18188_ (.A(_10169_),
    .B(_10170_),
    .X(_10171_));
 sky130_fd_sc_hd__xnor2_2 _18189_ (.A(_10168_),
    .B(_10171_),
    .Y(_10172_));
 sky130_fd_sc_hd__o21ai_1 _18190_ (.A1(_10106_),
    .A2(_10108_),
    .B1(_10107_),
    .Y(_10173_));
 sky130_fd_sc_hd__a21bo_1 _18191_ (.A1(_10106_),
    .A2(_10108_),
    .B1_N(_10173_),
    .X(_10174_));
 sky130_fd_sc_hd__nand2_1 _18192_ (.A(net328),
    .B(net388),
    .Y(_10175_));
 sky130_fd_sc_hd__nand2_1 _18193_ (.A(net1023),
    .B(net395),
    .Y(_10176_));
 sky130_fd_sc_hd__nand2_1 _18194_ (.A(net325),
    .B(net394),
    .Y(_10177_));
 sky130_fd_sc_hd__xnor2_1 _18195_ (.A(_10176_),
    .B(_10177_),
    .Y(_10178_));
 sky130_fd_sc_hd__xnor2_1 _18196_ (.A(_10175_),
    .B(_10178_),
    .Y(_10179_));
 sky130_fd_sc_hd__nor2_1 _18197_ (.A(_10174_),
    .B(_10179_),
    .Y(_10180_));
 sky130_fd_sc_hd__nand2_1 _18198_ (.A(_10174_),
    .B(_10179_),
    .Y(_10181_));
 sky130_fd_sc_hd__or2b_1 _18199_ (.A(_10180_),
    .B_N(_10181_),
    .X(_10182_));
 sky130_fd_sc_hd__xor2_2 _18200_ (.A(_10172_),
    .B(_10182_),
    .X(_10183_));
 sky130_fd_sc_hd__o21a_1 _18201_ (.A1(_10105_),
    .A2(_10110_),
    .B1(_10102_),
    .X(_10184_));
 sky130_fd_sc_hd__a21o_1 _18202_ (.A1(_10105_),
    .A2(_10110_),
    .B1(_10184_),
    .X(_10185_));
 sky130_fd_sc_hd__nand2_1 _18203_ (.A(net350),
    .B(net366),
    .Y(_10186_));
 sky130_fd_sc_hd__nand2_1 _18204_ (.A(\top0.pid_d.mult0.b[4] ),
    .B(net372),
    .Y(_10187_));
 sky130_fd_sc_hd__nand2_1 _18205_ (.A(net345),
    .B(net370),
    .Y(_10188_));
 sky130_fd_sc_hd__xnor2_1 _18206_ (.A(_10187_),
    .B(_10188_),
    .Y(_10189_));
 sky130_fd_sc_hd__xnor2_1 _18207_ (.A(_10186_),
    .B(_10189_),
    .Y(_10190_));
 sky130_fd_sc_hd__o21a_1 _18208_ (.A1(_10115_),
    .A2(_10117_),
    .B1(_10116_),
    .X(_10191_));
 sky130_fd_sc_hd__a21oi_2 _18209_ (.A1(_10115_),
    .A2(_10117_),
    .B1(_10191_),
    .Y(_10192_));
 sky130_fd_sc_hd__o21a_1 _18210_ (.A1(_10098_),
    .A2(_10100_),
    .B1(_10099_),
    .X(_10193_));
 sky130_fd_sc_hd__a21oi_2 _18211_ (.A1(_10098_),
    .A2(_10100_),
    .B1(_10193_),
    .Y(_10194_));
 sky130_fd_sc_hd__xnor2_1 _18212_ (.A(_10192_),
    .B(_10194_),
    .Y(_10195_));
 sky130_fd_sc_hd__xnor2_1 _18213_ (.A(_10190_),
    .B(_10195_),
    .Y(_10196_));
 sky130_fd_sc_hd__nor2_1 _18214_ (.A(_10185_),
    .B(_10196_),
    .Y(_10197_));
 sky130_fd_sc_hd__and2_1 _18215_ (.A(_10185_),
    .B(_10196_),
    .X(_10198_));
 sky130_fd_sc_hd__or2_1 _18216_ (.A(_10197_),
    .B(_10198_),
    .X(_10199_));
 sky130_fd_sc_hd__xnor2_2 _18217_ (.A(_10183_),
    .B(_10199_),
    .Y(_10200_));
 sky130_fd_sc_hd__a21o_1 _18218_ (.A1(_10114_),
    .A2(_10125_),
    .B1(_10112_),
    .X(_10201_));
 sky130_fd_sc_hd__o21a_1 _18219_ (.A1(_10114_),
    .A2(_10125_),
    .B1(_10201_),
    .X(_10202_));
 sky130_fd_sc_hd__nor2_2 _18220_ (.A(net354),
    .B(net358),
    .Y(_10203_));
 sky130_fd_sc_hd__o21ai_1 _18221_ (.A1(net405),
    .A2(_10203_),
    .B1(_09363_),
    .Y(_10204_));
 sky130_fd_sc_hd__and3_1 _18222_ (.A(net405),
    .B(_09353_),
    .C(_09363_),
    .X(_10205_));
 sky130_fd_sc_hd__a31o_1 _18223_ (.A1(net400),
    .A2(net366),
    .A3(_10204_),
    .B1(_10205_),
    .X(_10206_));
 sky130_fd_sc_hd__nand2_1 _18224_ (.A(net401),
    .B(net319),
    .Y(_10207_));
 sky130_fd_sc_hd__o21ai_4 _18225_ (.A1(net356),
    .A2(net360),
    .B1(net365),
    .Y(_10208_));
 sky130_fd_sc_hd__a22o_2 _18226_ (.A1(net319),
    .A2(_10206_),
    .B1(_10207_),
    .B2(_10208_),
    .X(_10209_));
 sky130_fd_sc_hd__nand2_1 _18227_ (.A(net405),
    .B(net315),
    .Y(_10210_));
 sky130_fd_sc_hd__nand2_1 _18228_ (.A(net410),
    .B(net313),
    .Y(_10211_));
 sky130_fd_sc_hd__xnor2_2 _18229_ (.A(_10210_),
    .B(_10211_),
    .Y(_10212_));
 sky130_fd_sc_hd__nand2_2 _18230_ (.A(net415),
    .B(\top0.pid_d.mult0.b[14] ),
    .Y(_10213_));
 sky130_fd_sc_hd__xnor2_4 _18231_ (.A(_10212_),
    .B(_10213_),
    .Y(_10214_));
 sky130_fd_sc_hd__xor2_4 _18232_ (.A(_10209_),
    .B(_10214_),
    .X(_10215_));
 sky130_fd_sc_hd__o21ai_1 _18233_ (.A1(_10077_),
    .A2(_10085_),
    .B1(_10086_),
    .Y(_10216_));
 sky130_fd_sc_hd__a21bo_1 _18234_ (.A1(_10121_),
    .A2(_10123_),
    .B1_N(_10119_),
    .X(_10217_));
 sky130_fd_sc_hd__o21a_1 _18235_ (.A1(_10121_),
    .A2(_10123_),
    .B1(_10217_),
    .X(_10218_));
 sky130_fd_sc_hd__xnor2_1 _18236_ (.A(_10216_),
    .B(_10218_),
    .Y(_10219_));
 sky130_fd_sc_hd__xnor2_2 _18237_ (.A(_10215_),
    .B(_10219_),
    .Y(_10220_));
 sky130_fd_sc_hd__xnor2_1 _18238_ (.A(_10202_),
    .B(_10220_),
    .Y(_10221_));
 sky130_fd_sc_hd__xnor2_2 _18239_ (.A(_10200_),
    .B(_10221_),
    .Y(_10222_));
 sky130_fd_sc_hd__or2_1 _18240_ (.A(_10097_),
    .B(_10127_),
    .X(_10223_));
 sky130_fd_sc_hd__a21o_1 _18241_ (.A1(_10095_),
    .A2(_10223_),
    .B1(_10129_),
    .X(_10224_));
 sky130_fd_sc_hd__a21bo_1 _18242_ (.A1(_10088_),
    .A2(_10093_),
    .B1_N(_10092_),
    .X(_10225_));
 sky130_fd_sc_hd__a32o_1 _18243_ (.A1(net416),
    .A2(net410),
    .A3(_09967_),
    .B1(\top0.pid_d.mult0.b[15] ),
    .B2(_09567_),
    .X(_10226_));
 sky130_fd_sc_hd__a31o_1 _18244_ (.A1(net421),
    .A2(net310),
    .A3(_10082_),
    .B1(_10226_),
    .X(_10227_));
 sky130_fd_sc_hd__nand2_2 _18245_ (.A(net307),
    .B(_09967_),
    .Y(_10228_));
 sky130_fd_sc_hd__or4bb_2 _18246_ (.A(net421),
    .B(_10228_),
    .C_N(net416),
    .D_N(net411),
    .X(_10229_));
 sky130_fd_sc_hd__nand2_1 _18247_ (.A(_10227_),
    .B(_10229_),
    .Y(_10230_));
 sky130_fd_sc_hd__xor2_1 _18248_ (.A(_10141_),
    .B(_10230_),
    .X(_10231_));
 sky130_fd_sc_hd__xnor2_1 _18249_ (.A(_10225_),
    .B(_10231_),
    .Y(_10232_));
 sky130_fd_sc_hd__and2_1 _18250_ (.A(_10224_),
    .B(_10232_),
    .X(_10233_));
 sky130_fd_sc_hd__or2_1 _18251_ (.A(_10224_),
    .B(_10232_),
    .X(_10234_));
 sky130_fd_sc_hd__and2b_1 _18252_ (.A_N(_10233_),
    .B(_10234_),
    .X(_10235_));
 sky130_fd_sc_hd__xnor2_2 _18253_ (.A(_10222_),
    .B(_10235_),
    .Y(_10236_));
 sky130_fd_sc_hd__a21o_1 _18254_ (.A1(_10131_),
    .A2(_10147_),
    .B1(_10133_),
    .X(_10237_));
 sky130_fd_sc_hd__o21ai_2 _18255_ (.A1(_10131_),
    .A2(_10147_),
    .B1(_10237_),
    .Y(_10238_));
 sky130_fd_sc_hd__a21o_1 _18256_ (.A1(_10135_),
    .A2(_10145_),
    .B1(_10144_),
    .X(_10239_));
 sky130_fd_sc_hd__xor2_1 _18257_ (.A(_10238_),
    .B(_10239_),
    .X(_10240_));
 sky130_fd_sc_hd__xnor2_2 _18258_ (.A(_10236_),
    .B(_10240_),
    .Y(_10241_));
 sky130_fd_sc_hd__xnor2_1 _18259_ (.A(_10167_),
    .B(_10241_),
    .Y(_10242_));
 sky130_fd_sc_hd__xnor2_1 _18260_ (.A(_10165_),
    .B(_10242_),
    .Y(_10243_));
 sky130_fd_sc_hd__a221o_1 _18261_ (.A1(net434),
    .A2(_10161_),
    .B1(_10243_),
    .B2(net436),
    .C1(_07138_),
    .X(_10244_));
 sky130_fd_sc_hd__o211a_1 _18262_ (.A1(\top0.pid_d.out[4] ),
    .A2(_09339_),
    .B1(_10244_),
    .C1(_10067_),
    .X(_00249_));
 sky130_fd_sc_hd__a21o_1 _18263_ (.A1(\top0.pid_d.curr_int[4] ),
    .A2(_10159_),
    .B1(\top0.pid_d.out[4] ),
    .X(_10245_));
 sky130_fd_sc_hd__o21ai_2 _18264_ (.A1(\top0.pid_d.curr_int[4] ),
    .A2(_10159_),
    .B1(_10245_),
    .Y(_10246_));
 sky130_fd_sc_hd__xnor2_1 _18265_ (.A(\top0.pid_d.out[5] ),
    .B(\top0.pid_d.curr_int[5] ),
    .Y(_10247_));
 sky130_fd_sc_hd__nand2_1 _18266_ (.A(_10246_),
    .B(_10247_),
    .Y(_10248_));
 sky130_fd_sc_hd__or2_1 _18267_ (.A(_10246_),
    .B(_10247_),
    .X(_10249_));
 sky130_fd_sc_hd__nand2_1 _18268_ (.A(_10167_),
    .B(_10241_),
    .Y(_10250_));
 sky130_fd_sc_hd__nor2_1 _18269_ (.A(_10167_),
    .B(_10241_),
    .Y(_10251_));
 sky130_fd_sc_hd__a21o_1 _18270_ (.A1(_10165_),
    .A2(_10250_),
    .B1(_10251_),
    .X(_10252_));
 sky130_fd_sc_hd__nor2_1 _18271_ (.A(_09353_),
    .B(_09364_),
    .Y(_10253_));
 sky130_fd_sc_hd__a31o_1 _18272_ (.A1(net406),
    .A2(_09353_),
    .A3(_10074_),
    .B1(_10253_),
    .X(_10254_));
 sky130_fd_sc_hd__and2_2 _18273_ (.A(net318),
    .B(net365),
    .X(_10255_));
 sky130_fd_sc_hd__o2bb2a_1 _18274_ (.A1_N(_10254_),
    .A2_N(_10255_),
    .B1(_10214_),
    .B2(_10209_),
    .X(_10256_));
 sky130_fd_sc_hd__o21ai_1 _18275_ (.A1(net401),
    .A2(_10203_),
    .B1(_09363_),
    .Y(_10257_));
 sky130_fd_sc_hd__a32o_1 _18276_ (.A1(net397),
    .A2(net366),
    .A3(_10257_),
    .B1(_09399_),
    .B2(_09363_),
    .X(_10258_));
 sky130_fd_sc_hd__nand2_1 _18277_ (.A(net396),
    .B(net317),
    .Y(_10259_));
 sky130_fd_sc_hd__a22o_1 _18278_ (.A1(net317),
    .A2(_10258_),
    .B1(_10259_),
    .B2(_10208_),
    .X(_10260_));
 sky130_fd_sc_hd__nand2_1 _18279_ (.A(net406),
    .B(net312),
    .Y(_10261_));
 sky130_fd_sc_hd__nand2_1 _18280_ (.A(net402),
    .B(net314),
    .Y(_10262_));
 sky130_fd_sc_hd__xor2_2 _18281_ (.A(_10261_),
    .B(_10262_),
    .X(_10263_));
 sky130_fd_sc_hd__nand2_1 _18282_ (.A(net411),
    .B(net310),
    .Y(_10264_));
 sky130_fd_sc_hd__xor2_2 _18283_ (.A(_10263_),
    .B(_10264_),
    .X(_10265_));
 sky130_fd_sc_hd__xor2_2 _18284_ (.A(_10260_),
    .B(_10265_),
    .X(_10266_));
 sky130_fd_sc_hd__a21bo_1 _18285_ (.A1(_10192_),
    .A2(_10194_),
    .B1_N(_10190_),
    .X(_10267_));
 sky130_fd_sc_hd__o21a_1 _18286_ (.A1(_10192_),
    .A2(_10194_),
    .B1(_10267_),
    .X(_10268_));
 sky130_fd_sc_hd__xnor2_1 _18287_ (.A(_10266_),
    .B(_10268_),
    .Y(_10269_));
 sky130_fd_sc_hd__xnor2_1 _18288_ (.A(_10256_),
    .B(_10269_),
    .Y(_10270_));
 sky130_fd_sc_hd__nand2_1 _18289_ (.A(net338),
    .B(net373),
    .Y(_10271_));
 sky130_fd_sc_hd__nand2_1 _18290_ (.A(net331),
    .B(net378),
    .Y(_10272_));
 sky130_fd_sc_hd__nand2_1 _18291_ (.A(net334),
    .B(net376),
    .Y(_10273_));
 sky130_fd_sc_hd__xor2_1 _18292_ (.A(_10272_),
    .B(_10273_),
    .X(_10274_));
 sky130_fd_sc_hd__xnor2_2 _18293_ (.A(_10271_),
    .B(_10274_),
    .Y(_10275_));
 sky130_fd_sc_hd__o21ai_1 _18294_ (.A1(_10175_),
    .A2(_10177_),
    .B1(_10176_),
    .Y(_10276_));
 sky130_fd_sc_hd__a21bo_1 _18295_ (.A1(_10175_),
    .A2(_10177_),
    .B1_N(_10276_),
    .X(_10277_));
 sky130_fd_sc_hd__nand2_1 _18296_ (.A(net329),
    .B(net382),
    .Y(_10278_));
 sky130_fd_sc_hd__nand2_1 _18297_ (.A(net1023),
    .B(net391),
    .Y(_10279_));
 sky130_fd_sc_hd__nand2_1 _18298_ (.A(net325),
    .B(net386),
    .Y(_10280_));
 sky130_fd_sc_hd__xnor2_1 _18299_ (.A(_10279_),
    .B(_10280_),
    .Y(_10281_));
 sky130_fd_sc_hd__xnor2_1 _18300_ (.A(_10278_),
    .B(_10281_),
    .Y(_10282_));
 sky130_fd_sc_hd__nor2_1 _18301_ (.A(_10277_),
    .B(_10282_),
    .Y(_10283_));
 sky130_fd_sc_hd__nand2_1 _18302_ (.A(_10277_),
    .B(_10282_),
    .Y(_10284_));
 sky130_fd_sc_hd__or2b_1 _18303_ (.A(_10283_),
    .B_N(_10284_),
    .X(_10285_));
 sky130_fd_sc_hd__xnor2_2 _18304_ (.A(_10275_),
    .B(_10285_),
    .Y(_10286_));
 sky130_fd_sc_hd__o21ai_2 _18305_ (.A1(_10172_),
    .A2(_10180_),
    .B1(_10181_),
    .Y(_10287_));
 sky130_fd_sc_hd__nand2_1 _18306_ (.A(net341),
    .B(net369),
    .Y(_10288_));
 sky130_fd_sc_hd__xor2_1 _18307_ (.A(net344),
    .B(net348),
    .X(_10289_));
 sky130_fd_sc_hd__nand2_1 _18308_ (.A(net364),
    .B(_10289_),
    .Y(_10290_));
 sky130_fd_sc_hd__xor2_2 _18309_ (.A(_10288_),
    .B(_10290_),
    .X(_10291_));
 sky130_fd_sc_hd__o21a_1 _18310_ (.A1(_10186_),
    .A2(_10188_),
    .B1(_10187_),
    .X(_10292_));
 sky130_fd_sc_hd__a21o_1 _18311_ (.A1(_10186_),
    .A2(_10188_),
    .B1(_10292_),
    .X(_10293_));
 sky130_fd_sc_hd__o21a_1 _18312_ (.A1(_10168_),
    .A2(_10170_),
    .B1(_10169_),
    .X(_10294_));
 sky130_fd_sc_hd__a21o_1 _18313_ (.A1(_10168_),
    .A2(_10170_),
    .B1(_10294_),
    .X(_10295_));
 sky130_fd_sc_hd__xnor2_1 _18314_ (.A(_10293_),
    .B(_10295_),
    .Y(_10296_));
 sky130_fd_sc_hd__xnor2_2 _18315_ (.A(_10291_),
    .B(_10296_),
    .Y(_10297_));
 sky130_fd_sc_hd__xor2_1 _18316_ (.A(_10287_),
    .B(_10297_),
    .X(_10298_));
 sky130_fd_sc_hd__xnor2_1 _18317_ (.A(_10286_),
    .B(_10298_),
    .Y(_10299_));
 sky130_fd_sc_hd__o21bai_1 _18318_ (.A1(_10183_),
    .A2(_10198_),
    .B1_N(_10197_),
    .Y(_10300_));
 sky130_fd_sc_hd__nor2_1 _18319_ (.A(_10299_),
    .B(_10300_),
    .Y(_10301_));
 sky130_fd_sc_hd__nand2_1 _18320_ (.A(_10299_),
    .B(_10300_),
    .Y(_10302_));
 sky130_fd_sc_hd__or2b_1 _18321_ (.A(_10301_),
    .B_N(_10302_),
    .X(_10303_));
 sky130_fd_sc_hd__xnor2_1 _18322_ (.A(_10270_),
    .B(_10303_),
    .Y(_10304_));
 sky130_fd_sc_hd__o21a_1 _18323_ (.A1(_10202_),
    .A2(_10220_),
    .B1(_10200_),
    .X(_10305_));
 sky130_fd_sc_hd__a21oi_2 _18324_ (.A1(_10202_),
    .A2(_10220_),
    .B1(_10305_),
    .Y(_10306_));
 sky130_fd_sc_hd__a21bo_1 _18325_ (.A1(_10215_),
    .A2(_10218_),
    .B1_N(_10216_),
    .X(_10307_));
 sky130_fd_sc_hd__o21ai_2 _18326_ (.A1(_10215_),
    .A2(_10218_),
    .B1(_10307_),
    .Y(_10308_));
 sky130_fd_sc_hd__and3_1 _18327_ (.A(net411),
    .B(net406),
    .C(_09967_),
    .X(_10309_));
 sky130_fd_sc_hd__xnor2_1 _18328_ (.A(_10103_),
    .B(_10309_),
    .Y(_10310_));
 sky130_fd_sc_hd__inv_2 _18329_ (.A(net310),
    .Y(_10311_));
 sky130_fd_sc_hd__o21ai_1 _18330_ (.A1(_10311_),
    .A2(_10210_),
    .B1(_10211_),
    .Y(_10312_));
 sky130_fd_sc_hd__a21boi_1 _18331_ (.A1(_10311_),
    .A2(_10210_),
    .B1_N(_10312_),
    .Y(_10313_));
 sky130_fd_sc_hd__mux2_1 _18332_ (.A0(_10310_),
    .A1(_10313_),
    .S(net416),
    .X(_10314_));
 sky130_fd_sc_hd__xnor2_1 _18333_ (.A(_10229_),
    .B(_10314_),
    .Y(_10315_));
 sky130_fd_sc_hd__xnor2_2 _18334_ (.A(_10308_),
    .B(_10315_),
    .Y(_10316_));
 sky130_fd_sc_hd__xnor2_1 _18335_ (.A(_10306_),
    .B(_10316_),
    .Y(_10317_));
 sky130_fd_sc_hd__xnor2_1 _18336_ (.A(_10304_),
    .B(_10317_),
    .Y(_10318_));
 sky130_fd_sc_hd__a21o_1 _18337_ (.A1(_10222_),
    .A2(_10234_),
    .B1(_10233_),
    .X(_10319_));
 sky130_fd_sc_hd__o21ba_1 _18338_ (.A1(_10225_),
    .A2(_10230_),
    .B1_N(_10141_),
    .X(_10320_));
 sky130_fd_sc_hd__a21o_1 _18339_ (.A1(_10225_),
    .A2(_10230_),
    .B1(_10320_),
    .X(_10321_));
 sky130_fd_sc_hd__or2_1 _18340_ (.A(_10319_),
    .B(_10321_),
    .X(_10322_));
 sky130_fd_sc_hd__nand2_1 _18341_ (.A(_10319_),
    .B(_10321_),
    .Y(_10323_));
 sky130_fd_sc_hd__nand2_1 _18342_ (.A(_10322_),
    .B(_10323_),
    .Y(_10324_));
 sky130_fd_sc_hd__xnor2_1 _18343_ (.A(_10318_),
    .B(_10324_),
    .Y(_10325_));
 sky130_fd_sc_hd__inv_2 _18344_ (.A(_10325_),
    .Y(_10326_));
 sky130_fd_sc_hd__o21ba_1 _18345_ (.A1(_10238_),
    .A2(_10239_),
    .B1_N(_10236_),
    .X(_10327_));
 sky130_fd_sc_hd__a21o_1 _18346_ (.A1(_10238_),
    .A2(_10239_),
    .B1(_10327_),
    .X(_10328_));
 sky130_fd_sc_hd__inv_2 _18347_ (.A(_10328_),
    .Y(_10329_));
 sky130_fd_sc_hd__nor2_1 _18348_ (.A(_10326_),
    .B(_10329_),
    .Y(_10330_));
 sky130_fd_sc_hd__nor2_1 _18349_ (.A(_10325_),
    .B(_10328_),
    .Y(_10331_));
 sky130_fd_sc_hd__or2_1 _18350_ (.A(_10330_),
    .B(_10331_),
    .X(_10332_));
 sky130_fd_sc_hd__xnor2_1 _18351_ (.A(_10252_),
    .B(_10332_),
    .Y(_10333_));
 sky130_fd_sc_hd__a32o_1 _18352_ (.A1(net434),
    .A2(_10248_),
    .A3(_10249_),
    .B1(_10333_),
    .B2(net436),
    .X(_10334_));
 sky130_fd_sc_hd__mux2_1 _18353_ (.A0(\top0.pid_d.out[5] ),
    .A1(_10334_),
    .S(net14),
    .X(_10335_));
 sky130_fd_sc_hd__and2_1 _18354_ (.A(net1018),
    .B(_10335_),
    .X(_10336_));
 sky130_fd_sc_hd__clkbuf_1 _18355_ (.A(_10336_),
    .X(_00250_));
 sky130_fd_sc_hd__inv_2 _18356_ (.A(\top0.pid_d.curr_int[5] ),
    .Y(_10337_));
 sky130_fd_sc_hd__o21ba_1 _18357_ (.A1(_10337_),
    .A2(_10246_),
    .B1_N(\top0.pid_d.out[5] ),
    .X(_10338_));
 sky130_fd_sc_hd__a21o_1 _18358_ (.A1(_10337_),
    .A2(_10246_),
    .B1(_10338_),
    .X(_10339_));
 sky130_fd_sc_hd__xnor2_1 _18359_ (.A(\top0.pid_d.out[6] ),
    .B(\top0.pid_d.curr_int[6] ),
    .Y(_10340_));
 sky130_fd_sc_hd__nand2_1 _18360_ (.A(_10339_),
    .B(_10340_),
    .Y(_10341_));
 sky130_fd_sc_hd__or2_1 _18361_ (.A(_10339_),
    .B(_10340_),
    .X(_10342_));
 sky130_fd_sc_hd__o221a_1 _18362_ (.A1(_10165_),
    .A2(_10251_),
    .B1(_10326_),
    .B2(_10329_),
    .C1(_10250_),
    .X(_10343_));
 sky130_fd_sc_hd__nor2_1 _18363_ (.A(_10331_),
    .B(_10343_),
    .Y(_10344_));
 sky130_fd_sc_hd__a21bo_1 _18364_ (.A1(_10306_),
    .A2(_10316_),
    .B1_N(_10304_),
    .X(_10345_));
 sky130_fd_sc_hd__o21a_1 _18365_ (.A1(_10306_),
    .A2(_10316_),
    .B1(_10345_),
    .X(_10346_));
 sky130_fd_sc_hd__a22o_1 _18366_ (.A1(net396),
    .A2(_09518_),
    .B1(_09399_),
    .B2(_10074_),
    .X(_10347_));
 sky130_fd_sc_hd__a2bb2o_1 _18367_ (.A1_N(_10260_),
    .A2_N(_10265_),
    .B1(_10347_),
    .B2(_10255_),
    .X(_10348_));
 sky130_fd_sc_hd__o21ai_1 _18368_ (.A1(net397),
    .A2(_10203_),
    .B1(_09363_),
    .Y(_10349_));
 sky130_fd_sc_hd__a32o_1 _18369_ (.A1(net390),
    .A2(net364),
    .A3(_10349_),
    .B1(_09429_),
    .B2(_09363_),
    .X(_10350_));
 sky130_fd_sc_hd__nand2_1 _18370_ (.A(net391),
    .B(net317),
    .Y(_10351_));
 sky130_fd_sc_hd__a22o_1 _18371_ (.A1(net319),
    .A2(_10350_),
    .B1(_10351_),
    .B2(_10208_),
    .X(_10352_));
 sky130_fd_sc_hd__nand2_1 _18372_ (.A(net401),
    .B(net312),
    .Y(_10353_));
 sky130_fd_sc_hd__nand2_1 _18373_ (.A(net396),
    .B(net314),
    .Y(_10354_));
 sky130_fd_sc_hd__xor2_1 _18374_ (.A(_10353_),
    .B(_10354_),
    .X(_10355_));
 sky130_fd_sc_hd__nand2_1 _18375_ (.A(net405),
    .B(net310),
    .Y(_10356_));
 sky130_fd_sc_hd__xor2_1 _18376_ (.A(_10355_),
    .B(_10356_),
    .X(_10357_));
 sky130_fd_sc_hd__xnor2_1 _18377_ (.A(_10352_),
    .B(_10357_),
    .Y(_10358_));
 sky130_fd_sc_hd__o21ba_1 _18378_ (.A1(_10293_),
    .A2(_10295_),
    .B1_N(_10291_),
    .X(_10359_));
 sky130_fd_sc_hd__a21o_1 _18379_ (.A1(_10293_),
    .A2(_10295_),
    .B1(_10359_),
    .X(_10360_));
 sky130_fd_sc_hd__nor2_1 _18380_ (.A(_10358_),
    .B(_10360_),
    .Y(_10361_));
 sky130_fd_sc_hd__nand2_1 _18381_ (.A(_10358_),
    .B(_10360_),
    .Y(_10362_));
 sky130_fd_sc_hd__or2b_1 _18382_ (.A(_10361_),
    .B_N(_10362_),
    .X(_10363_));
 sky130_fd_sc_hd__xnor2_1 _18383_ (.A(_10348_),
    .B(_10363_),
    .Y(_10364_));
 sky130_fd_sc_hd__nand2_2 _18384_ (.A(net338),
    .B(net369),
    .Y(_10365_));
 sky130_fd_sc_hd__nand2_1 _18385_ (.A(net331),
    .B(net376),
    .Y(_10366_));
 sky130_fd_sc_hd__nand2_1 _18386_ (.A(net334),
    .B(net373),
    .Y(_10367_));
 sky130_fd_sc_hd__xor2_1 _18387_ (.A(_10366_),
    .B(_10367_),
    .X(_10368_));
 sky130_fd_sc_hd__xnor2_2 _18388_ (.A(_10365_),
    .B(_10368_),
    .Y(_10369_));
 sky130_fd_sc_hd__o21ai_1 _18389_ (.A1(_10278_),
    .A2(_10280_),
    .B1(_10279_),
    .Y(_10370_));
 sky130_fd_sc_hd__a21bo_1 _18390_ (.A1(_10278_),
    .A2(_10280_),
    .B1_N(_10370_),
    .X(_10371_));
 sky130_fd_sc_hd__nand2_1 _18391_ (.A(net1022),
    .B(net378),
    .Y(_10372_));
 sky130_fd_sc_hd__nand2_1 _18392_ (.A(net1023),
    .B(net386),
    .Y(_10373_));
 sky130_fd_sc_hd__nand2_1 _18393_ (.A(net324),
    .B(net381),
    .Y(_10374_));
 sky130_fd_sc_hd__xnor2_1 _18394_ (.A(_10373_),
    .B(_10374_),
    .Y(_10375_));
 sky130_fd_sc_hd__xnor2_1 _18395_ (.A(_10372_),
    .B(_10375_),
    .Y(_10376_));
 sky130_fd_sc_hd__nor2_1 _18396_ (.A(_10371_),
    .B(_10376_),
    .Y(_10377_));
 sky130_fd_sc_hd__nand2_1 _18397_ (.A(_10371_),
    .B(_10376_),
    .Y(_10378_));
 sky130_fd_sc_hd__and2b_1 _18398_ (.A_N(_10377_),
    .B(_10378_),
    .X(_10379_));
 sky130_fd_sc_hd__xnor2_2 _18399_ (.A(_10369_),
    .B(_10379_),
    .Y(_10380_));
 sky130_fd_sc_hd__a21oi_1 _18400_ (.A1(_10275_),
    .A2(_10284_),
    .B1(_10283_),
    .Y(_10381_));
 sky130_fd_sc_hd__o21ai_1 _18401_ (.A1(_10271_),
    .A2(_10273_),
    .B1(_10272_),
    .Y(_10382_));
 sky130_fd_sc_hd__a21boi_1 _18402_ (.A1(_10271_),
    .A2(_10273_),
    .B1_N(_10382_),
    .Y(_10383_));
 sky130_fd_sc_hd__inv_2 _18403_ (.A(net368),
    .Y(_10384_));
 sky130_fd_sc_hd__o21a_1 _18404_ (.A1(net348),
    .A2(_10384_),
    .B1(net344),
    .X(_10385_));
 sky130_fd_sc_hd__a21o_1 _18405_ (.A1(net348),
    .A2(_10384_),
    .B1(_10385_),
    .X(_10386_));
 sky130_fd_sc_hd__or3_1 _18406_ (.A(net341),
    .B(net344),
    .C(net348),
    .X(_10387_));
 sky130_fd_sc_hd__nand2_1 _18407_ (.A(net364),
    .B(_10387_),
    .Y(_10388_));
 sky130_fd_sc_hd__a21oi_1 _18408_ (.A1(net341),
    .A2(_10386_),
    .B1(_10388_),
    .Y(_10389_));
 sky130_fd_sc_hd__xnor2_1 _18409_ (.A(_10383_),
    .B(_10389_),
    .Y(_10390_));
 sky130_fd_sc_hd__and2_1 _18410_ (.A(_10381_),
    .B(_10390_),
    .X(_10391_));
 sky130_fd_sc_hd__or2_1 _18411_ (.A(_10381_),
    .B(_10390_),
    .X(_10392_));
 sky130_fd_sc_hd__or2b_1 _18412_ (.A(_10391_),
    .B_N(_10392_),
    .X(_10393_));
 sky130_fd_sc_hd__xor2_2 _18413_ (.A(_10380_),
    .B(_10393_),
    .X(_10394_));
 sky130_fd_sc_hd__inv_2 _18414_ (.A(_10287_),
    .Y(_10395_));
 sky130_fd_sc_hd__a21o_1 _18415_ (.A1(_10395_),
    .A2(_10297_),
    .B1(_10286_),
    .X(_10396_));
 sky130_fd_sc_hd__o21a_1 _18416_ (.A1(_10395_),
    .A2(_10297_),
    .B1(_10396_),
    .X(_10397_));
 sky130_fd_sc_hd__xnor2_1 _18417_ (.A(_10394_),
    .B(_10397_),
    .Y(_10398_));
 sky130_fd_sc_hd__xnor2_1 _18418_ (.A(_10364_),
    .B(_10398_),
    .Y(_10399_));
 sky130_fd_sc_hd__a21oi_2 _18419_ (.A1(_10270_),
    .A2(_10302_),
    .B1(_10301_),
    .Y(_10400_));
 sky130_fd_sc_hd__o21ba_1 _18420_ (.A1(_10266_),
    .A2(_10268_),
    .B1_N(_10256_),
    .X(_10401_));
 sky130_fd_sc_hd__a21oi_2 _18421_ (.A1(_10266_),
    .A2(_10268_),
    .B1(_10401_),
    .Y(_10402_));
 sky130_fd_sc_hd__and3_1 _18422_ (.A(net406),
    .B(net402),
    .C(_09967_),
    .X(_10403_));
 sky130_fd_sc_hd__xnor2_1 _18423_ (.A(net307),
    .B(_10403_),
    .Y(_10404_));
 sky130_fd_sc_hd__a21oi_1 _18424_ (.A1(net310),
    .A2(_10263_),
    .B1(_10403_),
    .Y(_10405_));
 sky130_fd_sc_hd__mux2_1 _18425_ (.A0(_10404_),
    .A1(_10405_),
    .S(net411),
    .X(_10406_));
 sky130_fd_sc_hd__or3_2 _18426_ (.A(net416),
    .B(_09365_),
    .C(_10228_),
    .X(_10407_));
 sky130_fd_sc_hd__xor2_1 _18427_ (.A(_10406_),
    .B(_10407_),
    .X(_10408_));
 sky130_fd_sc_hd__xnor2_2 _18428_ (.A(_10402_),
    .B(_10408_),
    .Y(_10409_));
 sky130_fd_sc_hd__xnor2_1 _18429_ (.A(_10400_),
    .B(_10409_),
    .Y(_10410_));
 sky130_fd_sc_hd__xnor2_1 _18430_ (.A(_10399_),
    .B(_10410_),
    .Y(_10411_));
 sky130_fd_sc_hd__inv_2 _18431_ (.A(_10314_),
    .Y(_10412_));
 sky130_fd_sc_hd__o21a_1 _18432_ (.A1(_10308_),
    .A2(_10412_),
    .B1(_10229_),
    .X(_10413_));
 sky130_fd_sc_hd__a21oi_1 _18433_ (.A1(_10308_),
    .A2(_10412_),
    .B1(_10413_),
    .Y(_10414_));
 sky130_fd_sc_hd__or2_1 _18434_ (.A(_10411_),
    .B(_10414_),
    .X(_10415_));
 sky130_fd_sc_hd__nand2_1 _18435_ (.A(_10411_),
    .B(_10414_),
    .Y(_10416_));
 sky130_fd_sc_hd__nand2_1 _18436_ (.A(_10415_),
    .B(_10416_),
    .Y(_10417_));
 sky130_fd_sc_hd__xnor2_1 _18437_ (.A(_10346_),
    .B(_10417_),
    .Y(_10418_));
 sky130_fd_sc_hd__nand2_1 _18438_ (.A(_10318_),
    .B(_10322_),
    .Y(_10419_));
 sky130_fd_sc_hd__and3_1 _18439_ (.A(_10323_),
    .B(_10418_),
    .C(_10419_),
    .X(_10420_));
 sky130_fd_sc_hd__a21o_1 _18440_ (.A1(_10323_),
    .A2(_10419_),
    .B1(_10418_),
    .X(_10421_));
 sky130_fd_sc_hd__and2b_1 _18441_ (.A_N(_10420_),
    .B(_10421_),
    .X(_10422_));
 sky130_fd_sc_hd__xnor2_1 _18442_ (.A(_10344_),
    .B(_10422_),
    .Y(_10423_));
 sky130_fd_sc_hd__a32o_1 _18443_ (.A1(net434),
    .A2(_10341_),
    .A3(_10342_),
    .B1(_10423_),
    .B2(net436),
    .X(_10424_));
 sky130_fd_sc_hd__mux2_1 _18444_ (.A0(\top0.pid_d.out[6] ),
    .A1(_10424_),
    .S(net14),
    .X(_10425_));
 sky130_fd_sc_hd__and2_1 _18445_ (.A(_05449_),
    .B(_10425_),
    .X(_10426_));
 sky130_fd_sc_hd__clkbuf_1 _18446_ (.A(_10426_),
    .X(_00251_));
 sky130_fd_sc_hd__inv_2 _18447_ (.A(\top0.pid_d.curr_int[6] ),
    .Y(_10427_));
 sky130_fd_sc_hd__o21ba_1 _18448_ (.A1(_10427_),
    .A2(_10339_),
    .B1_N(\top0.pid_d.out[6] ),
    .X(_10428_));
 sky130_fd_sc_hd__a21o_1 _18449_ (.A1(_10427_),
    .A2(_10339_),
    .B1(_10428_),
    .X(_10429_));
 sky130_fd_sc_hd__xnor2_1 _18450_ (.A(\top0.pid_d.out[7] ),
    .B(\top0.pid_d.curr_int[7] ),
    .Y(_10430_));
 sky130_fd_sc_hd__nand2_1 _18451_ (.A(_10429_),
    .B(_10430_),
    .Y(_10431_));
 sky130_fd_sc_hd__or2_1 _18452_ (.A(_10429_),
    .B(_10430_),
    .X(_10432_));
 sky130_fd_sc_hd__or3_2 _18453_ (.A(_10331_),
    .B(_10343_),
    .C(_10420_),
    .X(_10433_));
 sky130_fd_sc_hd__nand2_1 _18454_ (.A(_10421_),
    .B(_10433_),
    .Y(_10434_));
 sky130_fd_sc_hd__a21o_1 _18455_ (.A1(_10406_),
    .A2(_10407_),
    .B1(_10402_),
    .X(_10435_));
 sky130_fd_sc_hd__o21ai_2 _18456_ (.A1(_10406_),
    .A2(_10407_),
    .B1(_10435_),
    .Y(_10436_));
 sky130_fd_sc_hd__a21o_1 _18457_ (.A1(_10400_),
    .A2(_10409_),
    .B1(_10399_),
    .X(_10437_));
 sky130_fd_sc_hd__o21a_1 _18458_ (.A1(_10400_),
    .A2(_10409_),
    .B1(_10437_),
    .X(_10438_));
 sky130_fd_sc_hd__nor2_1 _18459_ (.A(_10436_),
    .B(_10438_),
    .Y(_10439_));
 sky130_fd_sc_hd__and2_1 _18460_ (.A(_10436_),
    .B(_10438_),
    .X(_10440_));
 sky130_fd_sc_hd__or2_1 _18461_ (.A(_10439_),
    .B(_10440_),
    .X(_10441_));
 sky130_fd_sc_hd__nand2_1 _18462_ (.A(_10346_),
    .B(_10415_),
    .Y(_10442_));
 sky130_fd_sc_hd__and2_2 _18463_ (.A(_10416_),
    .B(_10442_),
    .X(_10443_));
 sky130_fd_sc_hd__a22o_1 _18464_ (.A1(net390),
    .A2(_09518_),
    .B1(_09429_),
    .B2(_10074_),
    .X(_10444_));
 sky130_fd_sc_hd__a2bb2o_1 _18465_ (.A1_N(_10352_),
    .A2_N(_10357_),
    .B1(_10444_),
    .B2(_10255_),
    .X(_10445_));
 sky130_fd_sc_hd__o21ai_1 _18466_ (.A1(net392),
    .A2(_10203_),
    .B1(_09362_),
    .Y(_10446_));
 sky130_fd_sc_hd__a32o_1 _18467_ (.A1(net385),
    .A2(net364),
    .A3(_10446_),
    .B1(_09494_),
    .B2(_09363_),
    .X(_10447_));
 sky130_fd_sc_hd__nand2_1 _18468_ (.A(net385),
    .B(net317),
    .Y(_10448_));
 sky130_fd_sc_hd__a22o_1 _18469_ (.A1(net317),
    .A2(_10447_),
    .B1(_10448_),
    .B2(_10208_),
    .X(_10449_));
 sky130_fd_sc_hd__nand2_1 _18470_ (.A(net396),
    .B(net312),
    .Y(_10450_));
 sky130_fd_sc_hd__nand2_1 _18471_ (.A(net393),
    .B(net315),
    .Y(_10451_));
 sky130_fd_sc_hd__xor2_2 _18472_ (.A(_10450_),
    .B(_10451_),
    .X(_10452_));
 sky130_fd_sc_hd__nand2_1 _18473_ (.A(net401),
    .B(net309),
    .Y(_10453_));
 sky130_fd_sc_hd__xor2_1 _18474_ (.A(_10452_),
    .B(_10453_),
    .X(_10454_));
 sky130_fd_sc_hd__xnor2_1 _18475_ (.A(_10449_),
    .B(_10454_),
    .Y(_10455_));
 sky130_fd_sc_hd__nor2_1 _18476_ (.A(net344),
    .B(net348),
    .Y(_10456_));
 sky130_fd_sc_hd__or3b_1 _18477_ (.A(net369),
    .B(_10456_),
    .C_N(net341),
    .X(_10457_));
 sky130_fd_sc_hd__and2_2 _18478_ (.A(net344),
    .B(net348),
    .X(_10458_));
 sky130_fd_sc_hd__a32o_1 _18479_ (.A1(_10383_),
    .A2(_10387_),
    .A3(_10457_),
    .B1(_10458_),
    .B2(net341),
    .X(_10459_));
 sky130_fd_sc_hd__nand2_1 _18480_ (.A(net364),
    .B(_10459_),
    .Y(_10460_));
 sky130_fd_sc_hd__nor2_1 _18481_ (.A(_10455_),
    .B(_10460_),
    .Y(_10461_));
 sky130_fd_sc_hd__nand2_1 _18482_ (.A(_10455_),
    .B(_10460_),
    .Y(_10462_));
 sky130_fd_sc_hd__and2b_1 _18483_ (.A_N(_10461_),
    .B(_10462_),
    .X(_10463_));
 sky130_fd_sc_hd__xnor2_2 _18484_ (.A(_10445_),
    .B(_10463_),
    .Y(_10464_));
 sky130_fd_sc_hd__nand2_2 _18485_ (.A(net327),
    .B(net376),
    .Y(_10465_));
 sky130_fd_sc_hd__nand2_1 _18486_ (.A(net320),
    .B(net381),
    .Y(_10466_));
 sky130_fd_sc_hd__nand2_1 _18487_ (.A(net323),
    .B(net379),
    .Y(_10467_));
 sky130_fd_sc_hd__xor2_1 _18488_ (.A(_10466_),
    .B(_10467_),
    .X(_10468_));
 sky130_fd_sc_hd__xnor2_2 _18489_ (.A(_10465_),
    .B(_10468_),
    .Y(_10469_));
 sky130_fd_sc_hd__o21ai_1 _18490_ (.A1(_10372_),
    .A2(_10374_),
    .B1(_10373_),
    .Y(_10470_));
 sky130_fd_sc_hd__a21bo_1 _18491_ (.A1(_10372_),
    .A2(_10374_),
    .B1_N(_10470_),
    .X(_10471_));
 sky130_fd_sc_hd__nand2_1 _18492_ (.A(net338),
    .B(net364),
    .Y(_10472_));
 sky130_fd_sc_hd__nand2_1 _18493_ (.A(net331),
    .B(net373),
    .Y(_10473_));
 sky130_fd_sc_hd__nand2_1 _18494_ (.A(net334),
    .B(net369),
    .Y(_10474_));
 sky130_fd_sc_hd__xnor2_1 _18495_ (.A(_10473_),
    .B(_10474_),
    .Y(_10475_));
 sky130_fd_sc_hd__xnor2_1 _18496_ (.A(_10472_),
    .B(_10475_),
    .Y(_10476_));
 sky130_fd_sc_hd__nor2_1 _18497_ (.A(_10471_),
    .B(_10476_),
    .Y(_10477_));
 sky130_fd_sc_hd__nand2_1 _18498_ (.A(_10471_),
    .B(_10476_),
    .Y(_10478_));
 sky130_fd_sc_hd__and2b_1 _18499_ (.A_N(_10477_),
    .B(_10478_),
    .X(_10479_));
 sky130_fd_sc_hd__xnor2_1 _18500_ (.A(_10469_),
    .B(_10479_),
    .Y(_10480_));
 sky130_fd_sc_hd__a21oi_2 _18501_ (.A1(_10369_),
    .A2(_10378_),
    .B1(_10377_),
    .Y(_10481_));
 sky130_fd_sc_hd__o21a_1 _18502_ (.A1(_10365_),
    .A2(_10367_),
    .B1(_10366_),
    .X(_10482_));
 sky130_fd_sc_hd__a21oi_2 _18503_ (.A1(_10365_),
    .A2(_10367_),
    .B1(_10482_),
    .Y(_10483_));
 sky130_fd_sc_hd__a21oi_4 _18504_ (.A1(net341),
    .A2(_10458_),
    .B1(_10388_),
    .Y(_10484_));
 sky130_fd_sc_hd__xnor2_2 _18505_ (.A(_10483_),
    .B(_10484_),
    .Y(_10485_));
 sky130_fd_sc_hd__xor2_1 _18506_ (.A(_10481_),
    .B(_10485_),
    .X(_10486_));
 sky130_fd_sc_hd__xnor2_1 _18507_ (.A(_10480_),
    .B(_10486_),
    .Y(_10487_));
 sky130_fd_sc_hd__a21o_1 _18508_ (.A1(_10380_),
    .A2(_10392_),
    .B1(_10391_),
    .X(_10488_));
 sky130_fd_sc_hd__xor2_1 _18509_ (.A(_10487_),
    .B(_10488_),
    .X(_10489_));
 sky130_fd_sc_hd__xnor2_2 _18510_ (.A(_10464_),
    .B(_10489_),
    .Y(_10490_));
 sky130_fd_sc_hd__a21o_1 _18511_ (.A1(_10394_),
    .A2(_10397_),
    .B1(_10364_),
    .X(_10491_));
 sky130_fd_sc_hd__o21a_1 _18512_ (.A1(_10394_),
    .A2(_10397_),
    .B1(_10491_),
    .X(_10492_));
 sky130_fd_sc_hd__o21ai_2 _18513_ (.A1(_10348_),
    .A2(_10361_),
    .B1(_10362_),
    .Y(_10493_));
 sky130_fd_sc_hd__clkbuf_4 _18514_ (.A(_10103_),
    .X(_10494_));
 sky130_fd_sc_hd__buf_2 _18515_ (.A(_09967_),
    .X(_10495_));
 sky130_fd_sc_hd__and3_1 _18516_ (.A(net401),
    .B(net396),
    .C(_10495_),
    .X(_10496_));
 sky130_fd_sc_hd__xnor2_1 _18517_ (.A(_10494_),
    .B(_10496_),
    .Y(_10497_));
 sky130_fd_sc_hd__a211o_1 _18518_ (.A1(net310),
    .A2(_10355_),
    .B1(_10496_),
    .C1(_09401_),
    .X(_10498_));
 sky130_fd_sc_hd__o21ai_2 _18519_ (.A1(net405),
    .A2(_10497_),
    .B1(_10498_),
    .Y(_10499_));
 sky130_fd_sc_hd__or3_1 _18520_ (.A(net410),
    .B(_09460_),
    .C(_10228_),
    .X(_10500_));
 sky130_fd_sc_hd__xnor2_1 _18521_ (.A(_10499_),
    .B(_10500_),
    .Y(_10501_));
 sky130_fd_sc_hd__xnor2_2 _18522_ (.A(_10493_),
    .B(_10501_),
    .Y(_10502_));
 sky130_fd_sc_hd__xor2_1 _18523_ (.A(_10492_),
    .B(_10502_),
    .X(_10503_));
 sky130_fd_sc_hd__xnor2_2 _18524_ (.A(_10490_),
    .B(_10503_),
    .Y(_10504_));
 sky130_fd_sc_hd__inv_2 _18525_ (.A(_10504_),
    .Y(_10505_));
 sky130_fd_sc_hd__xnor2_1 _18526_ (.A(_10443_),
    .B(_10505_),
    .Y(_10506_));
 sky130_fd_sc_hd__xnor2_1 _18527_ (.A(_10441_),
    .B(_10506_),
    .Y(_10507_));
 sky130_fd_sc_hd__xnor2_1 _18528_ (.A(_10434_),
    .B(_10507_),
    .Y(_10508_));
 sky130_fd_sc_hd__a32o_1 _18529_ (.A1(net434),
    .A2(_10431_),
    .A3(_10432_),
    .B1(_10508_),
    .B2(net436),
    .X(_10509_));
 sky130_fd_sc_hd__mux2_1 _18530_ (.A0(\top0.pid_d.out[7] ),
    .A1(_10509_),
    .S(net14),
    .X(_10510_));
 sky130_fd_sc_hd__and2_1 _18531_ (.A(_05449_),
    .B(_10510_),
    .X(_10511_));
 sky130_fd_sc_hd__clkbuf_1 _18532_ (.A(_10511_),
    .X(_00252_));
 sky130_fd_sc_hd__inv_2 _18533_ (.A(\top0.pid_d.curr_int[7] ),
    .Y(_10512_));
 sky130_fd_sc_hd__o21ba_1 _18534_ (.A1(_10512_),
    .A2(_10429_),
    .B1_N(\top0.pid_d.out[7] ),
    .X(_10513_));
 sky130_fd_sc_hd__a21o_1 _18535_ (.A1(_10512_),
    .A2(_10429_),
    .B1(_10513_),
    .X(_10514_));
 sky130_fd_sc_hd__xnor2_1 _18536_ (.A(\top0.pid_d.out[8] ),
    .B(\top0.pid_d.curr_int[8] ),
    .Y(_10515_));
 sky130_fd_sc_hd__nand2_1 _18537_ (.A(_10514_),
    .B(_10515_),
    .Y(_10516_));
 sky130_fd_sc_hd__or2_1 _18538_ (.A(_10514_),
    .B(_10515_),
    .X(_10517_));
 sky130_fd_sc_hd__a22o_1 _18539_ (.A1(net385),
    .A2(_09518_),
    .B1(_09494_),
    .B2(_10074_),
    .X(_10518_));
 sky130_fd_sc_hd__o2bb2a_2 _18540_ (.A1_N(_10255_),
    .A2_N(_10518_),
    .B1(_10454_),
    .B2(_10449_),
    .X(_10519_));
 sky130_fd_sc_hd__o21ai_1 _18541_ (.A1(net387),
    .A2(_10203_),
    .B1(_09364_),
    .Y(_10520_));
 sky130_fd_sc_hd__a32o_1 _18542_ (.A1(net382),
    .A2(net367),
    .A3(_10520_),
    .B1(_09689_),
    .B2(_09364_),
    .X(_10521_));
 sky130_fd_sc_hd__nand2_1 _18543_ (.A(net382),
    .B(net317),
    .Y(_10522_));
 sky130_fd_sc_hd__a22o_1 _18544_ (.A1(net317),
    .A2(_10521_),
    .B1(_10522_),
    .B2(_10208_),
    .X(_10523_));
 sky130_fd_sc_hd__nand2_1 _18545_ (.A(net390),
    .B(net312),
    .Y(_10524_));
 sky130_fd_sc_hd__nand2_1 _18546_ (.A(net387),
    .B(net314),
    .Y(_10525_));
 sky130_fd_sc_hd__xor2_1 _18547_ (.A(_10524_),
    .B(_10525_),
    .X(_10526_));
 sky130_fd_sc_hd__nand2_1 _18548_ (.A(net396),
    .B(net309),
    .Y(_10527_));
 sky130_fd_sc_hd__xor2_1 _18549_ (.A(_10526_),
    .B(_10527_),
    .X(_10528_));
 sky130_fd_sc_hd__xor2_1 _18550_ (.A(_10523_),
    .B(_10528_),
    .X(_10529_));
 sky130_fd_sc_hd__o21a_1 _18551_ (.A1(_10483_),
    .A2(_10458_),
    .B1(net341),
    .X(_10530_));
 sky130_fd_sc_hd__and2b_1 _18552_ (.A_N(_10456_),
    .B(_10483_),
    .X(_10531_));
 sky130_fd_sc_hd__o21a_1 _18553_ (.A1(_10530_),
    .A2(_10531_),
    .B1(net364),
    .X(_10532_));
 sky130_fd_sc_hd__nor2_1 _18554_ (.A(_10529_),
    .B(_10532_),
    .Y(_10533_));
 sky130_fd_sc_hd__nand2_1 _18555_ (.A(_10529_),
    .B(_10532_),
    .Y(_10534_));
 sky130_fd_sc_hd__or2b_2 _18556_ (.A(_10533_),
    .B_N(_10534_),
    .X(_10535_));
 sky130_fd_sc_hd__xnor2_4 _18557_ (.A(_10519_),
    .B(_10535_),
    .Y(_10536_));
 sky130_fd_sc_hd__nand2_2 _18558_ (.A(net327),
    .B(net373),
    .Y(_10537_));
 sky130_fd_sc_hd__nand2_1 _18559_ (.A(net320),
    .B(net379),
    .Y(_10538_));
 sky130_fd_sc_hd__nand2_1 _18560_ (.A(net323),
    .B(net376),
    .Y(_10539_));
 sky130_fd_sc_hd__xor2_1 _18561_ (.A(_10538_),
    .B(_10539_),
    .X(_10540_));
 sky130_fd_sc_hd__xnor2_2 _18562_ (.A(_10537_),
    .B(_10540_),
    .Y(_10541_));
 sky130_fd_sc_hd__o21a_1 _18563_ (.A1(_10465_),
    .A2(_10467_),
    .B1(_10466_),
    .X(_10542_));
 sky130_fd_sc_hd__a21oi_1 _18564_ (.A1(_10465_),
    .A2(_10467_),
    .B1(_10542_),
    .Y(_10543_));
 sky130_fd_sc_hd__nand2_1 _18565_ (.A(net331),
    .B(net368),
    .Y(_10544_));
 sky130_fd_sc_hd__xor2_4 _18566_ (.A(net334),
    .B(net338),
    .X(_10545_));
 sky130_fd_sc_hd__nand2_1 _18567_ (.A(net362),
    .B(_10545_),
    .Y(_10546_));
 sky130_fd_sc_hd__xor2_2 _18568_ (.A(_10544_),
    .B(_10546_),
    .X(_10547_));
 sky130_fd_sc_hd__xnor2_1 _18569_ (.A(_10543_),
    .B(_10547_),
    .Y(_10548_));
 sky130_fd_sc_hd__xnor2_2 _18570_ (.A(_10541_),
    .B(_10548_),
    .Y(_10549_));
 sky130_fd_sc_hd__a21oi_2 _18571_ (.A1(_10469_),
    .A2(_10478_),
    .B1(_10477_),
    .Y(_10550_));
 sky130_fd_sc_hd__o21a_1 _18572_ (.A1(_10472_),
    .A2(_10474_),
    .B1(_10473_),
    .X(_10551_));
 sky130_fd_sc_hd__a21oi_2 _18573_ (.A1(_10472_),
    .A2(_10474_),
    .B1(_10551_),
    .Y(_10552_));
 sky130_fd_sc_hd__xnor2_2 _18574_ (.A(_10484_),
    .B(_10552_),
    .Y(_10553_));
 sky130_fd_sc_hd__xor2_1 _18575_ (.A(_10550_),
    .B(_10553_),
    .X(_10554_));
 sky130_fd_sc_hd__xnor2_2 _18576_ (.A(_10549_),
    .B(_10554_),
    .Y(_10555_));
 sky130_fd_sc_hd__a21o_1 _18577_ (.A1(_10481_),
    .A2(_10485_),
    .B1(_10480_),
    .X(_10556_));
 sky130_fd_sc_hd__o21a_1 _18578_ (.A1(_10481_),
    .A2(_10485_),
    .B1(_10556_),
    .X(_10557_));
 sky130_fd_sc_hd__xnor2_2 _18579_ (.A(_10555_),
    .B(_10557_),
    .Y(_10558_));
 sky130_fd_sc_hd__xnor2_4 _18580_ (.A(_10536_),
    .B(_10558_),
    .Y(_10559_));
 sky130_fd_sc_hd__o21ba_1 _18581_ (.A1(_10464_),
    .A2(_10488_),
    .B1_N(_10487_),
    .X(_10560_));
 sky130_fd_sc_hd__a21o_1 _18582_ (.A1(_10464_),
    .A2(_10488_),
    .B1(_10560_),
    .X(_10561_));
 sky130_fd_sc_hd__a21oi_2 _18583_ (.A1(_10445_),
    .A2(_10462_),
    .B1(_10461_),
    .Y(_10562_));
 sky130_fd_sc_hd__and3_1 _18584_ (.A(net397),
    .B(net393),
    .C(_09967_),
    .X(_10563_));
 sky130_fd_sc_hd__xnor2_1 _18585_ (.A(_10103_),
    .B(_10563_),
    .Y(_10564_));
 sky130_fd_sc_hd__a211o_1 _18586_ (.A1(net309),
    .A2(_10452_),
    .B1(_10563_),
    .C1(_09353_),
    .X(_10565_));
 sky130_fd_sc_hd__o21ai_2 _18587_ (.A1(net402),
    .A2(_10564_),
    .B1(_10565_),
    .Y(_10566_));
 sky130_fd_sc_hd__or4_2 _18588_ (.A(net406),
    .B(_09353_),
    .C(_09351_),
    .D(_10228_),
    .X(_10567_));
 sky130_fd_sc_hd__xnor2_1 _18589_ (.A(_10566_),
    .B(_10567_),
    .Y(_10568_));
 sky130_fd_sc_hd__xnor2_1 _18590_ (.A(_10562_),
    .B(_10568_),
    .Y(_10569_));
 sky130_fd_sc_hd__and2_1 _18591_ (.A(_10561_),
    .B(_10569_),
    .X(_10570_));
 sky130_fd_sc_hd__or2_1 _18592_ (.A(_10561_),
    .B(_10569_),
    .X(_10571_));
 sky130_fd_sc_hd__and2b_1 _18593_ (.A_N(_10570_),
    .B(_10571_),
    .X(_10572_));
 sky130_fd_sc_hd__xor2_4 _18594_ (.A(_10559_),
    .B(_10572_),
    .X(_10573_));
 sky130_fd_sc_hd__o21ba_1 _18595_ (.A1(_10490_),
    .A2(_10502_),
    .B1_N(_10492_),
    .X(_10574_));
 sky130_fd_sc_hd__a21o_1 _18596_ (.A1(_10490_),
    .A2(_10502_),
    .B1(_10574_),
    .X(_10575_));
 sky130_fd_sc_hd__o21a_1 _18597_ (.A1(_10499_),
    .A2(_10500_),
    .B1(_10493_),
    .X(_10576_));
 sky130_fd_sc_hd__a21o_1 _18598_ (.A1(_10499_),
    .A2(_10500_),
    .B1(_10576_),
    .X(_10577_));
 sky130_fd_sc_hd__xor2_2 _18599_ (.A(_10575_),
    .B(_10577_),
    .X(_10578_));
 sky130_fd_sc_hd__xnor2_4 _18600_ (.A(_10573_),
    .B(_10578_),
    .Y(_10579_));
 sky130_fd_sc_hd__and3_1 _18601_ (.A(_10421_),
    .B(_10433_),
    .C(_10436_),
    .X(_10580_));
 sky130_fd_sc_hd__and2_1 _18602_ (.A(_10438_),
    .B(_10580_),
    .X(_10581_));
 sky130_fd_sc_hd__a21o_1 _18603_ (.A1(_10421_),
    .A2(_10433_),
    .B1(_10436_),
    .X(_10582_));
 sky130_fd_sc_hd__a21o_1 _18604_ (.A1(_10438_),
    .A2(_10582_),
    .B1(_10580_),
    .X(_10583_));
 sky130_fd_sc_hd__a21o_1 _18605_ (.A1(_10505_),
    .A2(_10583_),
    .B1(_10581_),
    .X(_10584_));
 sky130_fd_sc_hd__inv_2 _18606_ (.A(_10443_),
    .Y(_10585_));
 sky130_fd_sc_hd__o21ai_1 _18607_ (.A1(_10438_),
    .A2(_10580_),
    .B1(_10582_),
    .Y(_10586_));
 sky130_fd_sc_hd__a211oi_1 _18608_ (.A1(_10585_),
    .A2(_10505_),
    .B1(_10582_),
    .C1(_10438_),
    .Y(_10587_));
 sky130_fd_sc_hd__a31o_1 _18609_ (.A1(_10443_),
    .A2(_10504_),
    .A3(_10586_),
    .B1(_10587_),
    .X(_10588_));
 sky130_fd_sc_hd__a221o_1 _18610_ (.A1(_10505_),
    .A2(_10581_),
    .B1(_10584_),
    .B2(_10585_),
    .C1(_10588_),
    .X(_10589_));
 sky130_fd_sc_hd__xnor2_1 _18611_ (.A(_10579_),
    .B(_10589_),
    .Y(_10590_));
 sky130_fd_sc_hd__a32o_1 _18612_ (.A1(net432),
    .A2(_10516_),
    .A3(_10517_),
    .B1(_10590_),
    .B2(net436),
    .X(_10591_));
 sky130_fd_sc_hd__mux2_1 _18613_ (.A0(\top0.pid_d.out[8] ),
    .A1(_10591_),
    .S(net14),
    .X(_10592_));
 sky130_fd_sc_hd__and2_1 _18614_ (.A(_05449_),
    .B(_10592_),
    .X(_10593_));
 sky130_fd_sc_hd__clkbuf_1 _18615_ (.A(_10593_),
    .X(_00253_));
 sky130_fd_sc_hd__inv_2 _18616_ (.A(\top0.pid_d.curr_int[8] ),
    .Y(_10594_));
 sky130_fd_sc_hd__o21ba_1 _18617_ (.A1(_10594_),
    .A2(_10514_),
    .B1_N(\top0.pid_d.out[8] ),
    .X(_10595_));
 sky130_fd_sc_hd__a21o_1 _18618_ (.A1(_10594_),
    .A2(_10514_),
    .B1(_10595_),
    .X(_10596_));
 sky130_fd_sc_hd__xnor2_1 _18619_ (.A(\top0.pid_d.out[9] ),
    .B(\top0.pid_d.curr_int[9] ),
    .Y(_10597_));
 sky130_fd_sc_hd__nand2_1 _18620_ (.A(_10596_),
    .B(_10597_),
    .Y(_10598_));
 sky130_fd_sc_hd__or2_1 _18621_ (.A(_10596_),
    .B(_10597_),
    .X(_10599_));
 sky130_fd_sc_hd__o21bai_1 _18622_ (.A1(_10439_),
    .A2(_10504_),
    .B1_N(_10440_),
    .Y(_10600_));
 sky130_fd_sc_hd__o211a_1 _18623_ (.A1(_10579_),
    .A2(_10600_),
    .B1(_10421_),
    .C1(_10507_),
    .X(_10601_));
 sky130_fd_sc_hd__inv_2 _18624_ (.A(_10579_),
    .Y(_10602_));
 sky130_fd_sc_hd__nor2_1 _18625_ (.A(_10440_),
    .B(_10579_),
    .Y(_10603_));
 sky130_fd_sc_hd__o22a_1 _18626_ (.A1(_10439_),
    .A2(_10602_),
    .B1(_10603_),
    .B2(_10504_),
    .X(_10604_));
 sky130_fd_sc_hd__nor2_1 _18627_ (.A(_10443_),
    .B(_10604_),
    .Y(_10605_));
 sky130_fd_sc_hd__a221o_2 _18628_ (.A1(_10579_),
    .A2(_10600_),
    .B1(_10601_),
    .B2(_10433_),
    .C1(_10605_),
    .X(_10606_));
 sky130_fd_sc_hd__o21a_1 _18629_ (.A1(_10573_),
    .A2(_10577_),
    .B1(_10575_),
    .X(_10607_));
 sky130_fd_sc_hd__a21oi_1 _18630_ (.A1(_10573_),
    .A2(_10577_),
    .B1(_10607_),
    .Y(_10608_));
 sky130_fd_sc_hd__a22o_1 _18631_ (.A1(net382),
    .A2(_09518_),
    .B1(_09689_),
    .B2(_10074_),
    .X(_10609_));
 sky130_fd_sc_hd__a2bb2o_2 _18632_ (.A1_N(_10523_),
    .A2_N(_10528_),
    .B1(_10609_),
    .B2(_10255_),
    .X(_10610_));
 sky130_fd_sc_hd__o21ai_1 _18633_ (.A1(net381),
    .A2(_10203_),
    .B1(_09364_),
    .Y(_10611_));
 sky130_fd_sc_hd__nor2_1 _18634_ (.A(_09706_),
    .B(net377),
    .Y(_10612_));
 sky130_fd_sc_hd__a32o_1 _18635_ (.A1(net377),
    .A2(net364),
    .A3(_10611_),
    .B1(_10612_),
    .B2(_09364_),
    .X(_10613_));
 sky130_fd_sc_hd__nand2_1 _18636_ (.A(net377),
    .B(net316),
    .Y(_10614_));
 sky130_fd_sc_hd__a22o_1 _18637_ (.A1(net316),
    .A2(_10613_),
    .B1(_10614_),
    .B2(_10208_),
    .X(_10615_));
 sky130_fd_sc_hd__nand2_1 _18638_ (.A(net381),
    .B(net314),
    .Y(_10616_));
 sky130_fd_sc_hd__nand2_1 _18639_ (.A(net387),
    .B(net311),
    .Y(_10617_));
 sky130_fd_sc_hd__xnor2_1 _18640_ (.A(_10616_),
    .B(_10617_),
    .Y(_10618_));
 sky130_fd_sc_hd__nand2_1 _18641_ (.A(net390),
    .B(net309),
    .Y(_10619_));
 sky130_fd_sc_hd__xnor2_1 _18642_ (.A(_10618_),
    .B(_10619_),
    .Y(_10620_));
 sky130_fd_sc_hd__xnor2_1 _18643_ (.A(_10615_),
    .B(_10620_),
    .Y(_10621_));
 sky130_fd_sc_hd__o21a_1 _18644_ (.A1(_10458_),
    .A2(_10552_),
    .B1(net341),
    .X(_10622_));
 sky130_fd_sc_hd__and2b_1 _18645_ (.A_N(_10456_),
    .B(_10552_),
    .X(_10623_));
 sky130_fd_sc_hd__o21ai_1 _18646_ (.A1(_10622_),
    .A2(_10623_),
    .B1(net364),
    .Y(_10624_));
 sky130_fd_sc_hd__nand2_1 _18647_ (.A(_10621_),
    .B(_10624_),
    .Y(_10625_));
 sky130_fd_sc_hd__inv_2 _18648_ (.A(_10625_),
    .Y(_10626_));
 sky130_fd_sc_hd__nor2_1 _18649_ (.A(_10621_),
    .B(_10624_),
    .Y(_10627_));
 sky130_fd_sc_hd__nor2_1 _18650_ (.A(_10626_),
    .B(_10627_),
    .Y(_10628_));
 sky130_fd_sc_hd__xor2_2 _18651_ (.A(_10610_),
    .B(_10628_),
    .X(_10629_));
 sky130_fd_sc_hd__a21o_1 _18652_ (.A1(_10543_),
    .A2(_10547_),
    .B1(_10541_),
    .X(_10630_));
 sky130_fd_sc_hd__o21a_1 _18653_ (.A1(_10543_),
    .A2(_10547_),
    .B1(_10630_),
    .X(_10631_));
 sky130_fd_sc_hd__xor2_4 _18654_ (.A(net331),
    .B(_10545_),
    .X(_10632_));
 sky130_fd_sc_hd__nand2_4 _18655_ (.A(net362),
    .B(_10632_),
    .Y(_10633_));
 sky130_fd_sc_hd__o21ai_1 _18656_ (.A1(_10537_),
    .A2(_10539_),
    .B1(_10538_),
    .Y(_10634_));
 sky130_fd_sc_hd__a21bo_1 _18657_ (.A1(_10537_),
    .A2(_10539_),
    .B1_N(_10634_),
    .X(_10635_));
 sky130_fd_sc_hd__nand2_1 _18658_ (.A(net327),
    .B(net368),
    .Y(_10636_));
 sky130_fd_sc_hd__nand2_1 _18659_ (.A(net320),
    .B(net376),
    .Y(_10637_));
 sky130_fd_sc_hd__nand2_1 _18660_ (.A(net323),
    .B(net373),
    .Y(_10638_));
 sky130_fd_sc_hd__xnor2_1 _18661_ (.A(_10637_),
    .B(_10638_),
    .Y(_10639_));
 sky130_fd_sc_hd__xnor2_1 _18662_ (.A(_10636_),
    .B(_10639_),
    .Y(_10640_));
 sky130_fd_sc_hd__xnor2_1 _18663_ (.A(_10635_),
    .B(_10640_),
    .Y(_10641_));
 sky130_fd_sc_hd__xnor2_1 _18664_ (.A(_10633_),
    .B(_10641_),
    .Y(_10642_));
 sky130_fd_sc_hd__o211a_1 _18665_ (.A1(net334),
    .A2(net338),
    .B1(net369),
    .C1(net331),
    .X(_10643_));
 sky130_fd_sc_hd__o21a_1 _18666_ (.A1(_09377_),
    .A2(_10643_),
    .B1(net364),
    .X(_10644_));
 sky130_fd_sc_hd__xnor2_1 _18667_ (.A(_10484_),
    .B(_10644_),
    .Y(_10645_));
 sky130_fd_sc_hd__nor2_1 _18668_ (.A(_10642_),
    .B(_10645_),
    .Y(_10646_));
 sky130_fd_sc_hd__nand2_1 _18669_ (.A(_10642_),
    .B(_10645_),
    .Y(_10647_));
 sky130_fd_sc_hd__and2b_1 _18670_ (.A_N(_10646_),
    .B(_10647_),
    .X(_10648_));
 sky130_fd_sc_hd__xnor2_1 _18671_ (.A(_10631_),
    .B(_10648_),
    .Y(_10649_));
 sky130_fd_sc_hd__o21ba_1 _18672_ (.A1(_10550_),
    .A2(_10553_),
    .B1_N(_10549_),
    .X(_10650_));
 sky130_fd_sc_hd__a21o_1 _18673_ (.A1(_10550_),
    .A2(_10553_),
    .B1(_10650_),
    .X(_10651_));
 sky130_fd_sc_hd__nor2_1 _18674_ (.A(_10649_),
    .B(_10651_),
    .Y(_10652_));
 sky130_fd_sc_hd__nand2_1 _18675_ (.A(_10649_),
    .B(_10651_),
    .Y(_10653_));
 sky130_fd_sc_hd__or2b_1 _18676_ (.A(_10652_),
    .B_N(_10653_),
    .X(_10654_));
 sky130_fd_sc_hd__xnor2_2 _18677_ (.A(_10629_),
    .B(_10654_),
    .Y(_10655_));
 sky130_fd_sc_hd__o21a_1 _18678_ (.A1(_10555_),
    .A2(_10557_),
    .B1(_10536_),
    .X(_10656_));
 sky130_fd_sc_hd__a21o_1 _18679_ (.A1(_10555_),
    .A2(_10557_),
    .B1(_10656_),
    .X(_10657_));
 sky130_fd_sc_hd__a21oi_1 _18680_ (.A1(_10519_),
    .A2(_10534_),
    .B1(_10533_),
    .Y(_10658_));
 sky130_fd_sc_hd__and3_1 _18681_ (.A(net390),
    .B(net387),
    .C(_10495_),
    .X(_10659_));
 sky130_fd_sc_hd__xnor2_1 _18682_ (.A(_10494_),
    .B(_10659_),
    .Y(_10660_));
 sky130_fd_sc_hd__a211o_1 _18683_ (.A1(net309),
    .A2(_10526_),
    .B1(_10659_),
    .C1(_09351_),
    .X(_10661_));
 sky130_fd_sc_hd__o21ai_2 _18684_ (.A1(net396),
    .A2(_10660_),
    .B1(_10661_),
    .Y(_10662_));
 sky130_fd_sc_hd__or3_2 _18685_ (.A(net401),
    .B(_09433_),
    .C(_10228_),
    .X(_10663_));
 sky130_fd_sc_hd__xor2_1 _18686_ (.A(_10662_),
    .B(_10663_),
    .X(_10664_));
 sky130_fd_sc_hd__xnor2_1 _18687_ (.A(_10658_),
    .B(_10664_),
    .Y(_10665_));
 sky130_fd_sc_hd__nand2_1 _18688_ (.A(_10657_),
    .B(_10665_),
    .Y(_10666_));
 sky130_fd_sc_hd__inv_2 _18689_ (.A(_10666_),
    .Y(_10667_));
 sky130_fd_sc_hd__nor2_1 _18690_ (.A(_10657_),
    .B(_10665_),
    .Y(_10668_));
 sky130_fd_sc_hd__nor2_1 _18691_ (.A(_10667_),
    .B(_10668_),
    .Y(_10669_));
 sky130_fd_sc_hd__xnor2_2 _18692_ (.A(_10655_),
    .B(_10669_),
    .Y(_10670_));
 sky130_fd_sc_hd__a21o_1 _18693_ (.A1(_10559_),
    .A2(_10571_),
    .B1(_10570_),
    .X(_10671_));
 sky130_fd_sc_hd__o21a_1 _18694_ (.A1(_10566_),
    .A2(_10567_),
    .B1(_10562_),
    .X(_10672_));
 sky130_fd_sc_hd__a21o_1 _18695_ (.A1(_10566_),
    .A2(_10567_),
    .B1(_10672_),
    .X(_10673_));
 sky130_fd_sc_hd__xor2_1 _18696_ (.A(_10671_),
    .B(_10673_),
    .X(_10674_));
 sky130_fd_sc_hd__xnor2_1 _18697_ (.A(_10670_),
    .B(_10674_),
    .Y(_10675_));
 sky130_fd_sc_hd__nor2_1 _18698_ (.A(_10608_),
    .B(_10675_),
    .Y(_10676_));
 sky130_fd_sc_hd__and2_1 _18699_ (.A(_10608_),
    .B(_10675_),
    .X(_10677_));
 sky130_fd_sc_hd__or2_1 _18700_ (.A(_10676_),
    .B(_10677_),
    .X(_10678_));
 sky130_fd_sc_hd__xnor2_2 _18701_ (.A(_10606_),
    .B(_10678_),
    .Y(_10679_));
 sky130_fd_sc_hd__a32o_1 _18702_ (.A1(net432),
    .A2(_10598_),
    .A3(_10599_),
    .B1(_10679_),
    .B2(net437),
    .X(_10680_));
 sky130_fd_sc_hd__mux2_1 _18703_ (.A0(\top0.pid_d.out[9] ),
    .A1(_10680_),
    .S(_07141_),
    .X(_10681_));
 sky130_fd_sc_hd__and2_1 _18704_ (.A(_05449_),
    .B(_10681_),
    .X(_10682_));
 sky130_fd_sc_hd__clkbuf_1 _18705_ (.A(_10682_),
    .X(_00254_));
 sky130_fd_sc_hd__inv_2 _18706_ (.A(_10676_),
    .Y(_10683_));
 sky130_fd_sc_hd__o21ai_2 _18707_ (.A1(_10606_),
    .A2(_10677_),
    .B1(_10683_),
    .Y(_10684_));
 sky130_fd_sc_hd__o21a_1 _18708_ (.A1(_10671_),
    .A2(_10673_),
    .B1(_10670_),
    .X(_10685_));
 sky130_fd_sc_hd__a21o_1 _18709_ (.A1(_10671_),
    .A2(_10673_),
    .B1(_10685_),
    .X(_10686_));
 sky130_fd_sc_hd__a22o_1 _18710_ (.A1(net377),
    .A2(_09518_),
    .B1(_10074_),
    .B2(_10612_),
    .X(_10687_));
 sky130_fd_sc_hd__o2bb2a_2 _18711_ (.A1_N(_10255_),
    .A2_N(_10687_),
    .B1(_10615_),
    .B2(_10620_),
    .X(_10688_));
 sky130_fd_sc_hd__o21ai_1 _18712_ (.A1(net377),
    .A2(_10203_),
    .B1(_09364_),
    .Y(_10689_));
 sky130_fd_sc_hd__inv_2 _18713_ (.A(net374),
    .Y(_10690_));
 sky130_fd_sc_hd__and3_1 _18714_ (.A(net377),
    .B(_10690_),
    .C(_09364_),
    .X(_10691_));
 sky130_fd_sc_hd__a31o_1 _18715_ (.A1(net374),
    .A2(net365),
    .A3(_10689_),
    .B1(_10691_),
    .X(_10692_));
 sky130_fd_sc_hd__nand2_1 _18716_ (.A(net376),
    .B(net316),
    .Y(_10693_));
 sky130_fd_sc_hd__a22o_1 _18717_ (.A1(net317),
    .A2(_10692_),
    .B1(_10693_),
    .B2(_10208_),
    .X(_10694_));
 sky130_fd_sc_hd__nand2_1 _18718_ (.A(net381),
    .B(net312),
    .Y(_10695_));
 sky130_fd_sc_hd__nand2_1 _18719_ (.A(net377),
    .B(net314),
    .Y(_10696_));
 sky130_fd_sc_hd__xor2_1 _18720_ (.A(_10695_),
    .B(_10696_),
    .X(_10697_));
 sky130_fd_sc_hd__nand2_1 _18721_ (.A(net389),
    .B(net308),
    .Y(_10698_));
 sky130_fd_sc_hd__xor2_1 _18722_ (.A(_10697_),
    .B(_10698_),
    .X(_10699_));
 sky130_fd_sc_hd__xor2_1 _18723_ (.A(_10694_),
    .B(_10699_),
    .X(_10700_));
 sky130_fd_sc_hd__o21a_1 _18724_ (.A1(_10458_),
    .A2(_10644_),
    .B1(net341),
    .X(_10701_));
 sky130_fd_sc_hd__and2b_1 _18725_ (.A_N(_10456_),
    .B(_10644_),
    .X(_10702_));
 sky130_fd_sc_hd__o21a_1 _18726_ (.A1(_10701_),
    .A2(_10702_),
    .B1(net362),
    .X(_10703_));
 sky130_fd_sc_hd__nor2_1 _18727_ (.A(_10700_),
    .B(_10703_),
    .Y(_10704_));
 sky130_fd_sc_hd__nand2_1 _18728_ (.A(_10700_),
    .B(_10703_),
    .Y(_10705_));
 sky130_fd_sc_hd__and2b_1 _18729_ (.A_N(_10704_),
    .B(_10705_),
    .X(_10706_));
 sky130_fd_sc_hd__xnor2_4 _18730_ (.A(_10688_),
    .B(_10706_),
    .Y(_10707_));
 sky130_fd_sc_hd__o21ai_1 _18731_ (.A1(_10636_),
    .A2(_10638_),
    .B1(_10637_),
    .Y(_10708_));
 sky130_fd_sc_hd__a21bo_1 _18732_ (.A1(_10636_),
    .A2(_10638_),
    .B1_N(_10708_),
    .X(_10709_));
 sky130_fd_sc_hd__nand2_1 _18733_ (.A(net327),
    .B(net362),
    .Y(_10710_));
 sky130_fd_sc_hd__nand2_1 _18734_ (.A(net320),
    .B(net373),
    .Y(_10711_));
 sky130_fd_sc_hd__nand2_2 _18735_ (.A(net323),
    .B(net368),
    .Y(_10712_));
 sky130_fd_sc_hd__xnor2_1 _18736_ (.A(_10711_),
    .B(_10712_),
    .Y(_10713_));
 sky130_fd_sc_hd__xnor2_2 _18737_ (.A(_10710_),
    .B(_10713_),
    .Y(_10714_));
 sky130_fd_sc_hd__xnor2_1 _18738_ (.A(_10709_),
    .B(_10714_),
    .Y(_10715_));
 sky130_fd_sc_hd__xnor2_2 _18739_ (.A(_10633_),
    .B(_10715_),
    .Y(_10716_));
 sky130_fd_sc_hd__o21a_1 _18740_ (.A1(_10635_),
    .A2(_10640_),
    .B1(_10633_),
    .X(_10717_));
 sky130_fd_sc_hd__a21o_1 _18741_ (.A1(_10635_),
    .A2(_10640_),
    .B1(_10717_),
    .X(_10718_));
 sky130_fd_sc_hd__o21a_1 _18742_ (.A1(net334),
    .A2(net338),
    .B1(net331),
    .X(_10719_));
 sky130_fd_sc_hd__or2_1 _18743_ (.A(_09377_),
    .B(_10719_),
    .X(_10720_));
 sky130_fd_sc_hd__nand2_1 _18744_ (.A(net362),
    .B(_10720_),
    .Y(_10721_));
 sky130_fd_sc_hd__xor2_2 _18745_ (.A(_10484_),
    .B(_10721_),
    .X(_10722_));
 sky130_fd_sc_hd__inv_2 _18746_ (.A(_10722_),
    .Y(_10723_));
 sky130_fd_sc_hd__xnor2_1 _18747_ (.A(_10718_),
    .B(_10723_),
    .Y(_10724_));
 sky130_fd_sc_hd__xnor2_1 _18748_ (.A(_10716_),
    .B(_10724_),
    .Y(_10725_));
 sky130_fd_sc_hd__o21a_1 _18749_ (.A1(_10631_),
    .A2(_10646_),
    .B1(_10647_),
    .X(_10726_));
 sky130_fd_sc_hd__or2_1 _18750_ (.A(_10725_),
    .B(_10726_),
    .X(_10727_));
 sky130_fd_sc_hd__inv_2 _18751_ (.A(_10727_),
    .Y(_10728_));
 sky130_fd_sc_hd__and2_1 _18752_ (.A(_10725_),
    .B(_10726_),
    .X(_10729_));
 sky130_fd_sc_hd__nor2_2 _18753_ (.A(_10728_),
    .B(_10729_),
    .Y(_10730_));
 sky130_fd_sc_hd__xnor2_4 _18754_ (.A(_10707_),
    .B(_10730_),
    .Y(_10731_));
 sky130_fd_sc_hd__a21oi_1 _18755_ (.A1(_10629_),
    .A2(_10653_),
    .B1(_10652_),
    .Y(_10732_));
 sky130_fd_sc_hd__a21oi_2 _18756_ (.A1(_10610_),
    .A2(_10625_),
    .B1(_10627_),
    .Y(_10733_));
 sky130_fd_sc_hd__a21oi_1 _18757_ (.A1(_09771_),
    .A2(_10495_),
    .B1(_10494_),
    .Y(_10734_));
 sky130_fd_sc_hd__and3_1 _18758_ (.A(_10494_),
    .B(_09771_),
    .C(_10495_),
    .X(_10735_));
 sky130_fd_sc_hd__nand2_1 _18759_ (.A(_10616_),
    .B(_10617_),
    .Y(_10736_));
 sky130_fd_sc_hd__a221o_1 _18760_ (.A1(_09771_),
    .A2(_10495_),
    .B1(_10736_),
    .B2(net309),
    .C1(_09493_),
    .X(_10737_));
 sky130_fd_sc_hd__o31ai_4 _18761_ (.A1(net390),
    .A2(_10734_),
    .A3(_10735_),
    .B1(_10737_),
    .Y(_10738_));
 sky130_fd_sc_hd__or3_2 _18762_ (.A(_09688_),
    .B(_09459_),
    .C(_10228_),
    .X(_10739_));
 sky130_fd_sc_hd__xnor2_1 _18763_ (.A(_10738_),
    .B(_10739_),
    .Y(_10740_));
 sky130_fd_sc_hd__xnor2_2 _18764_ (.A(_10733_),
    .B(_10740_),
    .Y(_10741_));
 sky130_fd_sc_hd__xor2_1 _18765_ (.A(_10732_),
    .B(_10741_),
    .X(_10742_));
 sky130_fd_sc_hd__xnor2_2 _18766_ (.A(_10731_),
    .B(_10742_),
    .Y(_10743_));
 sky130_fd_sc_hd__o21ai_1 _18767_ (.A1(_10655_),
    .A2(_10668_),
    .B1(_10666_),
    .Y(_10744_));
 sky130_fd_sc_hd__o21ba_1 _18768_ (.A1(_10662_),
    .A2(_10663_),
    .B1_N(_10658_),
    .X(_10745_));
 sky130_fd_sc_hd__a21oi_1 _18769_ (.A1(_10662_),
    .A2(_10663_),
    .B1(_10745_),
    .Y(_10746_));
 sky130_fd_sc_hd__and2b_1 _18770_ (.A_N(_10744_),
    .B(_10746_),
    .X(_10747_));
 sky130_fd_sc_hd__or2b_1 _18771_ (.A(_10746_),
    .B_N(_10744_),
    .X(_10748_));
 sky130_fd_sc_hd__and2b_1 _18772_ (.A_N(_10747_),
    .B(_10748_),
    .X(_10749_));
 sky130_fd_sc_hd__xnor2_1 _18773_ (.A(_10743_),
    .B(_10749_),
    .Y(_10750_));
 sky130_fd_sc_hd__and2_1 _18774_ (.A(_10686_),
    .B(_10750_),
    .X(_10751_));
 sky130_fd_sc_hd__or2_1 _18775_ (.A(_10686_),
    .B(_10750_),
    .X(_10752_));
 sky130_fd_sc_hd__or2b_1 _18776_ (.A(_10751_),
    .B_N(_10752_),
    .X(_10753_));
 sky130_fd_sc_hd__xor2_2 _18777_ (.A(_10684_),
    .B(_10753_),
    .X(_10754_));
 sky130_fd_sc_hd__nor2_1 _18778_ (.A(\top0.pid_d.out[10] ),
    .B(_07137_),
    .Y(_10755_));
 sky130_fd_sc_hd__inv_2 _18779_ (.A(\top0.pid_d.curr_int[9] ),
    .Y(_10756_));
 sky130_fd_sc_hd__o21ba_1 _18780_ (.A1(_10756_),
    .A2(_10596_),
    .B1_N(\top0.pid_d.out[9] ),
    .X(_10757_));
 sky130_fd_sc_hd__a21o_1 _18781_ (.A1(_10756_),
    .A2(_10596_),
    .B1(_10757_),
    .X(_10758_));
 sky130_fd_sc_hd__xnor2_1 _18782_ (.A(\top0.pid_d.curr_int[10] ),
    .B(_10758_),
    .Y(_10759_));
 sky130_fd_sc_hd__mux2_1 _18783_ (.A0(\top0.pid_d.out[10] ),
    .A1(_10755_),
    .S(_10759_),
    .X(_10760_));
 sky130_fd_sc_hd__a22o_1 _18784_ (.A1(\top0.pid_d.out[10] ),
    .A2(_07137_),
    .B1(_10760_),
    .B2(net432),
    .X(_10761_));
 sky130_fd_sc_hd__a31o_1 _18785_ (.A1(net437),
    .A2(_09339_),
    .A3(_10754_),
    .B1(_10761_),
    .X(_10762_));
 sky130_fd_sc_hd__and2_1 _18786_ (.A(_05449_),
    .B(_10762_),
    .X(_10763_));
 sky130_fd_sc_hd__clkbuf_1 _18787_ (.A(_10763_),
    .X(_00255_));
 sky130_fd_sc_hd__a21oi_1 _18788_ (.A1(_10684_),
    .A2(_10752_),
    .B1(_10751_),
    .Y(_10764_));
 sky130_fd_sc_hd__a21o_1 _18789_ (.A1(_10731_),
    .A2(_10741_),
    .B1(_10732_),
    .X(_10765_));
 sky130_fd_sc_hd__o21ai_4 _18790_ (.A1(_10731_),
    .A2(_10741_),
    .B1(_10765_),
    .Y(_10766_));
 sky130_fd_sc_hd__nor2_1 _18791_ (.A(_09356_),
    .B(_09758_),
    .Y(_10767_));
 sky130_fd_sc_hd__a31o_1 _18792_ (.A1(net377),
    .A2(_10690_),
    .A3(_10074_),
    .B1(_10767_),
    .X(_10768_));
 sky130_fd_sc_hd__o2bb2a_2 _18793_ (.A1_N(_10255_),
    .A2_N(_10768_),
    .B1(_10699_),
    .B2(_10694_),
    .X(_10769_));
 sky130_fd_sc_hd__o21a_1 _18794_ (.A1(_10458_),
    .A2(_10720_),
    .B1(net341),
    .X(_10770_));
 sky130_fd_sc_hd__and2b_1 _18795_ (.A_N(_10456_),
    .B(_10720_),
    .X(_10771_));
 sky130_fd_sc_hd__o21ai_4 _18796_ (.A1(_10770_),
    .A2(_10771_),
    .B1(net362),
    .Y(_10772_));
 sky130_fd_sc_hd__nand2_1 _18797_ (.A(net377),
    .B(net311),
    .Y(_10773_));
 sky130_fd_sc_hd__nand2_1 _18798_ (.A(net374),
    .B(net314),
    .Y(_10774_));
 sky130_fd_sc_hd__xor2_2 _18799_ (.A(_10773_),
    .B(_10774_),
    .X(_10775_));
 sky130_fd_sc_hd__nand2_1 _18800_ (.A(net383),
    .B(net309),
    .Y(_10776_));
 sky130_fd_sc_hd__xor2_2 _18801_ (.A(_10775_),
    .B(_10776_),
    .X(_10777_));
 sky130_fd_sc_hd__nand2_1 _18802_ (.A(net371),
    .B(net318),
    .Y(_10778_));
 sky130_fd_sc_hd__a21oi_1 _18803_ (.A1(net374),
    .A2(_09395_),
    .B1(_09356_),
    .Y(_10779_));
 sky130_fd_sc_hd__a21o_1 _18804_ (.A1(_10690_),
    .A2(net360),
    .B1(_10779_),
    .X(_10780_));
 sky130_fd_sc_hd__nor2_1 _18805_ (.A(_10690_),
    .B(net371),
    .Y(_10781_));
 sky130_fd_sc_hd__a32o_1 _18806_ (.A1(net371),
    .A2(net366),
    .A3(_10780_),
    .B1(_10781_),
    .B2(_09364_),
    .X(_10782_));
 sky130_fd_sc_hd__a22o_1 _18807_ (.A1(_10208_),
    .A2(_10778_),
    .B1(_10782_),
    .B2(net316),
    .X(_10783_));
 sky130_fd_sc_hd__xor2_2 _18808_ (.A(_10777_),
    .B(_10783_),
    .X(_10784_));
 sky130_fd_sc_hd__xnor2_2 _18809_ (.A(_10772_),
    .B(_10784_),
    .Y(_10785_));
 sky130_fd_sc_hd__xnor2_4 _18810_ (.A(_10769_),
    .B(_10785_),
    .Y(_10786_));
 sky130_fd_sc_hd__inv_2 _18811_ (.A(_10786_),
    .Y(_10787_));
 sky130_fd_sc_hd__nor3_1 _18812_ (.A(_10718_),
    .B(_10716_),
    .C(_10723_),
    .Y(_10788_));
 sky130_fd_sc_hd__a31o_1 _18813_ (.A1(_10718_),
    .A2(_10716_),
    .A3(_10723_),
    .B1(_10788_),
    .X(_10789_));
 sky130_fd_sc_hd__inv_2 _18814_ (.A(net373),
    .Y(_10790_));
 sky130_fd_sc_hd__a21o_1 _18815_ (.A1(_10790_),
    .A2(net368),
    .B1(net327),
    .X(_10791_));
 sky130_fd_sc_hd__o21ai_1 _18816_ (.A1(net368),
    .A2(_10711_),
    .B1(_10791_),
    .Y(_10792_));
 sky130_fd_sc_hd__and2_1 _18817_ (.A(net327),
    .B(_10790_),
    .X(_10793_));
 sky130_fd_sc_hd__nor2_1 _18818_ (.A(net323),
    .B(net368),
    .Y(_10794_));
 sky130_fd_sc_hd__or2b_1 _18819_ (.A(net323),
    .B_N(net327),
    .X(_10795_));
 sky130_fd_sc_hd__a21oi_1 _18820_ (.A1(_10712_),
    .A2(_10795_),
    .B1(net320),
    .Y(_10796_));
 sky130_fd_sc_hd__a221o_1 _18821_ (.A1(net323),
    .A2(_10792_),
    .B1(_10793_),
    .B2(_10794_),
    .C1(_10796_),
    .X(_10797_));
 sky130_fd_sc_hd__nand2_1 _18822_ (.A(net320),
    .B(net368),
    .Y(_10798_));
 sky130_fd_sc_hd__o22a_1 _18823_ (.A1(net373),
    .A2(net362),
    .B1(_10793_),
    .B2(net323),
    .X(_10799_));
 sky130_fd_sc_hd__o2bb2a_1 _18824_ (.A1_N(net362),
    .A2_N(_10797_),
    .B1(_10798_),
    .B2(_10799_),
    .X(_10800_));
 sky130_fd_sc_hd__xnor2_1 _18825_ (.A(_10633_),
    .B(_10800_),
    .Y(_10801_));
 sky130_fd_sc_hd__o21a_1 _18826_ (.A1(_10709_),
    .A2(_10714_),
    .B1(_10633_),
    .X(_10802_));
 sky130_fd_sc_hd__a21o_1 _18827_ (.A1(_10709_),
    .A2(_10714_),
    .B1(_10802_),
    .X(_10803_));
 sky130_fd_sc_hd__nand2_1 _18828_ (.A(_10801_),
    .B(_10803_),
    .Y(_10804_));
 sky130_fd_sc_hd__or2_1 _18829_ (.A(_10801_),
    .B(_10803_),
    .X(_10805_));
 sky130_fd_sc_hd__nand2_1 _18830_ (.A(_10804_),
    .B(_10805_),
    .Y(_10806_));
 sky130_fd_sc_hd__xnor2_1 _18831_ (.A(_10789_),
    .B(_10806_),
    .Y(_10807_));
 sky130_fd_sc_hd__xnor2_1 _18832_ (.A(_10787_),
    .B(_10807_),
    .Y(_10808_));
 sky130_fd_sc_hd__a21o_1 _18833_ (.A1(_10688_),
    .A2(_10705_),
    .B1(_10704_),
    .X(_10809_));
 sky130_fd_sc_hd__and3_1 _18834_ (.A(net383),
    .B(net379),
    .C(_10495_),
    .X(_10810_));
 sky130_fd_sc_hd__xnor2_1 _18835_ (.A(_10494_),
    .B(_10810_),
    .Y(_10811_));
 sky130_fd_sc_hd__a211o_1 _18836_ (.A1(net308),
    .A2(_10697_),
    .B1(_10810_),
    .C1(_09688_),
    .X(_10812_));
 sky130_fd_sc_hd__o21ai_2 _18837_ (.A1(net387),
    .A2(_10811_),
    .B1(_10812_),
    .Y(_10813_));
 sky130_fd_sc_hd__or3_2 _18838_ (.A(net391),
    .B(_09692_),
    .C(_10228_),
    .X(_10814_));
 sky130_fd_sc_hd__xor2_1 _18839_ (.A(_10813_),
    .B(_10814_),
    .X(_10815_));
 sky130_fd_sc_hd__xnor2_1 _18840_ (.A(_10809_),
    .B(_10815_),
    .Y(_10816_));
 sky130_fd_sc_hd__o21a_1 _18841_ (.A1(_10707_),
    .A2(_10729_),
    .B1(_10727_),
    .X(_10817_));
 sky130_fd_sc_hd__nor2_1 _18842_ (.A(_10816_),
    .B(_10817_),
    .Y(_10818_));
 sky130_fd_sc_hd__and2_1 _18843_ (.A(_10816_),
    .B(_10817_),
    .X(_10819_));
 sky130_fd_sc_hd__nor2_1 _18844_ (.A(_10818_),
    .B(_10819_),
    .Y(_10820_));
 sky130_fd_sc_hd__xnor2_1 _18845_ (.A(_10808_),
    .B(_10820_),
    .Y(_10821_));
 sky130_fd_sc_hd__a21o_1 _18846_ (.A1(_10738_),
    .A2(_10739_),
    .B1(_10733_),
    .X(_10822_));
 sky130_fd_sc_hd__or2_1 _18847_ (.A(_10738_),
    .B(_10739_),
    .X(_10823_));
 sky130_fd_sc_hd__nand3_2 _18848_ (.A(_10821_),
    .B(_10822_),
    .C(_10823_),
    .Y(_10824_));
 sky130_fd_sc_hd__inv_2 _18849_ (.A(_10824_),
    .Y(_10825_));
 sky130_fd_sc_hd__a21oi_2 _18850_ (.A1(_10822_),
    .A2(_10823_),
    .B1(_10821_),
    .Y(_10826_));
 sky130_fd_sc_hd__nor2_2 _18851_ (.A(_10825_),
    .B(_10826_),
    .Y(_10827_));
 sky130_fd_sc_hd__xnor2_4 _18852_ (.A(_10766_),
    .B(_10827_),
    .Y(_10828_));
 sky130_fd_sc_hd__o21ai_4 _18853_ (.A1(_10743_),
    .A2(_10747_),
    .B1(_10748_),
    .Y(_10829_));
 sky130_fd_sc_hd__xnor2_1 _18854_ (.A(_10828_),
    .B(_10829_),
    .Y(_10830_));
 sky130_fd_sc_hd__xnor2_1 _18855_ (.A(_10764_),
    .B(_10830_),
    .Y(_10831_));
 sky130_fd_sc_hd__and3_1 _18856_ (.A(net435),
    .B(_09339_),
    .C(_10831_),
    .X(_10832_));
 sky130_fd_sc_hd__nor2_1 _18857_ (.A(\top0.pid_d.out[11] ),
    .B(_07138_),
    .Y(_10833_));
 sky130_fd_sc_hd__inv_2 _18858_ (.A(\top0.pid_d.curr_int[10] ),
    .Y(_10834_));
 sky130_fd_sc_hd__o21ba_1 _18859_ (.A1(_10834_),
    .A2(_10758_),
    .B1_N(\top0.pid_d.out[10] ),
    .X(_10835_));
 sky130_fd_sc_hd__a21o_1 _18860_ (.A1(_10834_),
    .A2(_10758_),
    .B1(_10835_),
    .X(_10836_));
 sky130_fd_sc_hd__xnor2_1 _18861_ (.A(\top0.pid_d.curr_int[11] ),
    .B(_10836_),
    .Y(_10837_));
 sky130_fd_sc_hd__mux2_1 _18862_ (.A0(\top0.pid_d.out[11] ),
    .A1(_10833_),
    .S(_10837_),
    .X(_10838_));
 sky130_fd_sc_hd__a22o_1 _18863_ (.A1(\top0.pid_d.out[11] ),
    .A2(_07138_),
    .B1(_10838_),
    .B2(net432),
    .X(_10839_));
 sky130_fd_sc_hd__o21a_1 _18864_ (.A1(_10832_),
    .A2(_10839_),
    .B1(_07710_),
    .X(_00256_));
 sky130_fd_sc_hd__a21oi_1 _18865_ (.A1(_10606_),
    .A2(_10683_),
    .B1(_10677_),
    .Y(_10840_));
 sky130_fd_sc_hd__o21ai_1 _18866_ (.A1(_10751_),
    .A2(_10840_),
    .B1(_10752_),
    .Y(_10841_));
 sky130_fd_sc_hd__o22a_1 _18867_ (.A1(_10718_),
    .A2(_10716_),
    .B1(_10787_),
    .B2(_10806_),
    .X(_10842_));
 sky130_fd_sc_hd__a21oi_1 _18868_ (.A1(_10787_),
    .A2(_10806_),
    .B1(_10842_),
    .Y(_10843_));
 sky130_fd_sc_hd__nand2_1 _18869_ (.A(_10718_),
    .B(_10716_),
    .Y(_10844_));
 sky130_fd_sc_hd__clkbuf_4 _18870_ (.A(_10722_),
    .X(_10845_));
 sky130_fd_sc_hd__a211o_1 _18871_ (.A1(_10786_),
    .A2(_10844_),
    .B1(_10806_),
    .C1(_10845_),
    .X(_10846_));
 sky130_fd_sc_hd__o221ai_4 _18872_ (.A1(_10723_),
    .A2(_10843_),
    .B1(_10844_),
    .B2(_10786_),
    .C1(_10846_),
    .Y(_10847_));
 sky130_fd_sc_hd__inv_2 _18873_ (.A(_10772_),
    .Y(_10848_));
 sky130_fd_sc_hd__o21ba_1 _18874_ (.A1(_10848_),
    .A2(_10784_),
    .B1_N(_10769_),
    .X(_10849_));
 sky130_fd_sc_hd__a21o_1 _18875_ (.A1(_10848_),
    .A2(_10784_),
    .B1(_10849_),
    .X(_10850_));
 sky130_fd_sc_hd__and3_1 _18876_ (.A(net380),
    .B(net374),
    .C(_10495_),
    .X(_10851_));
 sky130_fd_sc_hd__xnor2_1 _18877_ (.A(_10494_),
    .B(_10851_),
    .Y(_10852_));
 sky130_fd_sc_hd__a211o_1 _18878_ (.A1(net308),
    .A2(_10775_),
    .B1(_10851_),
    .C1(_09706_),
    .X(_10853_));
 sky130_fd_sc_hd__o21ai_2 _18879_ (.A1(net383),
    .A2(_10852_),
    .B1(_10853_),
    .Y(_10854_));
 sky130_fd_sc_hd__or3b_2 _18880_ (.A(net389),
    .B(_10494_),
    .C_N(_10810_),
    .X(_10855_));
 sky130_fd_sc_hd__xnor2_1 _18881_ (.A(_10854_),
    .B(_10855_),
    .Y(_10856_));
 sky130_fd_sc_hd__xnor2_1 _18882_ (.A(_10850_),
    .B(_10856_),
    .Y(_10857_));
 sky130_fd_sc_hd__nand2_1 _18883_ (.A(_09395_),
    .B(_10781_),
    .Y(_10858_));
 sky130_fd_sc_hd__a21oi_1 _18884_ (.A1(_09863_),
    .A2(_10858_),
    .B1(_09356_),
    .Y(_10859_));
 sky130_fd_sc_hd__a31o_1 _18885_ (.A1(_09356_),
    .A2(net360),
    .A3(_10781_),
    .B1(_10859_),
    .X(_10860_));
 sky130_fd_sc_hd__a2bb2o_2 _18886_ (.A1_N(_10777_),
    .A2_N(_10783_),
    .B1(_10860_),
    .B2(_10255_),
    .X(_10861_));
 sky130_fd_sc_hd__a21o_1 _18887_ (.A1(_09395_),
    .A2(_10778_),
    .B1(_09356_),
    .X(_10862_));
 sky130_fd_sc_hd__o21ai_1 _18888_ (.A1(_09395_),
    .A2(_10778_),
    .B1(_10862_),
    .Y(_10863_));
 sky130_fd_sc_hd__nand2_1 _18889_ (.A(net365),
    .B(_10863_),
    .Y(_10864_));
 sky130_fd_sc_hd__nand2_1 _18890_ (.A(net371),
    .B(net314),
    .Y(_10865_));
 sky130_fd_sc_hd__nand2_1 _18891_ (.A(net374),
    .B(net312),
    .Y(_10866_));
 sky130_fd_sc_hd__xor2_1 _18892_ (.A(_10865_),
    .B(_10866_),
    .X(_10867_));
 sky130_fd_sc_hd__nand2_1 _18893_ (.A(net380),
    .B(net308),
    .Y(_10868_));
 sky130_fd_sc_hd__xnor2_2 _18894_ (.A(_10867_),
    .B(_10868_),
    .Y(_10869_));
 sky130_fd_sc_hd__nand2_1 _18895_ (.A(net318),
    .B(net370),
    .Y(_10870_));
 sky130_fd_sc_hd__xor2_2 _18896_ (.A(_10075_),
    .B(_10870_),
    .X(_10871_));
 sky130_fd_sc_hd__xor2_1 _18897_ (.A(_10869_),
    .B(_10871_),
    .X(_10872_));
 sky130_fd_sc_hd__xnor2_2 _18898_ (.A(_10864_),
    .B(_10872_),
    .Y(_10873_));
 sky130_fd_sc_hd__xnor2_2 _18899_ (.A(_10772_),
    .B(_10873_),
    .Y(_10874_));
 sky130_fd_sc_hd__xnor2_4 _18900_ (.A(_10861_),
    .B(_10874_),
    .Y(_10875_));
 sky130_fd_sc_hd__o21a_1 _18901_ (.A1(net324),
    .A2(net327),
    .B1(_10384_),
    .X(_10876_));
 sky130_fd_sc_hd__a21o_1 _18902_ (.A1(net323),
    .A2(net327),
    .B1(_10876_),
    .X(_10877_));
 sky130_fd_sc_hd__or3_1 _18903_ (.A(net320),
    .B(net324),
    .C(net327),
    .X(_10878_));
 sky130_fd_sc_hd__nand2_1 _18904_ (.A(net363),
    .B(_10878_),
    .Y(_10879_));
 sky130_fd_sc_hd__a21o_1 _18905_ (.A1(net320),
    .A2(_10877_),
    .B1(_10879_),
    .X(_10880_));
 sky130_fd_sc_hd__nor3_1 _18906_ (.A(_10790_),
    .B(net362),
    .C(_10712_),
    .Y(_10881_));
 sky130_fd_sc_hd__or3_1 _18907_ (.A(net323),
    .B(_10790_),
    .C(net368),
    .X(_10882_));
 sky130_fd_sc_hd__a21oi_1 _18908_ (.A1(_10712_),
    .A2(_10882_),
    .B1(_10710_),
    .Y(_10883_));
 sky130_fd_sc_hd__o21ai_1 _18909_ (.A1(_10881_),
    .A2(_10883_),
    .B1(net320),
    .Y(_10884_));
 sky130_fd_sc_hd__nand2_1 _18910_ (.A(_10800_),
    .B(_10884_),
    .Y(_10885_));
 sky130_fd_sc_hd__mux2_1 _18911_ (.A0(_10885_),
    .A1(_10884_),
    .S(_10633_),
    .X(_10886_));
 sky130_fd_sc_hd__xnor2_1 _18912_ (.A(_10880_),
    .B(_10886_),
    .Y(_10887_));
 sky130_fd_sc_hd__mux2_1 _18913_ (.A0(_10804_),
    .A1(_10805_),
    .S(_10722_),
    .X(_10888_));
 sky130_fd_sc_hd__xnor2_1 _18914_ (.A(_10887_),
    .B(_10888_),
    .Y(_10889_));
 sky130_fd_sc_hd__xnor2_2 _18915_ (.A(_10875_),
    .B(_10889_),
    .Y(_10890_));
 sky130_fd_sc_hd__xor2_1 _18916_ (.A(_10857_),
    .B(_10890_),
    .X(_10891_));
 sky130_fd_sc_hd__xnor2_1 _18917_ (.A(_10847_),
    .B(_10891_),
    .Y(_10892_));
 sky130_fd_sc_hd__o21a_1 _18918_ (.A1(_10813_),
    .A2(_10814_),
    .B1(_10809_),
    .X(_10893_));
 sky130_fd_sc_hd__a21oi_1 _18919_ (.A1(_10813_),
    .A2(_10814_),
    .B1(_10893_),
    .Y(_10894_));
 sky130_fd_sc_hd__inv_2 _18920_ (.A(_10818_),
    .Y(_10895_));
 sky130_fd_sc_hd__a21o_1 _18921_ (.A1(_10808_),
    .A2(_10895_),
    .B1(_10819_),
    .X(_10896_));
 sky130_fd_sc_hd__nor2_1 _18922_ (.A(_10894_),
    .B(_10896_),
    .Y(_10897_));
 sky130_fd_sc_hd__nand2_1 _18923_ (.A(_10894_),
    .B(_10896_),
    .Y(_10898_));
 sky130_fd_sc_hd__and2b_1 _18924_ (.A_N(_10897_),
    .B(_10898_),
    .X(_10899_));
 sky130_fd_sc_hd__xnor2_1 _18925_ (.A(_10892_),
    .B(_10899_),
    .Y(_10900_));
 sky130_fd_sc_hd__inv_2 _18926_ (.A(_10900_),
    .Y(_10901_));
 sky130_fd_sc_hd__o21ai_1 _18927_ (.A1(_10766_),
    .A2(_10826_),
    .B1(_10824_),
    .Y(_10902_));
 sky130_fd_sc_hd__nor2_1 _18928_ (.A(_10901_),
    .B(_10902_),
    .Y(_10903_));
 sky130_fd_sc_hd__and2_1 _18929_ (.A(_10901_),
    .B(_10902_),
    .X(_10904_));
 sky130_fd_sc_hd__or2_2 _18930_ (.A(_10903_),
    .B(_10904_),
    .X(_10905_));
 sky130_fd_sc_hd__nand2_1 _18931_ (.A(_10828_),
    .B(_10829_),
    .Y(_10906_));
 sky130_fd_sc_hd__nor2_1 _18932_ (.A(_10828_),
    .B(_10829_),
    .Y(_10907_));
 sky130_fd_sc_hd__nor3_1 _18933_ (.A(_10841_),
    .B(_10905_),
    .C(_10907_),
    .Y(_10908_));
 sky130_fd_sc_hd__a31o_1 _18934_ (.A1(_10841_),
    .A2(_10905_),
    .A3(_10906_),
    .B1(_10908_),
    .X(_10909_));
 sky130_fd_sc_hd__and2_1 _18935_ (.A(\top0.pid_d.out[12] ),
    .B(\top0.pid_d.curr_int[12] ),
    .X(_10910_));
 sky130_fd_sc_hd__or2_1 _18936_ (.A(\top0.pid_d.out[12] ),
    .B(\top0.pid_d.curr_int[12] ),
    .X(_10911_));
 sky130_fd_sc_hd__or2b_1 _18937_ (.A(_10910_),
    .B_N(_10911_),
    .X(_10912_));
 sky130_fd_sc_hd__nor2_1 _18938_ (.A(\top0.pid_d.out[11] ),
    .B(\top0.pid_d.curr_int[11] ),
    .Y(_10913_));
 sky130_fd_sc_hd__nand2_1 _18939_ (.A(\top0.pid_d.out[11] ),
    .B(\top0.pid_d.curr_int[11] ),
    .Y(_10914_));
 sky130_fd_sc_hd__o21ai_2 _18940_ (.A1(_10836_),
    .A2(_10913_),
    .B1(_10914_),
    .Y(_10915_));
 sky130_fd_sc_hd__xnor2_1 _18941_ (.A(_10912_),
    .B(_10915_),
    .Y(_10916_));
 sky130_fd_sc_hd__and3_1 _18942_ (.A(net435),
    .B(_10828_),
    .C(_10829_),
    .X(_10917_));
 sky130_fd_sc_hd__nor3b_1 _18943_ (.A(_10828_),
    .B(_10829_),
    .C_N(net435),
    .Y(_10918_));
 sky130_fd_sc_hd__mux2_1 _18944_ (.A0(_10917_),
    .A1(_10918_),
    .S(_10905_),
    .X(_10919_));
 sky130_fd_sc_hd__a221o_1 _18945_ (.A1(net436),
    .A2(_10909_),
    .B1(_10916_),
    .B2(net432),
    .C1(_10919_),
    .X(_10920_));
 sky130_fd_sc_hd__mux2_1 _18946_ (.A0(\top0.pid_d.out[12] ),
    .A1(_10920_),
    .S(_07141_),
    .X(_10921_));
 sky130_fd_sc_hd__and2_1 _18947_ (.A(_05449_),
    .B(_10921_),
    .X(_10922_));
 sky130_fd_sc_hd__clkbuf_1 _18948_ (.A(_10922_),
    .X(_00257_));
 sky130_fd_sc_hd__or2b_1 _18949_ (.A(_10829_),
    .B_N(_10841_),
    .X(_10923_));
 sky130_fd_sc_hd__o211a_1 _18950_ (.A1(_10751_),
    .A2(_10840_),
    .B1(_10829_),
    .C1(_10752_),
    .X(_10924_));
 sky130_fd_sc_hd__or2_1 _18951_ (.A(_10828_),
    .B(_10924_),
    .X(_10925_));
 sky130_fd_sc_hd__a21o_1 _18952_ (.A1(_10923_),
    .A2(_10925_),
    .B1(_10904_),
    .X(_10926_));
 sky130_fd_sc_hd__and2b_1 _18953_ (.A_N(_10903_),
    .B(_10926_),
    .X(_10927_));
 sky130_fd_sc_hd__and2b_1 _18954_ (.A_N(_10857_),
    .B(_10890_),
    .X(_10928_));
 sky130_fd_sc_hd__or2b_1 _18955_ (.A(_10890_),
    .B_N(_10857_),
    .X(_10929_));
 sky130_fd_sc_hd__o21ai_2 _18956_ (.A1(_10847_),
    .A2(_10928_),
    .B1(_10929_),
    .Y(_10930_));
 sky130_fd_sc_hd__xor2_1 _18957_ (.A(_10880_),
    .B(_10886_),
    .X(_10931_));
 sky130_fd_sc_hd__a21bo_1 _18958_ (.A1(_10875_),
    .A2(_10931_),
    .B1_N(_10804_),
    .X(_10932_));
 sky130_fd_sc_hd__o21a_1 _18959_ (.A1(_10875_),
    .A2(_10931_),
    .B1(_10932_),
    .X(_10933_));
 sky130_fd_sc_hd__a211o_1 _18960_ (.A1(_10805_),
    .A2(_10875_),
    .B1(_10887_),
    .C1(_10723_),
    .X(_10934_));
 sky130_fd_sc_hd__o221a_2 _18961_ (.A1(_10805_),
    .A2(_10875_),
    .B1(_10933_),
    .B2(_10845_),
    .C1(_10934_),
    .X(_10935_));
 sky130_fd_sc_hd__a21o_1 _18962_ (.A1(_10880_),
    .A2(_10884_),
    .B1(_10845_),
    .X(_10936_));
 sky130_fd_sc_hd__nand2_1 _18963_ (.A(_10633_),
    .B(_10936_),
    .Y(_10937_));
 sky130_fd_sc_hd__a21o_1 _18964_ (.A1(_10880_),
    .A2(_10885_),
    .B1(_10723_),
    .X(_10938_));
 sky130_fd_sc_hd__o211a_1 _18965_ (.A1(_10880_),
    .A2(_10886_),
    .B1(_10937_),
    .C1(_10938_),
    .X(_10939_));
 sky130_fd_sc_hd__o211a_1 _18966_ (.A1(_09965_),
    .A2(_10384_),
    .B1(net311),
    .C1(net373),
    .X(_10940_));
 sky130_fd_sc_hd__a211o_1 _18967_ (.A1(net373),
    .A2(net311),
    .B1(_10384_),
    .C1(_09965_),
    .X(_10941_));
 sky130_fd_sc_hd__or2b_1 _18968_ (.A(_10940_),
    .B_N(_10941_),
    .X(_10942_));
 sky130_fd_sc_hd__nand2_1 _18969_ (.A(net376),
    .B(net308),
    .Y(_10943_));
 sky130_fd_sc_hd__xor2_2 _18970_ (.A(_10942_),
    .B(_10943_),
    .X(_10944_));
 sky130_fd_sc_hd__a21oi_1 _18971_ (.A1(_09395_),
    .A2(net368),
    .B1(_09356_),
    .Y(_10945_));
 sky130_fd_sc_hd__a21o_1 _18972_ (.A1(net360),
    .A2(_10384_),
    .B1(_10945_),
    .X(_10946_));
 sky130_fd_sc_hd__or2_1 _18973_ (.A(net360),
    .B(net316),
    .X(_10947_));
 sky130_fd_sc_hd__o21ai_1 _18974_ (.A1(net356),
    .A2(_10947_),
    .B1(net363),
    .Y(_10948_));
 sky130_fd_sc_hd__a21oi_1 _18975_ (.A1(net316),
    .A2(_10946_),
    .B1(_10948_),
    .Y(_10949_));
 sky130_fd_sc_hd__xnor2_2 _18976_ (.A(_10944_),
    .B(_10949_),
    .Y(_10950_));
 sky130_fd_sc_hd__a22o_1 _18977_ (.A1(net365),
    .A2(_10863_),
    .B1(_10869_),
    .B2(_10871_),
    .X(_10951_));
 sky130_fd_sc_hd__o21a_1 _18978_ (.A1(_10869_),
    .A2(_10871_),
    .B1(_10951_),
    .X(_10952_));
 sky130_fd_sc_hd__xnor2_1 _18979_ (.A(_10848_),
    .B(_10952_),
    .Y(_10953_));
 sky130_fd_sc_hd__xnor2_2 _18980_ (.A(_10950_),
    .B(_10953_),
    .Y(_10954_));
 sky130_fd_sc_hd__o21ai_2 _18981_ (.A1(_10632_),
    .A2(_10878_),
    .B1(net363),
    .Y(_10955_));
 sky130_fd_sc_hd__and2_1 _18982_ (.A(net320),
    .B(_10632_),
    .X(_10956_));
 sky130_fd_sc_hd__and3_1 _18983_ (.A(net363),
    .B(_10877_),
    .C(_10956_),
    .X(_10957_));
 sky130_fd_sc_hd__nor2_1 _18984_ (.A(_10955_),
    .B(_10957_),
    .Y(_10958_));
 sky130_fd_sc_hd__xnor2_1 _18985_ (.A(_10845_),
    .B(_10958_),
    .Y(_10959_));
 sky130_fd_sc_hd__xnor2_1 _18986_ (.A(_10954_),
    .B(_10959_),
    .Y(_10960_));
 sky130_fd_sc_hd__xnor2_1 _18987_ (.A(_10939_),
    .B(_10960_),
    .Y(_10961_));
 sky130_fd_sc_hd__a21o_1 _18988_ (.A1(_10861_),
    .A2(_10873_),
    .B1(_10848_),
    .X(_10962_));
 sky130_fd_sc_hd__o21a_1 _18989_ (.A1(_10861_),
    .A2(_10873_),
    .B1(_10962_),
    .X(_10963_));
 sky130_fd_sc_hd__and3_1 _18990_ (.A(net374),
    .B(net371),
    .C(_10495_),
    .X(_10964_));
 sky130_fd_sc_hd__xnor2_1 _18991_ (.A(net307),
    .B(_10964_),
    .Y(_10965_));
 sky130_fd_sc_hd__nand2_1 _18992_ (.A(_10865_),
    .B(_10866_),
    .Y(_10966_));
 sky130_fd_sc_hd__a21oi_1 _18993_ (.A1(net309),
    .A2(_10966_),
    .B1(_10964_),
    .Y(_10967_));
 sky130_fd_sc_hd__mux2_1 _18994_ (.A0(_10965_),
    .A1(_10967_),
    .S(net380),
    .X(_10968_));
 sky130_fd_sc_hd__or3b_2 _18995_ (.A(net383),
    .B(_10494_),
    .C_N(_10851_),
    .X(_10969_));
 sky130_fd_sc_hd__xnor2_1 _18996_ (.A(_10968_),
    .B(_10969_),
    .Y(_10970_));
 sky130_fd_sc_hd__xnor2_1 _18997_ (.A(_10963_),
    .B(_10970_),
    .Y(_10971_));
 sky130_fd_sc_hd__nand2_1 _18998_ (.A(_10961_),
    .B(_10971_),
    .Y(_10972_));
 sky130_fd_sc_hd__nor2_1 _18999_ (.A(_10961_),
    .B(_10971_),
    .Y(_10973_));
 sky130_fd_sc_hd__inv_2 _19000_ (.A(_10973_),
    .Y(_10974_));
 sky130_fd_sc_hd__nand2_1 _19001_ (.A(_10972_),
    .B(_10974_),
    .Y(_10975_));
 sky130_fd_sc_hd__xnor2_1 _19002_ (.A(_10935_),
    .B(_10975_),
    .Y(_10976_));
 sky130_fd_sc_hd__a21bo_1 _19003_ (.A1(_10854_),
    .A2(_10855_),
    .B1_N(_10850_),
    .X(_10977_));
 sky130_fd_sc_hd__o21a_1 _19004_ (.A1(_10854_),
    .A2(_10855_),
    .B1(_10977_),
    .X(_10978_));
 sky130_fd_sc_hd__nor2_1 _19005_ (.A(_10976_),
    .B(_10978_),
    .Y(_10979_));
 sky130_fd_sc_hd__nand2_1 _19006_ (.A(_10976_),
    .B(_10978_),
    .Y(_10980_));
 sky130_fd_sc_hd__or2b_1 _19007_ (.A(_10979_),
    .B_N(_10980_),
    .X(_10981_));
 sky130_fd_sc_hd__xnor2_1 _19008_ (.A(_10930_),
    .B(_10981_),
    .Y(_10982_));
 sky130_fd_sc_hd__a21o_1 _19009_ (.A1(_10892_),
    .A2(_10898_),
    .B1(_10897_),
    .X(_10983_));
 sky130_fd_sc_hd__xnor2_1 _19010_ (.A(_10982_),
    .B(_10983_),
    .Y(_10984_));
 sky130_fd_sc_hd__xnor2_1 _19011_ (.A(_10927_),
    .B(_10984_),
    .Y(_10985_));
 sky130_fd_sc_hd__a21o_1 _19012_ (.A1(_10911_),
    .A2(_10915_),
    .B1(_10910_),
    .X(_10986_));
 sky130_fd_sc_hd__xnor2_1 _19013_ (.A(\top0.pid_d.out[13] ),
    .B(\top0.pid_d.curr_int[13] ),
    .Y(_10987_));
 sky130_fd_sc_hd__xnor2_1 _19014_ (.A(_10986_),
    .B(_10987_),
    .Y(_10988_));
 sky130_fd_sc_hd__a221o_1 _19015_ (.A1(net435),
    .A2(_10985_),
    .B1(_10988_),
    .B2(net432),
    .C1(_07138_),
    .X(_10989_));
 sky130_fd_sc_hd__o211a_1 _19016_ (.A1(\top0.pid_d.out[13] ),
    .A2(_09339_),
    .B1(_10989_),
    .C1(_10067_),
    .X(_00258_));
 sky130_fd_sc_hd__inv_2 _19017_ (.A(_10983_),
    .Y(_10990_));
 sky130_fd_sc_hd__a21oi_1 _19018_ (.A1(_10982_),
    .A2(_10990_),
    .B1(_10903_),
    .Y(_10991_));
 sky130_fd_sc_hd__a2bb2o_1 _19019_ (.A1_N(_10982_),
    .A2_N(_10990_),
    .B1(_10991_),
    .B2(_10926_),
    .X(_10992_));
 sky130_fd_sc_hd__o21ai_2 _19020_ (.A1(_10930_),
    .A2(_10979_),
    .B1(_10980_),
    .Y(_10993_));
 sky130_fd_sc_hd__a21oi_2 _19021_ (.A1(_10935_),
    .A2(_10972_),
    .B1(_10973_),
    .Y(_10994_));
 sky130_fd_sc_hd__a21bo_1 _19022_ (.A1(_10968_),
    .A2(_10969_),
    .B1_N(_10963_),
    .X(_10995_));
 sky130_fd_sc_hd__o21ai_2 _19023_ (.A1(_10968_),
    .A2(_10969_),
    .B1(_10995_),
    .Y(_10996_));
 sky130_fd_sc_hd__a21o_1 _19024_ (.A1(_10845_),
    .A2(_10958_),
    .B1(_10939_),
    .X(_10997_));
 sky130_fd_sc_hd__a21oi_1 _19025_ (.A1(_10954_),
    .A2(_10955_),
    .B1(_10957_),
    .Y(_10998_));
 sky130_fd_sc_hd__o2bb2a_1 _19026_ (.A1_N(_10954_),
    .A2_N(_10997_),
    .B1(_10998_),
    .B2(_10845_),
    .X(_10999_));
 sky130_fd_sc_hd__and2b_1 _19027_ (.A_N(_10944_),
    .B(_10947_),
    .X(_11000_));
 sky130_fd_sc_hd__nand3_1 _19028_ (.A(net316),
    .B(_10384_),
    .C(_10074_),
    .Y(_11001_));
 sky130_fd_sc_hd__a21bo_1 _19029_ (.A1(net360),
    .A2(net316),
    .B1_N(_10944_),
    .X(_11002_));
 sky130_fd_sc_hd__o2111a_2 _19030_ (.A1(net356),
    .A2(_11000_),
    .B1(_11001_),
    .C1(_11002_),
    .D1(net363),
    .X(_11003_));
 sky130_fd_sc_hd__nand2_1 _19031_ (.A(net314),
    .B(net365),
    .Y(_11004_));
 sky130_fd_sc_hd__and3_1 _19032_ (.A(net371),
    .B(net308),
    .C(_11004_),
    .X(_11005_));
 sky130_fd_sc_hd__a21oi_1 _19033_ (.A1(net371),
    .A2(net308),
    .B1(_11004_),
    .Y(_11006_));
 sky130_fd_sc_hd__a2bb2o_1 _19034_ (.A1_N(_11005_),
    .A2_N(_11006_),
    .B1(net311),
    .B2(net370),
    .X(_11007_));
 sky130_fd_sc_hd__o41a_2 _19035_ (.A1(_09966_),
    .A2(_10384_),
    .A3(_11005_),
    .A4(_11006_),
    .B1(_11007_),
    .X(_11008_));
 sky130_fd_sc_hd__a31o_1 _19036_ (.A1(net356),
    .A2(net360),
    .A3(net316),
    .B1(_10948_),
    .X(_11009_));
 sky130_fd_sc_hd__xor2_2 _19037_ (.A(_11008_),
    .B(_11009_),
    .X(_11010_));
 sky130_fd_sc_hd__xnor2_2 _19038_ (.A(_10772_),
    .B(_11010_),
    .Y(_11011_));
 sky130_fd_sc_hd__xnor2_4 _19039_ (.A(_11003_),
    .B(_11011_),
    .Y(_11012_));
 sky130_fd_sc_hd__mux2_2 _19040_ (.A0(_10957_),
    .A1(_10955_),
    .S(_10845_),
    .X(_11013_));
 sky130_fd_sc_hd__xnor2_4 _19041_ (.A(_11012_),
    .B(_11013_),
    .Y(_11014_));
 sky130_fd_sc_hd__o21a_1 _19042_ (.A1(_10950_),
    .A2(_10952_),
    .B1(_10848_),
    .X(_11015_));
 sky130_fd_sc_hd__a21o_1 _19043_ (.A1(_10950_),
    .A2(_10952_),
    .B1(_11015_),
    .X(_11016_));
 sky130_fd_sc_hd__or3b_2 _19044_ (.A(net377),
    .B(_10494_),
    .C_N(_10964_),
    .X(_11017_));
 sky130_fd_sc_hd__and3_1 _19045_ (.A(net371),
    .B(net370),
    .C(_10495_),
    .X(_11018_));
 sky130_fd_sc_hd__xnor2_1 _19046_ (.A(_10494_),
    .B(_11018_),
    .Y(_11019_));
 sky130_fd_sc_hd__a211o_1 _19047_ (.A1(net309),
    .A2(_10942_),
    .B1(_11018_),
    .C1(_10690_),
    .X(_11020_));
 sky130_fd_sc_hd__o21ai_2 _19048_ (.A1(net374),
    .A2(_11019_),
    .B1(_11020_),
    .Y(_11021_));
 sky130_fd_sc_hd__xnor2_1 _19049_ (.A(_11017_),
    .B(_11021_),
    .Y(_11022_));
 sky130_fd_sc_hd__xnor2_1 _19050_ (.A(_11016_),
    .B(_11022_),
    .Y(_11023_));
 sky130_fd_sc_hd__xnor2_1 _19051_ (.A(_11014_),
    .B(_11023_),
    .Y(_11024_));
 sky130_fd_sc_hd__xnor2_2 _19052_ (.A(_10999_),
    .B(_11024_),
    .Y(_11025_));
 sky130_fd_sc_hd__xor2_1 _19053_ (.A(_10996_),
    .B(_11025_),
    .X(_11026_));
 sky130_fd_sc_hd__xnor2_2 _19054_ (.A(_10994_),
    .B(_11026_),
    .Y(_11027_));
 sky130_fd_sc_hd__nor2_1 _19055_ (.A(_10993_),
    .B(_11027_),
    .Y(_11028_));
 sky130_fd_sc_hd__and2_1 _19056_ (.A(_10993_),
    .B(_11027_),
    .X(_11029_));
 sky130_fd_sc_hd__nor2_1 _19057_ (.A(_11028_),
    .B(_11029_),
    .Y(_11030_));
 sky130_fd_sc_hd__xnor2_1 _19058_ (.A(_10992_),
    .B(_11030_),
    .Y(_11031_));
 sky130_fd_sc_hd__a221o_1 _19059_ (.A1(\top0.pid_d.out[13] ),
    .A2(\top0.pid_d.curr_int[13] ),
    .B1(_10911_),
    .B2(_10915_),
    .C1(_10910_),
    .X(_11032_));
 sky130_fd_sc_hd__o21ai_2 _19060_ (.A1(\top0.pid_d.out[13] ),
    .A2(\top0.pid_d.curr_int[13] ),
    .B1(_11032_),
    .Y(_11033_));
 sky130_fd_sc_hd__xor2_1 _19061_ (.A(\top0.pid_d.out[14] ),
    .B(\top0.pid_d.curr_int[14] ),
    .X(_11034_));
 sky130_fd_sc_hd__xnor2_1 _19062_ (.A(_11033_),
    .B(_11034_),
    .Y(_11035_));
 sky130_fd_sc_hd__a221o_1 _19063_ (.A1(net435),
    .A2(_11031_),
    .B1(_11035_),
    .B2(net432),
    .C1(_07138_),
    .X(_11036_));
 sky130_fd_sc_hd__o211a_1 _19064_ (.A1(\top0.pid_d.out[14] ),
    .A2(_09339_),
    .B1(_11036_),
    .C1(_10067_),
    .X(_00259_));
 sky130_fd_sc_hd__inv_2 _19065_ (.A(_10992_),
    .Y(_11037_));
 sky130_fd_sc_hd__nor2_1 _19066_ (.A(_11017_),
    .B(_11021_),
    .Y(_11038_));
 sky130_fd_sc_hd__nand2_1 _19067_ (.A(_11016_),
    .B(_11038_),
    .Y(_11039_));
 sky130_fd_sc_hd__nand2_1 _19068_ (.A(_11017_),
    .B(_11021_),
    .Y(_11040_));
 sky130_fd_sc_hd__or3b_1 _19069_ (.A(_11016_),
    .B(_11040_),
    .C_N(_11014_),
    .X(_11041_));
 sky130_fd_sc_hd__o21ai_1 _19070_ (.A1(_11016_),
    .A2(_11038_),
    .B1(_11040_),
    .Y(_11042_));
 sky130_fd_sc_hd__o21a_1 _19071_ (.A1(_11014_),
    .A2(_11042_),
    .B1(_11039_),
    .X(_11043_));
 sky130_fd_sc_hd__o2bb2a_1 _19072_ (.A1_N(_11042_),
    .A2_N(_11014_),
    .B1(_11016_),
    .B2(_11040_),
    .X(_11044_));
 sky130_fd_sc_hd__mux2_1 _19073_ (.A0(_11043_),
    .A1(_11044_),
    .S(_10999_),
    .X(_11045_));
 sky130_fd_sc_hd__o211ai_4 _19074_ (.A1(_11014_),
    .A2(_11039_),
    .B1(_11041_),
    .C1(_11045_),
    .Y(_11046_));
 sky130_fd_sc_hd__and4_1 _19075_ (.A(net324),
    .B(net1022),
    .C(net362),
    .D(_10956_),
    .X(_11047_));
 sky130_fd_sc_hd__nor2_1 _19076_ (.A(_10957_),
    .B(_11012_),
    .Y(_11048_));
 sky130_fd_sc_hd__o21ai_1 _19077_ (.A1(_10955_),
    .A2(_11012_),
    .B1(_10845_),
    .Y(_11049_));
 sky130_fd_sc_hd__o31a_1 _19078_ (.A1(_10845_),
    .A2(_11047_),
    .A3(_11048_),
    .B1(_11049_),
    .X(_11050_));
 sky130_fd_sc_hd__a31o_1 _19079_ (.A1(_10690_),
    .A2(net370),
    .A3(_10495_),
    .B1(_10790_),
    .X(_11051_));
 sky130_fd_sc_hd__nand2_1 _19080_ (.A(net307),
    .B(_11051_),
    .Y(_11052_));
 sky130_fd_sc_hd__nand2_1 _19081_ (.A(net370),
    .B(net308),
    .Y(_11053_));
 sky130_fd_sc_hd__o32a_1 _19082_ (.A1(net311),
    .A2(net370),
    .A3(_11004_),
    .B1(_11053_),
    .B2(net365),
    .X(_11054_));
 sky130_fd_sc_hd__a211o_1 _19083_ (.A1(_10790_),
    .A2(net314),
    .B1(net311),
    .C1(_11053_),
    .X(_11055_));
 sky130_fd_sc_hd__a21o_1 _19084_ (.A1(_10384_),
    .A2(net308),
    .B1(_09965_),
    .X(_11056_));
 sky130_fd_sc_hd__a22o_1 _19085_ (.A1(net371),
    .A2(_11056_),
    .B1(_11053_),
    .B2(_09965_),
    .X(_11057_));
 sky130_fd_sc_hd__a211o_1 _19086_ (.A1(net311),
    .A2(_10384_),
    .B1(net308),
    .C1(_09965_),
    .X(_11058_));
 sky130_fd_sc_hd__a21bo_1 _19087_ (.A1(net311),
    .A2(_11057_),
    .B1_N(_11058_),
    .X(_11059_));
 sky130_fd_sc_hd__nand2_1 _19088_ (.A(net365),
    .B(_11059_),
    .Y(_11060_));
 sky130_fd_sc_hd__o211a_1 _19089_ (.A1(net371),
    .A2(_11054_),
    .B1(_11055_),
    .C1(_11060_),
    .X(_11061_));
 sky130_fd_sc_hd__xor2_1 _19090_ (.A(_11052_),
    .B(_11061_),
    .X(_11062_));
 sky130_fd_sc_hd__a21o_1 _19091_ (.A1(net360),
    .A2(net316),
    .B1(_11008_),
    .X(_11063_));
 sky130_fd_sc_hd__a22o_1 _19092_ (.A1(_10947_),
    .A2(_11008_),
    .B1(_11063_),
    .B2(net356),
    .X(_11064_));
 sky130_fd_sc_hd__nand2_1 _19093_ (.A(net363),
    .B(_11064_),
    .Y(_11065_));
 sky130_fd_sc_hd__mux2_1 _19094_ (.A0(_11047_),
    .A1(_10955_),
    .S(_10845_),
    .X(_11066_));
 sky130_fd_sc_hd__xnor2_1 _19095_ (.A(_11065_),
    .B(_11066_),
    .Y(_11067_));
 sky130_fd_sc_hd__xnor2_1 _19096_ (.A(_11062_),
    .B(_11067_),
    .Y(_11068_));
 sky130_fd_sc_hd__nand2_1 _19097_ (.A(_11003_),
    .B(_11010_),
    .Y(_11069_));
 sky130_fd_sc_hd__or3_1 _19098_ (.A(_10772_),
    .B(_11003_),
    .C(_11010_),
    .X(_11070_));
 sky130_fd_sc_hd__o21a_1 _19099_ (.A1(_10848_),
    .A2(_11069_),
    .B1(_11070_),
    .X(_11071_));
 sky130_fd_sc_hd__xnor2_1 _19100_ (.A(_11068_),
    .B(_11071_),
    .Y(_11072_));
 sky130_fd_sc_hd__xnor2_2 _19101_ (.A(_11050_),
    .B(_11072_),
    .Y(_11073_));
 sky130_fd_sc_hd__xnor2_4 _19102_ (.A(_11046_),
    .B(_11073_),
    .Y(_11074_));
 sky130_fd_sc_hd__a21o_1 _19103_ (.A1(_10996_),
    .A2(_11025_),
    .B1(_10994_),
    .X(_11075_));
 sky130_fd_sc_hd__o21a_1 _19104_ (.A1(_10996_),
    .A2(_11025_),
    .B1(_11075_),
    .X(_11076_));
 sky130_fd_sc_hd__xnor2_4 _19105_ (.A(_11074_),
    .B(_11076_),
    .Y(_11077_));
 sky130_fd_sc_hd__or3_1 _19106_ (.A(_11037_),
    .B(_11028_),
    .C(_11077_),
    .X(_11078_));
 sky130_fd_sc_hd__nand2_1 _19107_ (.A(_11028_),
    .B(_11077_),
    .Y(_11079_));
 sky130_fd_sc_hd__o21bai_1 _19108_ (.A1(_11029_),
    .A2(_11077_),
    .B1_N(_10992_),
    .Y(_11080_));
 sky130_fd_sc_hd__o2111a_1 _19109_ (.A1(\top0.pid_d.out[15] ),
    .A2(_09339_),
    .B1(_11080_),
    .C1(_05443_),
    .D1(net435),
    .X(_11081_));
 sky130_fd_sc_hd__xor2_2 _19110_ (.A(\top0.pid_d.out[15] ),
    .B(\top0.pid_d.curr_int[15] ),
    .X(_11082_));
 sky130_fd_sc_hd__o21ai_1 _19111_ (.A1(\top0.pid_d.out[14] ),
    .A2(\top0.pid_d.curr_int[14] ),
    .B1(_11082_),
    .Y(_11083_));
 sky130_fd_sc_hd__inv_2 _19112_ (.A(_11082_),
    .Y(_11084_));
 sky130_fd_sc_hd__a21oi_1 _19113_ (.A1(\top0.pid_d.out[14] ),
    .A2(\top0.pid_d.curr_int[14] ),
    .B1(_11084_),
    .Y(_11085_));
 sky130_fd_sc_hd__mux2_1 _19114_ (.A0(_11083_),
    .A1(_11085_),
    .S(_11033_),
    .X(_11086_));
 sky130_fd_sc_hd__o311a_1 _19115_ (.A1(\top0.pid_d.out[14] ),
    .A2(\top0.pid_d.curr_int[14] ),
    .A3(_11082_),
    .B1(_11086_),
    .C1(net432),
    .X(_11087_));
 sky130_fd_sc_hd__a41o_1 _19116_ (.A1(net432),
    .A2(\top0.pid_d.out[14] ),
    .A3(\top0.pid_d.curr_int[14] ),
    .A4(_11084_),
    .B1(_07137_),
    .X(_11088_));
 sky130_fd_sc_hd__a31o_1 _19117_ (.A1(net435),
    .A2(_11029_),
    .A3(_11077_),
    .B1(_11088_),
    .X(_11089_));
 sky130_fd_sc_hd__o221a_1 _19118_ (.A1(\top0.pid_d.out[15] ),
    .A2(_09339_),
    .B1(_11087_),
    .B2(_11089_),
    .C1(net1019),
    .X(_11090_));
 sky130_fd_sc_hd__a31o_1 _19119_ (.A1(_11078_),
    .A2(_11079_),
    .A3(_11081_),
    .B1(_11090_),
    .X(_00260_));
 sky130_fd_sc_hd__or3_1 _19120_ (.A(\top0.pid_d.state[3] ),
    .B(net438),
    .C(_07136_),
    .X(_11091_));
 sky130_fd_sc_hd__mux2_1 _19121_ (.A0(net433),
    .A1(\top0.pid_d.out_valid ),
    .S(_11091_),
    .X(_11092_));
 sky130_fd_sc_hd__and2_1 _19122_ (.A(_05449_),
    .B(_11092_),
    .X(_11093_));
 sky130_fd_sc_hd__clkbuf_1 _19123_ (.A(_11093_),
    .X(_00261_));
 sky130_fd_sc_hd__nor3_4 _19124_ (.A(\top0.pid_d.state[0] ),
    .B(net433),
    .C(_07136_),
    .Y(_11094_));
 sky130_fd_sc_hd__nor2_4 _19125_ (.A(_05430_),
    .B(_11094_),
    .Y(_11095_));
 sky130_fd_sc_hd__buf_2 _19126_ (.A(_11095_),
    .X(_11096_));
 sky130_fd_sc_hd__and3_2 _19127_ (.A(net437),
    .B(_05442_),
    .C(_11094_),
    .X(_11097_));
 sky130_fd_sc_hd__clkbuf_4 _19128_ (.A(_11097_),
    .X(_11098_));
 sky130_fd_sc_hd__and3_2 _19129_ (.A(\top0.pid_d.state[3] ),
    .B(_05442_),
    .C(_11094_),
    .X(_11099_));
 sky130_fd_sc_hd__buf_2 _19130_ (.A(_11099_),
    .X(_11100_));
 sky130_fd_sc_hd__a22o_1 _19131_ (.A1(\top0.kid[0] ),
    .A2(_11098_),
    .B1(_11100_),
    .B2(\top0.kpd[0] ),
    .X(_11101_));
 sky130_fd_sc_hd__a21o_1 _19132_ (.A1(\top0.pid_d.mult0.a[0] ),
    .A2(_11096_),
    .B1(_11101_),
    .X(_00262_));
 sky130_fd_sc_hd__a22o_1 _19133_ (.A1(\top0.kid[1] ),
    .A2(_11098_),
    .B1(_11100_),
    .B2(\top0.kpd[1] ),
    .X(_11102_));
 sky130_fd_sc_hd__a21o_1 _19134_ (.A1(net424),
    .A2(_11096_),
    .B1(_11102_),
    .X(_00263_));
 sky130_fd_sc_hd__a22o_1 _19135_ (.A1(\top0.kid[2] ),
    .A2(_11098_),
    .B1(_11100_),
    .B2(\top0.kpd[2] ),
    .X(_11103_));
 sky130_fd_sc_hd__a21o_1 _19136_ (.A1(net421),
    .A2(_11096_),
    .B1(_11103_),
    .X(_00264_));
 sky130_fd_sc_hd__a22o_1 _19137_ (.A1(\top0.kid[3] ),
    .A2(_11098_),
    .B1(_11100_),
    .B2(\top0.kpd[3] ),
    .X(_11104_));
 sky130_fd_sc_hd__a21o_1 _19138_ (.A1(net415),
    .A2(_11096_),
    .B1(_11104_),
    .X(_00265_));
 sky130_fd_sc_hd__a22o_1 _19139_ (.A1(\top0.kid[4] ),
    .A2(_11098_),
    .B1(_11100_),
    .B2(\top0.kpd[4] ),
    .X(_11105_));
 sky130_fd_sc_hd__a21o_1 _19140_ (.A1(net410),
    .A2(_11096_),
    .B1(_11105_),
    .X(_00266_));
 sky130_fd_sc_hd__a22o_1 _19141_ (.A1(\top0.kid[5] ),
    .A2(_11098_),
    .B1(_11100_),
    .B2(\top0.kpd[5] ),
    .X(_11106_));
 sky130_fd_sc_hd__a21o_1 _19142_ (.A1(net405),
    .A2(_11096_),
    .B1(_11106_),
    .X(_00267_));
 sky130_fd_sc_hd__a22o_1 _19143_ (.A1(\top0.kid[6] ),
    .A2(_11098_),
    .B1(_11100_),
    .B2(\top0.kpd[6] ),
    .X(_11107_));
 sky130_fd_sc_hd__a21o_1 _19144_ (.A1(net402),
    .A2(_11096_),
    .B1(_11107_),
    .X(_00268_));
 sky130_fd_sc_hd__a22o_1 _19145_ (.A1(\top0.kid[7] ),
    .A2(_11098_),
    .B1(_11100_),
    .B2(\top0.kpd[7] ),
    .X(_11108_));
 sky130_fd_sc_hd__a21o_1 _19146_ (.A1(net397),
    .A2(_11096_),
    .B1(_11108_),
    .X(_00269_));
 sky130_fd_sc_hd__a22o_1 _19147_ (.A1(\top0.kid[8] ),
    .A2(_11098_),
    .B1(_11100_),
    .B2(\top0.kpd[8] ),
    .X(_11109_));
 sky130_fd_sc_hd__a21o_1 _19148_ (.A1(net393),
    .A2(_11096_),
    .B1(_11109_),
    .X(_00270_));
 sky130_fd_sc_hd__a22o_1 _19149_ (.A1(\top0.kid[9] ),
    .A2(_11098_),
    .B1(_11100_),
    .B2(\top0.kpd[9] ),
    .X(_11110_));
 sky130_fd_sc_hd__a21o_1 _19150_ (.A1(net389),
    .A2(_11096_),
    .B1(_11110_),
    .X(_00271_));
 sky130_fd_sc_hd__a22o_1 _19151_ (.A1(\top0.kid[10] ),
    .A2(_11097_),
    .B1(_11099_),
    .B2(\top0.kpd[10] ),
    .X(_11111_));
 sky130_fd_sc_hd__a21o_1 _19152_ (.A1(net383),
    .A2(_11095_),
    .B1(_11111_),
    .X(_00272_));
 sky130_fd_sc_hd__a22o_1 _19153_ (.A1(\top0.kid[11] ),
    .A2(_11097_),
    .B1(_11099_),
    .B2(\top0.kpd[11] ),
    .X(_11112_));
 sky130_fd_sc_hd__a21o_1 _19154_ (.A1(net380),
    .A2(_11095_),
    .B1(_11112_),
    .X(_00273_));
 sky130_fd_sc_hd__a22o_1 _19155_ (.A1(\top0.kid[12] ),
    .A2(_11097_),
    .B1(_11099_),
    .B2(\top0.kpd[12] ),
    .X(_11113_));
 sky130_fd_sc_hd__a21o_1 _19156_ (.A1(net374),
    .A2(_11095_),
    .B1(_11113_),
    .X(_00274_));
 sky130_fd_sc_hd__a22o_1 _19157_ (.A1(\top0.kid[13] ),
    .A2(_11097_),
    .B1(_11099_),
    .B2(\top0.kpd[13] ),
    .X(_11114_));
 sky130_fd_sc_hd__a21o_1 _19158_ (.A1(net372),
    .A2(_11095_),
    .B1(_11114_),
    .X(_00275_));
 sky130_fd_sc_hd__a22o_1 _19159_ (.A1(\top0.kid[14] ),
    .A2(_11097_),
    .B1(_11099_),
    .B2(\top0.kpd[14] ),
    .X(_11115_));
 sky130_fd_sc_hd__a21o_1 _19160_ (.A1(net370),
    .A2(_11095_),
    .B1(_11115_),
    .X(_00276_));
 sky130_fd_sc_hd__a22o_1 _19161_ (.A1(\top0.kid[15] ),
    .A2(_11097_),
    .B1(_11099_),
    .B2(\top0.kpd[15] ),
    .X(_11116_));
 sky130_fd_sc_hd__a21o_1 _19162_ (.A1(net365),
    .A2(_11095_),
    .B1(_11116_),
    .X(_00277_));
 sky130_fd_sc_hd__clkbuf_4 _19163_ (.A(_11094_),
    .X(_11117_));
 sky130_fd_sc_hd__xor2_1 _19164_ (.A(\top0.pid_d.prev_error[0] ),
    .B(\top0.pid_d.curr_error[0] ),
    .X(_11118_));
 sky130_fd_sc_hd__and3_1 _19165_ (.A(\top0.matmul0.done_pass ),
    .B(\top0.matmul0.state[1] ),
    .C(\top0.pid_d.state[3] ),
    .X(_11119_));
 sky130_fd_sc_hd__buf_2 _19166_ (.A(_11119_),
    .X(_11120_));
 sky130_fd_sc_hd__clkbuf_4 _19167_ (.A(_11120_),
    .X(_11121_));
 sky130_fd_sc_hd__or3_1 _19168_ (.A(\top0.pid_d.state[0] ),
    .B(net433),
    .C(_07136_),
    .X(_11122_));
 sky130_fd_sc_hd__buf_2 _19169_ (.A(_11122_),
    .X(_11123_));
 sky130_fd_sc_hd__a221o_1 _19170_ (.A1(net440),
    .A2(_11118_),
    .B1(_11121_),
    .B2(\top0.matmul0.alpha_pass[0] ),
    .C1(_11123_),
    .X(_11124_));
 sky130_fd_sc_hd__o211a_1 _19171_ (.A1(net361),
    .A2(_11117_),
    .B1(_11124_),
    .C1(_10067_),
    .X(_00278_));
 sky130_fd_sc_hd__clkbuf_4 _19172_ (.A(_11123_),
    .X(_11125_));
 sky130_fd_sc_hd__xnor2_1 _19173_ (.A(\top0.pid_d.prev_error[1] ),
    .B(\top0.pid_d.curr_error[1] ),
    .Y(_11126_));
 sky130_fd_sc_hd__and3_1 _19174_ (.A(\top0.pid_d.prev_error[0] ),
    .B(\top0.pid_d.curr_error[0] ),
    .C(_11126_),
    .X(_11127_));
 sky130_fd_sc_hd__a21oi_1 _19175_ (.A1(\top0.pid_d.prev_error[0] ),
    .A2(\top0.pid_d.curr_error[0] ),
    .B1(_11126_),
    .Y(_11128_));
 sky130_fd_sc_hd__o21a_1 _19176_ (.A1(_11127_),
    .A2(_11128_),
    .B1(net439),
    .X(_11129_));
 sky130_fd_sc_hd__xor2_1 _19177_ (.A(\top0.matmul0.alpha_pass[0] ),
    .B(\top0.matmul0.alpha_pass[1] ),
    .X(_11130_));
 sky130_fd_sc_hd__and2_1 _19178_ (.A(_11120_),
    .B(_11130_),
    .X(_11131_));
 sky130_fd_sc_hd__nand2_1 _19179_ (.A(_09356_),
    .B(_11125_),
    .Y(_11132_));
 sky130_fd_sc_hd__o311a_1 _19180_ (.A1(_11125_),
    .A2(_11129_),
    .A3(_11131_),
    .B1(_11132_),
    .C1(_07800_),
    .X(_00279_));
 sky130_fd_sc_hd__or2_1 _19181_ (.A(\top0.pid_d.prev_error[1] ),
    .B(\top0.pid_d.curr_error[1] ),
    .X(_11133_));
 sky130_fd_sc_hd__a22o_1 _19182_ (.A1(\top0.pid_d.prev_error[0] ),
    .A2(\top0.pid_d.curr_error[0] ),
    .B1(\top0.pid_d.prev_error[1] ),
    .B2(\top0.pid_d.curr_error[1] ),
    .X(_11134_));
 sky130_fd_sc_hd__and2_1 _19183_ (.A(_11133_),
    .B(_11134_),
    .X(_11135_));
 sky130_fd_sc_hd__xor2_1 _19184_ (.A(\top0.pid_d.prev_error[2] ),
    .B(\top0.pid_d.curr_error[2] ),
    .X(_11136_));
 sky130_fd_sc_hd__or2_1 _19185_ (.A(_11135_),
    .B(_11136_),
    .X(_11137_));
 sky130_fd_sc_hd__nand2_1 _19186_ (.A(_11135_),
    .B(_11136_),
    .Y(_11138_));
 sky130_fd_sc_hd__and3_1 _19187_ (.A(net439),
    .B(_11137_),
    .C(_11138_),
    .X(_11139_));
 sky130_fd_sc_hd__o21ai_1 _19188_ (.A1(\top0.matmul0.alpha_pass[0] ),
    .A2(\top0.matmul0.alpha_pass[1] ),
    .B1(\top0.matmul0.alpha_pass[2] ),
    .Y(_11140_));
 sky130_fd_sc_hd__or3_1 _19189_ (.A(\top0.matmul0.alpha_pass[0] ),
    .B(\top0.matmul0.alpha_pass[1] ),
    .C(\top0.matmul0.alpha_pass[2] ),
    .X(_11141_));
 sky130_fd_sc_hd__and3_1 _19190_ (.A(_11120_),
    .B(_11140_),
    .C(_11141_),
    .X(_11142_));
 sky130_fd_sc_hd__or2_1 _19191_ (.A(net351),
    .B(_11094_),
    .X(_11143_));
 sky130_fd_sc_hd__o311a_1 _19192_ (.A1(_11125_),
    .A2(_11139_),
    .A3(_11142_),
    .B1(_11143_),
    .C1(_07800_),
    .X(_00280_));
 sky130_fd_sc_hd__a31o_1 _19193_ (.A1(\top0.pid_d.curr_error[2] ),
    .A2(_11133_),
    .A3(_11134_),
    .B1(\top0.pid_d.prev_error[2] ),
    .X(_11144_));
 sky130_fd_sc_hd__o21ai_2 _19194_ (.A1(\top0.pid_d.curr_error[2] ),
    .A2(_11135_),
    .B1(_11144_),
    .Y(_11145_));
 sky130_fd_sc_hd__xnor2_1 _19195_ (.A(\top0.pid_d.prev_error[3] ),
    .B(\top0.pid_d.curr_error[3] ),
    .Y(_11146_));
 sky130_fd_sc_hd__nand2_1 _19196_ (.A(_11145_),
    .B(_11146_),
    .Y(_11147_));
 sky130_fd_sc_hd__or2_1 _19197_ (.A(_11145_),
    .B(_11146_),
    .X(_11148_));
 sky130_fd_sc_hd__and3_1 _19198_ (.A(net439),
    .B(_11147_),
    .C(_11148_),
    .X(_11149_));
 sky130_fd_sc_hd__or2_2 _19199_ (.A(\top0.matmul0.alpha_pass[3] ),
    .B(_11141_),
    .X(_11150_));
 sky130_fd_sc_hd__nand2_1 _19200_ (.A(\top0.matmul0.alpha_pass[3] ),
    .B(_11141_),
    .Y(_11151_));
 sky130_fd_sc_hd__and3_1 _19201_ (.A(_11120_),
    .B(_11150_),
    .C(_11151_),
    .X(_11152_));
 sky130_fd_sc_hd__or2_1 _19202_ (.A(net346),
    .B(_11094_),
    .X(_11153_));
 sky130_fd_sc_hd__o311a_1 _19203_ (.A1(_11125_),
    .A2(_11149_),
    .A3(_11152_),
    .B1(_11153_),
    .C1(_07800_),
    .X(_00281_));
 sky130_fd_sc_hd__inv_2 _19204_ (.A(\top0.pid_d.curr_error[3] ),
    .Y(_11154_));
 sky130_fd_sc_hd__o21ba_1 _19205_ (.A1(_11154_),
    .A2(_11145_),
    .B1_N(\top0.pid_d.prev_error[3] ),
    .X(_11155_));
 sky130_fd_sc_hd__a21o_1 _19206_ (.A1(_11154_),
    .A2(_11145_),
    .B1(_11155_),
    .X(_11156_));
 sky130_fd_sc_hd__xnor2_1 _19207_ (.A(\top0.pid_d.prev_error[4] ),
    .B(\top0.pid_d.curr_error[4] ),
    .Y(_11157_));
 sky130_fd_sc_hd__xnor2_1 _19208_ (.A(_11156_),
    .B(_11157_),
    .Y(_11158_));
 sky130_fd_sc_hd__inv_2 _19209_ (.A(_11158_),
    .Y(_11159_));
 sky130_fd_sc_hd__nor2_1 _19210_ (.A(\top0.matmul0.alpha_pass[4] ),
    .B(_11150_),
    .Y(_11160_));
 sky130_fd_sc_hd__and2_1 _19211_ (.A(\top0.matmul0.alpha_pass[4] ),
    .B(_11150_),
    .X(_11161_));
 sky130_fd_sc_hd__nor2_1 _19212_ (.A(_11160_),
    .B(_11161_),
    .Y(_11162_));
 sky130_fd_sc_hd__a221o_1 _19213_ (.A1(net440),
    .A2(_11159_),
    .B1(_11162_),
    .B2(_11120_),
    .C1(_11123_),
    .X(_11163_));
 sky130_fd_sc_hd__o211a_1 _19214_ (.A1(net342),
    .A2(_11117_),
    .B1(_11163_),
    .C1(_10067_),
    .X(_00282_));
 sky130_fd_sc_hd__inv_2 _19215_ (.A(\top0.pid_d.curr_error[4] ),
    .Y(_11164_));
 sky130_fd_sc_hd__o21ba_1 _19216_ (.A1(_11164_),
    .A2(_11156_),
    .B1_N(\top0.pid_d.prev_error[4] ),
    .X(_11165_));
 sky130_fd_sc_hd__a21o_1 _19217_ (.A1(_11164_),
    .A2(_11156_),
    .B1(_11165_),
    .X(_11166_));
 sky130_fd_sc_hd__xnor2_1 _19218_ (.A(\top0.pid_d.prev_error[5] ),
    .B(\top0.pid_d.curr_error[5] ),
    .Y(_11167_));
 sky130_fd_sc_hd__nand2_1 _19219_ (.A(_11166_),
    .B(_11167_),
    .Y(_11168_));
 sky130_fd_sc_hd__or2_1 _19220_ (.A(_11166_),
    .B(_11167_),
    .X(_11169_));
 sky130_fd_sc_hd__and3_1 _19221_ (.A(net439),
    .B(_11168_),
    .C(_11169_),
    .X(_11170_));
 sky130_fd_sc_hd__xnor2_1 _19222_ (.A(net76),
    .B(_11160_),
    .Y(_11171_));
 sky130_fd_sc_hd__a21o_1 _19223_ (.A1(_11121_),
    .A2(_11171_),
    .B1(_11125_),
    .X(_11172_));
 sky130_fd_sc_hd__o221a_1 _19224_ (.A1(net339),
    .A2(_11117_),
    .B1(_11170_),
    .B2(_11172_),
    .C1(_08889_),
    .X(_00283_));
 sky130_fd_sc_hd__inv_2 _19225_ (.A(\top0.pid_d.curr_error[5] ),
    .Y(_11173_));
 sky130_fd_sc_hd__o21ba_1 _19226_ (.A1(_11173_),
    .A2(_11166_),
    .B1_N(\top0.pid_d.prev_error[5] ),
    .X(_11174_));
 sky130_fd_sc_hd__a21o_1 _19227_ (.A1(_11173_),
    .A2(_11166_),
    .B1(_11174_),
    .X(_11175_));
 sky130_fd_sc_hd__xnor2_1 _19228_ (.A(\top0.pid_d.prev_error[6] ),
    .B(\top0.pid_d.curr_error[6] ),
    .Y(_11176_));
 sky130_fd_sc_hd__nand2_1 _19229_ (.A(_11175_),
    .B(_11176_),
    .Y(_11177_));
 sky130_fd_sc_hd__or2_1 _19230_ (.A(_11175_),
    .B(_11176_),
    .X(_11178_));
 sky130_fd_sc_hd__and3_1 _19231_ (.A(net440),
    .B(_11177_),
    .C(_11178_),
    .X(_11179_));
 sky130_fd_sc_hd__or4_2 _19232_ (.A(\top0.matmul0.alpha_pass[4] ),
    .B(net76),
    .C(\top0.matmul0.alpha_pass[6] ),
    .D(_11150_),
    .X(_11180_));
 sky130_fd_sc_hd__o31ai_2 _19233_ (.A1(\top0.matmul0.alpha_pass[4] ),
    .A2(net76),
    .A3(_11150_),
    .B1(\top0.matmul0.alpha_pass[6] ),
    .Y(_11181_));
 sky130_fd_sc_hd__a31o_1 _19234_ (.A1(_11121_),
    .A2(_11180_),
    .A3(_11181_),
    .B1(_11123_),
    .X(_11182_));
 sky130_fd_sc_hd__o221a_1 _19235_ (.A1(net336),
    .A2(_11117_),
    .B1(_11179_),
    .B2(_11182_),
    .C1(_08889_),
    .X(_00284_));
 sky130_fd_sc_hd__inv_2 _19236_ (.A(\top0.pid_d.curr_error[6] ),
    .Y(_11183_));
 sky130_fd_sc_hd__o21ba_1 _19237_ (.A1(_11183_),
    .A2(_11175_),
    .B1_N(\top0.pid_d.prev_error[6] ),
    .X(_11184_));
 sky130_fd_sc_hd__a21o_1 _19238_ (.A1(_11183_),
    .A2(_11175_),
    .B1(_11184_),
    .X(_11185_));
 sky130_fd_sc_hd__xnor2_1 _19239_ (.A(\top0.pid_d.prev_error[7] ),
    .B(\top0.pid_d.curr_error[7] ),
    .Y(_11186_));
 sky130_fd_sc_hd__nand2_1 _19240_ (.A(_11185_),
    .B(_11186_),
    .Y(_11187_));
 sky130_fd_sc_hd__or2_1 _19241_ (.A(_11185_),
    .B(_11186_),
    .X(_11188_));
 sky130_fd_sc_hd__and3_1 _19242_ (.A(net440),
    .B(_11187_),
    .C(_11188_),
    .X(_11189_));
 sky130_fd_sc_hd__or2_1 _19243_ (.A(\top0.matmul0.alpha_pass[7] ),
    .B(_11180_),
    .X(_11190_));
 sky130_fd_sc_hd__nand2_1 _19244_ (.A(\top0.matmul0.alpha_pass[7] ),
    .B(_11180_),
    .Y(_11191_));
 sky130_fd_sc_hd__and2_1 _19245_ (.A(_11190_),
    .B(_11191_),
    .X(_11192_));
 sky130_fd_sc_hd__a21o_1 _19246_ (.A1(_11121_),
    .A2(_11192_),
    .B1(_11125_),
    .X(_11193_));
 sky130_fd_sc_hd__o221a_1 _19247_ (.A1(net332),
    .A2(_11117_),
    .B1(_11189_),
    .B2(_11193_),
    .C1(_08889_),
    .X(_00285_));
 sky130_fd_sc_hd__inv_2 _19248_ (.A(\top0.pid_d.curr_error[7] ),
    .Y(_11194_));
 sky130_fd_sc_hd__o21ba_1 _19249_ (.A1(_11194_),
    .A2(_11185_),
    .B1_N(\top0.pid_d.prev_error[7] ),
    .X(_11195_));
 sky130_fd_sc_hd__a21o_1 _19250_ (.A1(_11194_),
    .A2(_11185_),
    .B1(_11195_),
    .X(_11196_));
 sky130_fd_sc_hd__xnor2_1 _19251_ (.A(\top0.pid_d.prev_error[8] ),
    .B(\top0.pid_d.curr_error[8] ),
    .Y(_11197_));
 sky130_fd_sc_hd__nand2_1 _19252_ (.A(_11196_),
    .B(_11197_),
    .Y(_11198_));
 sky130_fd_sc_hd__or2_1 _19253_ (.A(_11196_),
    .B(_11197_),
    .X(_11199_));
 sky130_fd_sc_hd__and3_1 _19254_ (.A(net438),
    .B(_11198_),
    .C(_11199_),
    .X(_11200_));
 sky130_fd_sc_hd__xor2_1 _19255_ (.A(net1024),
    .B(_11190_),
    .X(_11201_));
 sky130_fd_sc_hd__a21o_1 _19256_ (.A1(_11121_),
    .A2(_11201_),
    .B1(_11125_),
    .X(_11202_));
 sky130_fd_sc_hd__o221a_1 _19257_ (.A1(net329),
    .A2(_11117_),
    .B1(_11200_),
    .B2(_11202_),
    .C1(_08889_),
    .X(_00286_));
 sky130_fd_sc_hd__inv_2 _19258_ (.A(\top0.pid_d.curr_error[8] ),
    .Y(_11203_));
 sky130_fd_sc_hd__o21ba_1 _19259_ (.A1(_11203_),
    .A2(_11196_),
    .B1_N(\top0.pid_d.prev_error[8] ),
    .X(_11204_));
 sky130_fd_sc_hd__a21o_1 _19260_ (.A1(_11203_),
    .A2(_11196_),
    .B1(_11204_),
    .X(_11205_));
 sky130_fd_sc_hd__xnor2_1 _19261_ (.A(\top0.pid_d.prev_error[9] ),
    .B(\top0.pid_d.curr_error[9] ),
    .Y(_11206_));
 sky130_fd_sc_hd__nand2_1 _19262_ (.A(_11205_),
    .B(_11206_),
    .Y(_11207_));
 sky130_fd_sc_hd__or2_1 _19263_ (.A(_11205_),
    .B(_11206_),
    .X(_11208_));
 sky130_fd_sc_hd__and3_1 _19264_ (.A(net439),
    .B(_11207_),
    .C(_11208_),
    .X(_11209_));
 sky130_fd_sc_hd__or3_1 _19265_ (.A(net1024),
    .B(\top0.matmul0.alpha_pass[9] ),
    .C(_11190_),
    .X(_11210_));
 sky130_fd_sc_hd__o21ai_1 _19266_ (.A1(net1024),
    .A2(_11190_),
    .B1(\top0.matmul0.alpha_pass[9] ),
    .Y(_11211_));
 sky130_fd_sc_hd__and3_1 _19267_ (.A(_11120_),
    .B(_11210_),
    .C(_11211_),
    .X(_11212_));
 sky130_fd_sc_hd__or2_1 _19268_ (.A(net326),
    .B(_11094_),
    .X(_11213_));
 sky130_fd_sc_hd__o311a_1 _19269_ (.A1(_11125_),
    .A2(_11209_),
    .A3(_11212_),
    .B1(_11213_),
    .C1(_07800_),
    .X(_00287_));
 sky130_fd_sc_hd__inv_2 _19270_ (.A(\top0.pid_d.curr_error[9] ),
    .Y(_11214_));
 sky130_fd_sc_hd__o21ba_1 _19271_ (.A1(_11214_),
    .A2(_11205_),
    .B1_N(\top0.pid_d.prev_error[9] ),
    .X(_11215_));
 sky130_fd_sc_hd__a21o_1 _19272_ (.A1(_11214_),
    .A2(_11205_),
    .B1(_11215_),
    .X(_11216_));
 sky130_fd_sc_hd__xnor2_1 _19273_ (.A(\top0.pid_d.prev_error[10] ),
    .B(\top0.pid_d.curr_error[10] ),
    .Y(_11217_));
 sky130_fd_sc_hd__nand2_1 _19274_ (.A(_11216_),
    .B(_11217_),
    .Y(_11218_));
 sky130_fd_sc_hd__or2_1 _19275_ (.A(_11216_),
    .B(_11217_),
    .X(_11219_));
 sky130_fd_sc_hd__and3_1 _19276_ (.A(net438),
    .B(_11218_),
    .C(_11219_),
    .X(_11220_));
 sky130_fd_sc_hd__or2_1 _19277_ (.A(\top0.matmul0.alpha_pass[10] ),
    .B(_11210_),
    .X(_11221_));
 sky130_fd_sc_hd__nand2_1 _19278_ (.A(\top0.matmul0.alpha_pass[10] ),
    .B(_11210_),
    .Y(_11222_));
 sky130_fd_sc_hd__and2_1 _19279_ (.A(_11221_),
    .B(_11222_),
    .X(_11223_));
 sky130_fd_sc_hd__a21o_1 _19280_ (.A1(_11121_),
    .A2(_11223_),
    .B1(_11123_),
    .X(_11224_));
 sky130_fd_sc_hd__o221a_1 _19281_ (.A1(net322),
    .A2(_11117_),
    .B1(_11220_),
    .B2(_11224_),
    .C1(_08889_),
    .X(_00288_));
 sky130_fd_sc_hd__inv_2 _19282_ (.A(\top0.pid_d.curr_error[10] ),
    .Y(_11225_));
 sky130_fd_sc_hd__o21ba_1 _19283_ (.A1(_11225_),
    .A2(_11216_),
    .B1_N(\top0.pid_d.prev_error[10] ),
    .X(_11226_));
 sky130_fd_sc_hd__a21o_1 _19284_ (.A1(_11225_),
    .A2(_11216_),
    .B1(_11226_),
    .X(_11227_));
 sky130_fd_sc_hd__xnor2_1 _19285_ (.A(\top0.pid_d.prev_error[11] ),
    .B(\top0.pid_d.curr_error[11] ),
    .Y(_11228_));
 sky130_fd_sc_hd__nand2_1 _19286_ (.A(_11227_),
    .B(_11228_),
    .Y(_11229_));
 sky130_fd_sc_hd__or2_1 _19287_ (.A(_11227_),
    .B(_11228_),
    .X(_11230_));
 sky130_fd_sc_hd__and3_1 _19288_ (.A(net437),
    .B(_11229_),
    .C(_11230_),
    .X(_11231_));
 sky130_fd_sc_hd__xor2_1 _19289_ (.A(\top0.matmul0.alpha_pass[11] ),
    .B(_11221_),
    .X(_11232_));
 sky130_fd_sc_hd__a21o_1 _19290_ (.A1(_11121_),
    .A2(_11232_),
    .B1(_11123_),
    .X(_11233_));
 sky130_fd_sc_hd__o221a_1 _19291_ (.A1(\top0.pid_d.mult0.b[11] ),
    .A2(_11094_),
    .B1(_11231_),
    .B2(_11233_),
    .C1(_08889_),
    .X(_00289_));
 sky130_fd_sc_hd__and2_1 _19292_ (.A(\top0.pid_d.prev_error[12] ),
    .B(\top0.pid_d.curr_error[12] ),
    .X(_11234_));
 sky130_fd_sc_hd__nor2_1 _19293_ (.A(\top0.pid_d.prev_error[12] ),
    .B(\top0.pid_d.curr_error[12] ),
    .Y(_11235_));
 sky130_fd_sc_hd__nor2_1 _19294_ (.A(_11234_),
    .B(_11235_),
    .Y(_11236_));
 sky130_fd_sc_hd__nor2_1 _19295_ (.A(\top0.pid_d.prev_error[11] ),
    .B(\top0.pid_d.curr_error[11] ),
    .Y(_11237_));
 sky130_fd_sc_hd__nand2_1 _19296_ (.A(\top0.pid_d.prev_error[11] ),
    .B(\top0.pid_d.curr_error[11] ),
    .Y(_11238_));
 sky130_fd_sc_hd__o21a_1 _19297_ (.A1(_11227_),
    .A2(_11237_),
    .B1(_11238_),
    .X(_11239_));
 sky130_fd_sc_hd__xnor2_1 _19298_ (.A(_11236_),
    .B(_11239_),
    .Y(_11240_));
 sky130_fd_sc_hd__or3_1 _19299_ (.A(\top0.matmul0.alpha_pass[11] ),
    .B(\top0.matmul0.alpha_pass[12] ),
    .C(_11221_),
    .X(_11241_));
 sky130_fd_sc_hd__o21ai_1 _19300_ (.A1(\top0.matmul0.alpha_pass[11] ),
    .A2(_11221_),
    .B1(\top0.matmul0.alpha_pass[12] ),
    .Y(_11242_));
 sky130_fd_sc_hd__and3_1 _19301_ (.A(_11120_),
    .B(_11241_),
    .C(_11242_),
    .X(_11243_));
 sky130_fd_sc_hd__a211o_1 _19302_ (.A1(net437),
    .A2(_11240_),
    .B1(_11243_),
    .C1(_11125_),
    .X(_11244_));
 sky130_fd_sc_hd__o211a_1 _19303_ (.A1(net315),
    .A2(_11117_),
    .B1(_11244_),
    .C1(_10067_),
    .X(_00290_));
 sky130_fd_sc_hd__or2_1 _19304_ (.A(\top0.matmul0.alpha_pass[13] ),
    .B(_11241_),
    .X(_11245_));
 sky130_fd_sc_hd__nand2_1 _19305_ (.A(\top0.matmul0.alpha_pass[13] ),
    .B(_11241_),
    .Y(_11246_));
 sky130_fd_sc_hd__and3_1 _19306_ (.A(_11119_),
    .B(_11245_),
    .C(_11246_),
    .X(_11247_));
 sky130_fd_sc_hd__nand2_1 _19307_ (.A(\top0.pid_d.prev_error[12] ),
    .B(\top0.pid_d.curr_error[12] ),
    .Y(_11248_));
 sky130_fd_sc_hd__a21o_1 _19308_ (.A1(_11248_),
    .A2(_11239_),
    .B1(_11235_),
    .X(_11249_));
 sky130_fd_sc_hd__xor2_1 _19309_ (.A(\top0.pid_d.prev_error[13] ),
    .B(\top0.pid_d.curr_error[13] ),
    .X(_11250_));
 sky130_fd_sc_hd__xnor2_1 _19310_ (.A(_11249_),
    .B(_11250_),
    .Y(_11251_));
 sky130_fd_sc_hd__nand2_1 _19311_ (.A(net437),
    .B(_11251_),
    .Y(_11252_));
 sky130_fd_sc_hd__or3b_1 _19312_ (.A(_11247_),
    .B(_11123_),
    .C_N(_11252_),
    .X(_11253_));
 sky130_fd_sc_hd__o211a_1 _19313_ (.A1(net313),
    .A2(_11117_),
    .B1(_11253_),
    .C1(_10067_),
    .X(_00291_));
 sky130_fd_sc_hd__and2_1 _19314_ (.A(\top0.pid_d.prev_error[14] ),
    .B(\top0.pid_d.curr_error[14] ),
    .X(_11254_));
 sky130_fd_sc_hd__nor2_1 _19315_ (.A(\top0.pid_d.prev_error[14] ),
    .B(\top0.pid_d.curr_error[14] ),
    .Y(_11255_));
 sky130_fd_sc_hd__nor2_1 _19316_ (.A(\top0.pid_d.prev_error[13] ),
    .B(\top0.pid_d.curr_error[13] ),
    .Y(_11256_));
 sky130_fd_sc_hd__nand2_1 _19317_ (.A(\top0.pid_d.prev_error[13] ),
    .B(\top0.pid_d.curr_error[13] ),
    .Y(_11257_));
 sky130_fd_sc_hd__o21ai_1 _19318_ (.A1(_11249_),
    .A2(_11256_),
    .B1(_11257_),
    .Y(_11258_));
 sky130_fd_sc_hd__o21ai_1 _19319_ (.A1(_11254_),
    .A2(_11255_),
    .B1(_11258_),
    .Y(_11259_));
 sky130_fd_sc_hd__or3_1 _19320_ (.A(_11258_),
    .B(_11254_),
    .C(_11255_),
    .X(_11260_));
 sky130_fd_sc_hd__a21bo_1 _19321_ (.A1(_11259_),
    .A2(_11260_),
    .B1_N(net437),
    .X(_11261_));
 sky130_fd_sc_hd__nor2_1 _19322_ (.A(\top0.matmul0.alpha_pass[14] ),
    .B(_11245_),
    .Y(_11262_));
 sky130_fd_sc_hd__and2_1 _19323_ (.A(\top0.matmul0.alpha_pass[14] ),
    .B(_11245_),
    .X(_11263_));
 sky130_fd_sc_hd__nor2_1 _19324_ (.A(_11262_),
    .B(_11263_),
    .Y(_11264_));
 sky130_fd_sc_hd__a21oi_1 _19325_ (.A1(_11121_),
    .A2(_11264_),
    .B1(_11123_),
    .Y(_11265_));
 sky130_fd_sc_hd__a221oi_2 _19326_ (.A1(_10311_),
    .A2(_11125_),
    .B1(_11261_),
    .B2(_11265_),
    .C1(_05430_),
    .Y(_00292_));
 sky130_fd_sc_hd__o21ba_1 _19327_ (.A1(_11258_),
    .A2(_11254_),
    .B1_N(_11255_),
    .X(_11266_));
 sky130_fd_sc_hd__xnor2_1 _19328_ (.A(\top0.pid_d.prev_error[15] ),
    .B(\top0.pid_d.curr_error[15] ),
    .Y(_11267_));
 sky130_fd_sc_hd__xnor2_2 _19329_ (.A(_11266_),
    .B(_11267_),
    .Y(_11268_));
 sky130_fd_sc_hd__xnor2_1 _19330_ (.A(\top0.matmul0.alpha_pass[15] ),
    .B(_11262_),
    .Y(_11269_));
 sky130_fd_sc_hd__a221o_1 _19331_ (.A1(net438),
    .A2(_11268_),
    .B1(_11269_),
    .B2(_11120_),
    .C1(_11123_),
    .X(_11270_));
 sky130_fd_sc_hd__o211a_1 _19332_ (.A1(net307),
    .A2(_11117_),
    .B1(_11270_),
    .C1(_10067_),
    .X(_00293_));
 sky130_fd_sc_hd__and3_1 _19333_ (.A(\top0.matmul0.alpha_pass[0] ),
    .B(_05443_),
    .C(_11120_),
    .X(_11271_));
 sky130_fd_sc_hd__or2_1 _19334_ (.A(_00006_),
    .B(_11095_),
    .X(_11272_));
 sky130_fd_sc_hd__buf_2 _19335_ (.A(_11272_),
    .X(_11273_));
 sky130_fd_sc_hd__mux2_1 _19336_ (.A0(_11271_),
    .A1(\top0.pid_d.curr_error[0] ),
    .S(_11273_),
    .X(_11274_));
 sky130_fd_sc_hd__clkbuf_1 _19337_ (.A(_11274_),
    .X(_00294_));
 sky130_fd_sc_hd__clkbuf_4 _19338_ (.A(_11273_),
    .X(_11275_));
 sky130_fd_sc_hd__nor2_1 _19339_ (.A(net438),
    .B(_11123_),
    .Y(_11276_));
 sky130_fd_sc_hd__and2_1 _19340_ (.A(_05442_),
    .B(_11276_),
    .X(_11277_));
 sky130_fd_sc_hd__buf_2 _19341_ (.A(_11277_),
    .X(_11278_));
 sky130_fd_sc_hd__a22o_1 _19342_ (.A1(\top0.pid_d.curr_error[1] ),
    .A2(_11275_),
    .B1(_11278_),
    .B2(_11131_),
    .X(_00295_));
 sky130_fd_sc_hd__a22o_1 _19343_ (.A1(net986),
    .A2(_11275_),
    .B1(_11278_),
    .B2(_11142_),
    .X(_00296_));
 sky130_fd_sc_hd__a22o_1 _19344_ (.A1(\top0.pid_d.curr_error[3] ),
    .A2(_11275_),
    .B1(_11278_),
    .B2(_11152_),
    .X(_00297_));
 sky130_fd_sc_hd__a32o_1 _19345_ (.A1(_11121_),
    .A2(_11162_),
    .A3(_11278_),
    .B1(_11273_),
    .B2(\top0.pid_d.curr_error[4] ),
    .X(_00298_));
 sky130_fd_sc_hd__and3_1 _19346_ (.A(_05439_),
    .B(_00003_),
    .C(_11276_),
    .X(_11279_));
 sky130_fd_sc_hd__a22o_1 _19347_ (.A1(\top0.pid_d.curr_error[5] ),
    .A2(_11275_),
    .B1(_11279_),
    .B2(_11171_),
    .X(_00299_));
 sky130_fd_sc_hd__a32o_1 _19348_ (.A1(_11180_),
    .A2(_11181_),
    .A3(_11279_),
    .B1(_11273_),
    .B2(\top0.pid_d.curr_error[6] ),
    .X(_00300_));
 sky130_fd_sc_hd__and3_1 _19349_ (.A(_05443_),
    .B(_11120_),
    .C(_11276_),
    .X(_11280_));
 sky130_fd_sc_hd__clkbuf_2 _19350_ (.A(_11280_),
    .X(_11281_));
 sky130_fd_sc_hd__a22o_1 _19351_ (.A1(net927),
    .A2(_11275_),
    .B1(_11281_),
    .B2(_11192_),
    .X(_00301_));
 sky130_fd_sc_hd__a22o_1 _19352_ (.A1(net923),
    .A2(_11275_),
    .B1(_11281_),
    .B2(_11201_),
    .X(_00302_));
 sky130_fd_sc_hd__a22o_1 _19353_ (.A1(\top0.pid_d.curr_error[9] ),
    .A2(_11275_),
    .B1(_11278_),
    .B2(_11212_),
    .X(_00303_));
 sky130_fd_sc_hd__a22o_1 _19354_ (.A1(net931),
    .A2(_11275_),
    .B1(_11281_),
    .B2(_11223_),
    .X(_00304_));
 sky130_fd_sc_hd__a22o_1 _19355_ (.A1(net760),
    .A2(_11275_),
    .B1(_11281_),
    .B2(_11232_),
    .X(_00305_));
 sky130_fd_sc_hd__mux2_1 _19356_ (.A0(\top0.pid_d.curr_error[12] ),
    .A1(_11243_),
    .S(_11276_),
    .X(_11282_));
 sky130_fd_sc_hd__and2_1 _19357_ (.A(_05449_),
    .B(_11282_),
    .X(_11283_));
 sky130_fd_sc_hd__clkbuf_1 _19358_ (.A(_11283_),
    .X(_00306_));
 sky130_fd_sc_hd__a22o_1 _19359_ (.A1(net910),
    .A2(_11275_),
    .B1(_11278_),
    .B2(_11247_),
    .X(_00307_));
 sky130_fd_sc_hd__a32o_1 _19360_ (.A1(_11121_),
    .A2(_11264_),
    .A3(_11278_),
    .B1(_11273_),
    .B2(net765),
    .X(_00308_));
 sky130_fd_sc_hd__a22o_1 _19361_ (.A1(net722),
    .A2(_11273_),
    .B1(_11281_),
    .B2(_11269_),
    .X(_00309_));
 sky130_fd_sc_hd__o21a_2 _19362_ (.A1(net433),
    .A2(_07137_),
    .B1(_05441_),
    .X(_11284_));
 sky130_fd_sc_hd__clkbuf_4 _19363_ (.A(_11284_),
    .X(_11285_));
 sky130_fd_sc_hd__and2b_1 _19364_ (.A_N(_11284_),
    .B(_00006_),
    .X(_11286_));
 sky130_fd_sc_hd__buf_2 _19365_ (.A(_11286_),
    .X(_11287_));
 sky130_fd_sc_hd__clkbuf_4 _19366_ (.A(_11287_),
    .X(_11288_));
 sky130_fd_sc_hd__a22o_1 _19367_ (.A1(\top0.pid_d.prev_error[0] ),
    .A2(_11285_),
    .B1(_11288_),
    .B2(net940),
    .X(_00310_));
 sky130_fd_sc_hd__a22o_1 _19368_ (.A1(net961),
    .A2(_11285_),
    .B1(_11288_),
    .B2(\top0.pid_d.curr_error[1] ),
    .X(_00311_));
 sky130_fd_sc_hd__a22o_1 _19369_ (.A1(net892),
    .A2(_11285_),
    .B1(_11288_),
    .B2(\top0.pid_d.curr_error[2] ),
    .X(_00312_));
 sky130_fd_sc_hd__a22o_1 _19370_ (.A1(net872),
    .A2(_11285_),
    .B1(_11288_),
    .B2(\top0.pid_d.curr_error[3] ),
    .X(_00313_));
 sky130_fd_sc_hd__a22o_1 _19371_ (.A1(net878),
    .A2(_11285_),
    .B1(_11288_),
    .B2(\top0.pid_d.curr_error[4] ),
    .X(_00314_));
 sky130_fd_sc_hd__a22o_1 _19372_ (.A1(net884),
    .A2(_11285_),
    .B1(_11288_),
    .B2(\top0.pid_d.curr_error[5] ),
    .X(_00315_));
 sky130_fd_sc_hd__a22o_1 _19373_ (.A1(net879),
    .A2(_11285_),
    .B1(_11288_),
    .B2(\top0.pid_d.curr_error[6] ),
    .X(_00316_));
 sky130_fd_sc_hd__a22o_1 _19374_ (.A1(net880),
    .A2(_11285_),
    .B1(_11288_),
    .B2(\top0.pid_d.curr_error[7] ),
    .X(_00317_));
 sky130_fd_sc_hd__a22o_1 _19375_ (.A1(net876),
    .A2(_11285_),
    .B1(_11288_),
    .B2(\top0.pid_d.curr_error[8] ),
    .X(_00318_));
 sky130_fd_sc_hd__a22o_1 _19376_ (.A1(net889),
    .A2(_11285_),
    .B1(_11288_),
    .B2(\top0.pid_d.curr_error[9] ),
    .X(_00319_));
 sky130_fd_sc_hd__a22o_1 _19377_ (.A1(net874),
    .A2(_11284_),
    .B1(_11287_),
    .B2(\top0.pid_d.curr_error[10] ),
    .X(_00320_));
 sky130_fd_sc_hd__a22o_1 _19378_ (.A1(\top0.pid_d.prev_error[11] ),
    .A2(_11284_),
    .B1(_11287_),
    .B2(net760),
    .X(_00321_));
 sky130_fd_sc_hd__a22o_1 _19379_ (.A1(net903),
    .A2(_11284_),
    .B1(_11287_),
    .B2(\top0.pid_d.curr_error[12] ),
    .X(_00322_));
 sky130_fd_sc_hd__a22o_1 _19380_ (.A1(\top0.pid_d.prev_error[13] ),
    .A2(_11284_),
    .B1(_11287_),
    .B2(net910),
    .X(_00323_));
 sky130_fd_sc_hd__a22o_1 _19381_ (.A1(\top0.pid_d.prev_error[14] ),
    .A2(_11284_),
    .B1(_11287_),
    .B2(net765),
    .X(_00324_));
 sky130_fd_sc_hd__a22o_1 _19382_ (.A1(\top0.pid_d.prev_error[15] ),
    .A2(_11284_),
    .B1(_11287_),
    .B2(net722),
    .X(_00325_));
 sky130_fd_sc_hd__o31a_4 _19383_ (.A1(\top0.pid_d.state[0] ),
    .A2(\top0.pid_d.state[3] ),
    .A3(net433),
    .B1(_05441_),
    .X(_11289_));
 sky130_fd_sc_hd__clkbuf_4 _19384_ (.A(_11289_),
    .X(_11290_));
 sky130_fd_sc_hd__o21ai_1 _19385_ (.A1(net437),
    .A2(_07136_),
    .B1(_05441_),
    .Y(_11291_));
 sky130_fd_sc_hd__nor2_2 _19386_ (.A(_11289_),
    .B(_11291_),
    .Y(_11292_));
 sky130_fd_sc_hd__clkbuf_4 _19387_ (.A(_11292_),
    .X(_11293_));
 sky130_fd_sc_hd__xor2_1 _19388_ (.A(\top0.pid_d.curr_int[0] ),
    .B(\top0.pid_d.prev_int[0] ),
    .X(_11294_));
 sky130_fd_sc_hd__a22o_1 _19389_ (.A1(net439),
    .A2(_11118_),
    .B1(_11294_),
    .B2(net442),
    .X(_11295_));
 sky130_fd_sc_hd__a31o_1 _19390_ (.A1(net431),
    .A2(_09892_),
    .A3(_09893_),
    .B1(_11295_),
    .X(_11296_));
 sky130_fd_sc_hd__a22o_1 _19391_ (.A1(\top0.pid_d.curr_int[0] ),
    .A2(_11290_),
    .B1(_11293_),
    .B2(_11296_),
    .X(_00326_));
 sky130_fd_sc_hd__nand2_1 _19392_ (.A(\top0.pid_d.curr_int[0] ),
    .B(\top0.pid_d.prev_int[0] ),
    .Y(_11297_));
 sky130_fd_sc_hd__xor2_1 _19393_ (.A(\top0.pid_d.curr_int[1] ),
    .B(\top0.pid_d.prev_int[1] ),
    .X(_11298_));
 sky130_fd_sc_hd__xnor2_1 _19394_ (.A(_11297_),
    .B(_11298_),
    .Y(_11299_));
 sky130_fd_sc_hd__a221o_1 _19395_ (.A1(net431),
    .A2(_09977_),
    .B1(_11299_),
    .B2(net442),
    .C1(_11129_),
    .X(_11300_));
 sky130_fd_sc_hd__a22o_1 _19396_ (.A1(\top0.pid_d.curr_int[1] ),
    .A2(_11290_),
    .B1(_11293_),
    .B2(_11300_),
    .X(_00327_));
 sky130_fd_sc_hd__nand2_1 _19397_ (.A(\top0.pid_d.curr_int[1] ),
    .B(\top0.pid_d.prev_int[1] ),
    .Y(_11301_));
 sky130_fd_sc_hd__o211ai_2 _19398_ (.A1(\top0.pid_d.curr_int[1] ),
    .A2(\top0.pid_d.prev_int[1] ),
    .B1(\top0.pid_d.prev_int[0] ),
    .C1(\top0.pid_d.curr_int[0] ),
    .Y(_11302_));
 sky130_fd_sc_hd__nand2_1 _19399_ (.A(_11301_),
    .B(_11302_),
    .Y(_11303_));
 sky130_fd_sc_hd__xnor2_1 _19400_ (.A(\top0.pid_d.curr_int[2] ),
    .B(\top0.pid_d.prev_int[2] ),
    .Y(_11304_));
 sky130_fd_sc_hd__xnor2_1 _19401_ (.A(_11303_),
    .B(_11304_),
    .Y(_11305_));
 sky130_fd_sc_hd__a221o_1 _19402_ (.A1(net431),
    .A2(_10065_),
    .B1(_11305_),
    .B2(net442),
    .C1(_11139_),
    .X(_11306_));
 sky130_fd_sc_hd__a22o_1 _19403_ (.A1(\top0.pid_d.curr_int[2] ),
    .A2(_11290_),
    .B1(_11293_),
    .B2(_11306_),
    .X(_00328_));
 sky130_fd_sc_hd__inv_2 _19404_ (.A(\top0.pid_d.prev_int[2] ),
    .Y(_11307_));
 sky130_fd_sc_hd__a21o_1 _19405_ (.A1(_11301_),
    .A2(_11302_),
    .B1(_11307_),
    .X(_11308_));
 sky130_fd_sc_hd__inv_2 _19406_ (.A(\top0.pid_d.curr_int[2] ),
    .Y(_11309_));
 sky130_fd_sc_hd__a31o_1 _19407_ (.A1(_11307_),
    .A2(_11301_),
    .A3(_11302_),
    .B1(_11309_),
    .X(_11310_));
 sky130_fd_sc_hd__nand2_1 _19408_ (.A(_11308_),
    .B(_11310_),
    .Y(_11311_));
 sky130_fd_sc_hd__xnor2_1 _19409_ (.A(\top0.pid_d.curr_int[3] ),
    .B(\top0.pid_d.prev_int[3] ),
    .Y(_11312_));
 sky130_fd_sc_hd__xnor2_1 _19410_ (.A(_11311_),
    .B(_11312_),
    .Y(_11313_));
 sky130_fd_sc_hd__a221o_1 _19411_ (.A1(net431),
    .A2(_10156_),
    .B1(_11313_),
    .B2(net442),
    .C1(_11149_),
    .X(_11314_));
 sky130_fd_sc_hd__a22o_1 _19412_ (.A1(\top0.pid_d.curr_int[3] ),
    .A2(_11290_),
    .B1(_11293_),
    .B2(_11314_),
    .X(_00329_));
 sky130_fd_sc_hd__inv_2 _19413_ (.A(\top0.pid_d.prev_int[3] ),
    .Y(_11315_));
 sky130_fd_sc_hd__inv_2 _19414_ (.A(\top0.pid_d.curr_int[3] ),
    .Y(_11316_));
 sky130_fd_sc_hd__a31o_1 _19415_ (.A1(_11315_),
    .A2(_11308_),
    .A3(_11310_),
    .B1(_11316_),
    .X(_11317_));
 sky130_fd_sc_hd__a21bo_1 _19416_ (.A1(\top0.pid_d.prev_int[3] ),
    .A2(_11311_),
    .B1_N(_11317_),
    .X(_11318_));
 sky130_fd_sc_hd__xor2_1 _19417_ (.A(\top0.pid_d.curr_int[4] ),
    .B(\top0.pid_d.prev_int[4] ),
    .X(_11319_));
 sky130_fd_sc_hd__or2_1 _19418_ (.A(_11318_),
    .B(_11319_),
    .X(_11320_));
 sky130_fd_sc_hd__nand2_1 _19419_ (.A(_11318_),
    .B(_11319_),
    .Y(_11321_));
 sky130_fd_sc_hd__a32o_1 _19420_ (.A1(net442),
    .A2(_11320_),
    .A3(_11321_),
    .B1(net436),
    .B2(_11159_),
    .X(_11322_));
 sky130_fd_sc_hd__a21o_1 _19421_ (.A1(net431),
    .A2(_10243_),
    .B1(_11322_),
    .X(_11323_));
 sky130_fd_sc_hd__a22o_1 _19422_ (.A1(\top0.pid_d.curr_int[4] ),
    .A2(_11290_),
    .B1(_11293_),
    .B2(_11323_),
    .X(_00330_));
 sky130_fd_sc_hd__a21o_1 _19423_ (.A1(\top0.pid_d.prev_int[4] ),
    .A2(_11318_),
    .B1(\top0.pid_d.curr_int[4] ),
    .X(_11324_));
 sky130_fd_sc_hd__o21a_1 _19424_ (.A1(\top0.pid_d.prev_int[4] ),
    .A2(_11318_),
    .B1(_11324_),
    .X(_11325_));
 sky130_fd_sc_hd__xnor2_1 _19425_ (.A(\top0.pid_d.curr_int[5] ),
    .B(\top0.pid_d.prev_int[5] ),
    .Y(_11326_));
 sky130_fd_sc_hd__xnor2_1 _19426_ (.A(_11325_),
    .B(_11326_),
    .Y(_11327_));
 sky130_fd_sc_hd__a221o_1 _19427_ (.A1(net431),
    .A2(_10333_),
    .B1(_11327_),
    .B2(net442),
    .C1(_11170_),
    .X(_11328_));
 sky130_fd_sc_hd__a22o_1 _19428_ (.A1(\top0.pid_d.curr_int[5] ),
    .A2(_11290_),
    .B1(_11293_),
    .B2(_11328_),
    .X(_00331_));
 sky130_fd_sc_hd__a21o_1 _19429_ (.A1(\top0.pid_d.prev_int[5] ),
    .A2(_11325_),
    .B1(\top0.pid_d.curr_int[5] ),
    .X(_11329_));
 sky130_fd_sc_hd__o21ai_2 _19430_ (.A1(\top0.pid_d.prev_int[5] ),
    .A2(_11325_),
    .B1(_11329_),
    .Y(_11330_));
 sky130_fd_sc_hd__xor2_1 _19431_ (.A(\top0.pid_d.curr_int[6] ),
    .B(\top0.pid_d.prev_int[6] ),
    .X(_11331_));
 sky130_fd_sc_hd__xnor2_1 _19432_ (.A(_11330_),
    .B(_11331_),
    .Y(_11332_));
 sky130_fd_sc_hd__a221o_1 _19433_ (.A1(net431),
    .A2(_10423_),
    .B1(_11332_),
    .B2(net442),
    .C1(_11179_),
    .X(_11333_));
 sky130_fd_sc_hd__a22o_1 _19434_ (.A1(\top0.pid_d.curr_int[6] ),
    .A2(_11290_),
    .B1(_11293_),
    .B2(_11333_),
    .X(_00332_));
 sky130_fd_sc_hd__inv_2 _19435_ (.A(\top0.pid_d.prev_int[6] ),
    .Y(_11334_));
 sky130_fd_sc_hd__o21a_1 _19436_ (.A1(_11334_),
    .A2(_11330_),
    .B1(_10427_),
    .X(_11335_));
 sky130_fd_sc_hd__a21o_1 _19437_ (.A1(_11334_),
    .A2(_11330_),
    .B1(_11335_),
    .X(_11336_));
 sky130_fd_sc_hd__xor2_1 _19438_ (.A(\top0.pid_d.curr_int[7] ),
    .B(\top0.pid_d.prev_int[7] ),
    .X(_11337_));
 sky130_fd_sc_hd__xnor2_1 _19439_ (.A(_11336_),
    .B(_11337_),
    .Y(_11338_));
 sky130_fd_sc_hd__a221o_1 _19440_ (.A1(\top0.pid_d.state[5] ),
    .A2(_10508_),
    .B1(_11338_),
    .B2(net442),
    .C1(_11189_),
    .X(_11339_));
 sky130_fd_sc_hd__a22o_1 _19441_ (.A1(\top0.pid_d.curr_int[7] ),
    .A2(_11290_),
    .B1(_11293_),
    .B2(_11339_),
    .X(_00333_));
 sky130_fd_sc_hd__and2_1 _19442_ (.A(net431),
    .B(_11292_),
    .X(_11340_));
 sky130_fd_sc_hd__buf_2 _19443_ (.A(_11340_),
    .X(_11341_));
 sky130_fd_sc_hd__inv_2 _19444_ (.A(\top0.pid_d.prev_int[7] ),
    .Y(_11342_));
 sky130_fd_sc_hd__nor2_1 _19445_ (.A(_11342_),
    .B(_11336_),
    .Y(_11343_));
 sky130_fd_sc_hd__nand2_1 _19446_ (.A(_11342_),
    .B(_11336_),
    .Y(_11344_));
 sky130_fd_sc_hd__o21ai_2 _19447_ (.A1(\top0.pid_d.curr_int[7] ),
    .A2(_11343_),
    .B1(_11344_),
    .Y(_11345_));
 sky130_fd_sc_hd__xnor2_1 _19448_ (.A(\top0.pid_d.curr_int[8] ),
    .B(\top0.pid_d.prev_int[8] ),
    .Y(_11346_));
 sky130_fd_sc_hd__nand2_1 _19449_ (.A(_11345_),
    .B(_11346_),
    .Y(_11347_));
 sky130_fd_sc_hd__or2_1 _19450_ (.A(_11345_),
    .B(_11346_),
    .X(_11348_));
 sky130_fd_sc_hd__a31o_1 _19451_ (.A1(net441),
    .A2(_11347_),
    .A3(_11348_),
    .B1(_11200_),
    .X(_11349_));
 sky130_fd_sc_hd__a22o_1 _19452_ (.A1(\top0.pid_d.curr_int[8] ),
    .A2(_11289_),
    .B1(_11292_),
    .B2(_11349_),
    .X(_11350_));
 sky130_fd_sc_hd__a21o_1 _19453_ (.A1(_10590_),
    .A2(_11341_),
    .B1(_11350_),
    .X(_00334_));
 sky130_fd_sc_hd__inv_2 _19454_ (.A(\top0.pid_d.prev_int[8] ),
    .Y(_11351_));
 sky130_fd_sc_hd__a21o_1 _19455_ (.A1(_11351_),
    .A2(_11345_),
    .B1(_10594_),
    .X(_11352_));
 sky130_fd_sc_hd__o21a_1 _19456_ (.A1(_11351_),
    .A2(_11345_),
    .B1(_11352_),
    .X(_11353_));
 sky130_fd_sc_hd__xor2_1 _19457_ (.A(\top0.pid_d.curr_int[9] ),
    .B(\top0.pid_d.prev_int[9] ),
    .X(_11354_));
 sky130_fd_sc_hd__xnor2_1 _19458_ (.A(_11353_),
    .B(_11354_),
    .Y(_11355_));
 sky130_fd_sc_hd__a221o_1 _19459_ (.A1(net431),
    .A2(_10679_),
    .B1(_11355_),
    .B2(net441),
    .C1(_11209_),
    .X(_11356_));
 sky130_fd_sc_hd__a22o_1 _19460_ (.A1(\top0.pid_d.curr_int[9] ),
    .A2(_11290_),
    .B1(_11293_),
    .B2(_11356_),
    .X(_00335_));
 sky130_fd_sc_hd__inv_2 _19461_ (.A(\top0.pid_d.prev_int[9] ),
    .Y(_11357_));
 sky130_fd_sc_hd__a21o_1 _19462_ (.A1(_11357_),
    .A2(_11353_),
    .B1(_10756_),
    .X(_11358_));
 sky130_fd_sc_hd__o21a_1 _19463_ (.A1(_11357_),
    .A2(_11353_),
    .B1(_11358_),
    .X(_11359_));
 sky130_fd_sc_hd__xnor2_1 _19464_ (.A(\top0.pid_d.curr_int[10] ),
    .B(\top0.pid_d.prev_int[10] ),
    .Y(_11360_));
 sky130_fd_sc_hd__nand2_1 _19465_ (.A(_11359_),
    .B(_11360_),
    .Y(_11361_));
 sky130_fd_sc_hd__or2_1 _19466_ (.A(_11359_),
    .B(_11360_),
    .X(_11362_));
 sky130_fd_sc_hd__a31o_1 _19467_ (.A1(net441),
    .A2(_11361_),
    .A3(_11362_),
    .B1(_11220_),
    .X(_11363_));
 sky130_fd_sc_hd__inv_2 _19468_ (.A(_11289_),
    .Y(_11364_));
 sky130_fd_sc_hd__nor2_1 _19469_ (.A(_10834_),
    .B(_11364_),
    .Y(_11365_));
 sky130_fd_sc_hd__a221o_1 _19470_ (.A1(_10754_),
    .A2(_11341_),
    .B1(_11363_),
    .B2(_11292_),
    .C1(_11365_),
    .X(_00336_));
 sky130_fd_sc_hd__inv_2 _19471_ (.A(\top0.pid_d.prev_int[10] ),
    .Y(_11366_));
 sky130_fd_sc_hd__a21o_1 _19472_ (.A1(_11366_),
    .A2(_11359_),
    .B1(_10834_),
    .X(_11367_));
 sky130_fd_sc_hd__o21a_1 _19473_ (.A1(_11366_),
    .A2(_11359_),
    .B1(_11367_),
    .X(_11368_));
 sky130_fd_sc_hd__xnor2_1 _19474_ (.A(\top0.pid_d.curr_int[11] ),
    .B(\top0.pid_d.prev_int[11] ),
    .Y(_11369_));
 sky130_fd_sc_hd__nand2_1 _19475_ (.A(_11368_),
    .B(_11369_),
    .Y(_11370_));
 sky130_fd_sc_hd__or2_1 _19476_ (.A(_11368_),
    .B(_11369_),
    .X(_11371_));
 sky130_fd_sc_hd__a31o_1 _19477_ (.A1(net441),
    .A2(_11370_),
    .A3(_11371_),
    .B1(_11231_),
    .X(_11372_));
 sky130_fd_sc_hd__and2_1 _19478_ (.A(_10831_),
    .B(_11341_),
    .X(_11373_));
 sky130_fd_sc_hd__a221o_1 _19479_ (.A1(\top0.pid_d.curr_int[11] ),
    .A2(_11290_),
    .B1(_11293_),
    .B2(_11372_),
    .C1(_11373_),
    .X(_00337_));
 sky130_fd_sc_hd__a21oi_1 _19480_ (.A1(_10828_),
    .A2(_10923_),
    .B1(_10924_),
    .Y(_11374_));
 sky130_fd_sc_hd__xnor2_1 _19481_ (.A(_10905_),
    .B(_11374_),
    .Y(_11375_));
 sky130_fd_sc_hd__xor2_1 _19482_ (.A(\top0.pid_d.curr_int[12] ),
    .B(\top0.pid_d.prev_int[12] ),
    .X(_11376_));
 sky130_fd_sc_hd__nand2_1 _19483_ (.A(\top0.pid_d.curr_int[11] ),
    .B(\top0.pid_d.prev_int[11] ),
    .Y(_11377_));
 sky130_fd_sc_hd__nor2_1 _19484_ (.A(\top0.pid_d.curr_int[11] ),
    .B(\top0.pid_d.prev_int[11] ),
    .Y(_11378_));
 sky130_fd_sc_hd__a21o_1 _19485_ (.A1(_11368_),
    .A2(_11377_),
    .B1(_11378_),
    .X(_11379_));
 sky130_fd_sc_hd__xnor2_1 _19486_ (.A(_11376_),
    .B(_11379_),
    .Y(_11380_));
 sky130_fd_sc_hd__a22o_1 _19487_ (.A1(net435),
    .A2(_11240_),
    .B1(_11380_),
    .B2(net441),
    .X(_11381_));
 sky130_fd_sc_hd__a22o_1 _19488_ (.A1(\top0.pid_d.curr_int[12] ),
    .A2(_11289_),
    .B1(_11292_),
    .B2(_11381_),
    .X(_11382_));
 sky130_fd_sc_hd__a21o_1 _19489_ (.A1(_11341_),
    .A2(_11375_),
    .B1(_11382_),
    .X(_00338_));
 sky130_fd_sc_hd__a21bo_1 _19490_ (.A1(\top0.pid_d.curr_int[12] ),
    .A2(\top0.pid_d.prev_int[12] ),
    .B1_N(_11379_),
    .X(_11383_));
 sky130_fd_sc_hd__o21a_1 _19491_ (.A1(\top0.pid_d.curr_int[12] ),
    .A2(\top0.pid_d.prev_int[12] ),
    .B1(_11383_),
    .X(_11384_));
 sky130_fd_sc_hd__xnor2_1 _19492_ (.A(\top0.pid_d.curr_int[13] ),
    .B(\top0.pid_d.prev_int[13] ),
    .Y(_11385_));
 sky130_fd_sc_hd__xnor2_1 _19493_ (.A(_11384_),
    .B(_11385_),
    .Y(_11386_));
 sky130_fd_sc_hd__nand2_1 _19494_ (.A(net441),
    .B(_11386_),
    .Y(_11387_));
 sky130_fd_sc_hd__or2_1 _19495_ (.A(_11289_),
    .B(_11291_),
    .X(_11388_));
 sky130_fd_sc_hd__a21oi_1 _19496_ (.A1(_11252_),
    .A2(_11387_),
    .B1(_11388_),
    .Y(_11389_));
 sky130_fd_sc_hd__a221o_1 _19497_ (.A1(\top0.pid_d.curr_int[13] ),
    .A2(_11289_),
    .B1(_11341_),
    .B2(_10985_),
    .C1(_11389_),
    .X(_00339_));
 sky130_fd_sc_hd__xnor2_1 _19498_ (.A(\top0.pid_d.curr_int[14] ),
    .B(\top0.pid_d.prev_int[14] ),
    .Y(_11390_));
 sky130_fd_sc_hd__or2_1 _19499_ (.A(\top0.pid_d.curr_int[13] ),
    .B(\top0.pid_d.prev_int[13] ),
    .X(_11391_));
 sky130_fd_sc_hd__and2_1 _19500_ (.A(\top0.pid_d.curr_int[13] ),
    .B(\top0.pid_d.prev_int[13] ),
    .X(_11392_));
 sky130_fd_sc_hd__a21o_1 _19501_ (.A1(_11384_),
    .A2(_11391_),
    .B1(_11392_),
    .X(_11393_));
 sky130_fd_sc_hd__xnor2_1 _19502_ (.A(_11390_),
    .B(_11393_),
    .Y(_11394_));
 sky130_fd_sc_hd__nand2_1 _19503_ (.A(net441),
    .B(_11394_),
    .Y(_11395_));
 sky130_fd_sc_hd__a21oi_1 _19504_ (.A1(_11261_),
    .A2(_11395_),
    .B1(_11388_),
    .Y(_11396_));
 sky130_fd_sc_hd__a221o_1 _19505_ (.A1(\top0.pid_d.curr_int[14] ),
    .A2(_11289_),
    .B1(_11341_),
    .B2(_11031_),
    .C1(_11396_),
    .X(_00340_));
 sky130_fd_sc_hd__o21a_1 _19506_ (.A1(_10993_),
    .A2(_11027_),
    .B1(_11077_),
    .X(_11397_));
 sky130_fd_sc_hd__o21a_1 _19507_ (.A1(_11037_),
    .A2(_11397_),
    .B1(_11080_),
    .X(_11398_));
 sky130_fd_sc_hd__or2_1 _19508_ (.A(\top0.pid_d.curr_int[14] ),
    .B(\top0.pid_d.prev_int[14] ),
    .X(_11399_));
 sky130_fd_sc_hd__a21o_1 _19509_ (.A1(\top0.pid_d.curr_int[14] ),
    .A2(\top0.pid_d.prev_int[14] ),
    .B1(_11393_),
    .X(_11400_));
 sky130_fd_sc_hd__xor2_1 _19510_ (.A(\top0.pid_d.curr_int[15] ),
    .B(\top0.pid_d.prev_int[15] ),
    .X(_11401_));
 sky130_fd_sc_hd__a21o_1 _19511_ (.A1(_11399_),
    .A2(_11400_),
    .B1(_11401_),
    .X(_11402_));
 sky130_fd_sc_hd__nand3_1 _19512_ (.A(_11401_),
    .B(_11399_),
    .C(_11400_),
    .Y(_11403_));
 sky130_fd_sc_hd__a32o_1 _19513_ (.A1(net441),
    .A2(_11402_),
    .A3(_11403_),
    .B1(net435),
    .B2(_11268_),
    .X(_11404_));
 sky130_fd_sc_hd__mux2_1 _19514_ (.A0(_11028_),
    .A1(_11029_),
    .S(_11077_),
    .X(_11405_));
 sky130_fd_sc_hd__a22o_1 _19515_ (.A1(\top0.pid_d.curr_int[15] ),
    .A2(_11289_),
    .B1(_11341_),
    .B2(_11405_),
    .X(_11406_));
 sky130_fd_sc_hd__a221o_1 _19516_ (.A1(_11341_),
    .A2(_11398_),
    .B1(_11404_),
    .B2(_11292_),
    .C1(_11406_),
    .X(_00341_));
 sky130_fd_sc_hd__inv_2 _19517_ (.A(net303),
    .Y(_11407_));
 sky130_fd_sc_hd__buf_4 _19518_ (.A(_11407_),
    .X(_11408_));
 sky130_fd_sc_hd__inv_2 _19519_ (.A(net196),
    .Y(_11409_));
 sky130_fd_sc_hd__inv_2 _19520_ (.A(net201),
    .Y(_11410_));
 sky130_fd_sc_hd__nor2_1 _19521_ (.A(net183),
    .B(net189),
    .Y(_11411_));
 sky130_fd_sc_hd__and3_1 _19522_ (.A(_11409_),
    .B(_11410_),
    .C(_11411_),
    .X(_11412_));
 sky130_fd_sc_hd__buf_2 _19523_ (.A(_11412_),
    .X(_11413_));
 sky130_fd_sc_hd__mux2_1 _19524_ (.A0(net83),
    .A1(net88),
    .S(_11413_),
    .X(_11414_));
 sky130_fd_sc_hd__mux4_2 _19525_ (.A0(net108),
    .A1(net103),
    .A2(net98),
    .A3(net94),
    .S0(net199),
    .S1(net193),
    .X(_11415_));
 sky130_fd_sc_hd__mux4_1 _19526_ (.A0(net123),
    .A1(net120),
    .A2(net1031),
    .A3(net113),
    .S0(net197),
    .S1(net191),
    .X(_11416_));
 sky130_fd_sc_hd__mux4_1 _19527_ (.A0(net144),
    .A1(net138),
    .A2(net133),
    .A3(net128),
    .S0(net197),
    .S1(net191),
    .X(_11417_));
 sky130_fd_sc_hd__mux4_1 _19528_ (.A0(net165),
    .A1(net160),
    .A2(net157),
    .A3(\top0.cordic0.vec[1][3] ),
    .S0(net197),
    .S1(net191),
    .X(_11418_));
 sky130_fd_sc_hd__inv_2 _19529_ (.A(net187),
    .Y(_11419_));
 sky130_fd_sc_hd__inv_2 _19530_ (.A(net182),
    .Y(_11420_));
 sky130_fd_sc_hd__mux4_1 _19531_ (.A0(_11415_),
    .A1(_11416_),
    .A2(_11417_),
    .A3(_11418_),
    .S0(_11419_),
    .S1(_11420_),
    .X(_11421_));
 sky130_fd_sc_hd__inv_2 _19532_ (.A(net179),
    .Y(_11422_));
 sky130_fd_sc_hd__mux2_1 _19533_ (.A0(_11414_),
    .A1(_11421_),
    .S(_11422_),
    .X(_11423_));
 sky130_fd_sc_hd__clkbuf_4 _19534_ (.A(_11423_),
    .X(_11424_));
 sky130_fd_sc_hd__clkbuf_4 _19535_ (.A(_11422_),
    .X(_11425_));
 sky130_fd_sc_hd__buf_4 _19536_ (.A(_11425_),
    .X(_11426_));
 sky130_fd_sc_hd__or2_2 _19537_ (.A(net194),
    .B(net203),
    .X(_11427_));
 sky130_fd_sc_hd__or3_2 _19538_ (.A(net186),
    .B(net190),
    .C(_11427_),
    .X(_11428_));
 sky130_fd_sc_hd__nor2_1 _19539_ (.A(_11426_),
    .B(_11428_),
    .Y(_11429_));
 sky130_fd_sc_hd__clkbuf_4 _19540_ (.A(_11429_),
    .X(_11430_));
 sky130_fd_sc_hd__buf_4 _19541_ (.A(_11430_),
    .X(_11431_));
 sky130_fd_sc_hd__o21ai_1 _19542_ (.A1(_11424_),
    .A2(_11431_),
    .B1(net174),
    .Y(_11432_));
 sky130_fd_sc_hd__inv_2 _19543_ (.A(net176),
    .Y(_11433_));
 sky130_fd_sc_hd__nor2_1 _19544_ (.A(_11433_),
    .B(_11430_),
    .Y(_11434_));
 sky130_fd_sc_hd__clkbuf_4 _19545_ (.A(_11434_),
    .X(_11435_));
 sky130_fd_sc_hd__and3_1 _19546_ (.A(net306),
    .B(_11424_),
    .C(_11435_),
    .X(_11436_));
 sky130_fd_sc_hd__a21oi_1 _19547_ (.A1(_11408_),
    .A2(_11432_),
    .B1(_11436_),
    .Y(_00342_));
 sky130_fd_sc_hd__inv_2 _19548_ (.A(net299),
    .Y(_11437_));
 sky130_fd_sc_hd__buf_4 _19549_ (.A(_11437_),
    .X(_11438_));
 sky130_fd_sc_hd__clkbuf_2 _19550_ (.A(_11430_),
    .X(_11439_));
 sky130_fd_sc_hd__mux4_2 _19551_ (.A0(net103),
    .A1(net98),
    .A2(net94),
    .A3(net88),
    .S0(net199),
    .S1(\top0.cordic0.gm0.iter[1] ),
    .X(_11440_));
 sky130_fd_sc_hd__mux4_1 _19552_ (.A0(net121),
    .A1(net1031),
    .A2(net113),
    .A3(net108),
    .S0(net198),
    .S1(net191),
    .X(_11441_));
 sky130_fd_sc_hd__mux2_1 _19553_ (.A0(_11440_),
    .A1(_11441_),
    .S(_11419_),
    .X(_11442_));
 sky130_fd_sc_hd__or3_2 _19554_ (.A(_11420_),
    .B(net179),
    .C(_11442_),
    .X(_11443_));
 sky130_fd_sc_hd__inv_2 _19555_ (.A(net81),
    .Y(_11444_));
 sky130_fd_sc_hd__nand2_2 _19556_ (.A(net179),
    .B(_11444_),
    .Y(_11445_));
 sky130_fd_sc_hd__mux4_1 _19557_ (.A0(net138),
    .A1(net133),
    .A2(net129),
    .A3(net125),
    .S0(net197),
    .S1(net191),
    .X(_11446_));
 sky130_fd_sc_hd__or2_1 _19558_ (.A(net182),
    .B(net180),
    .X(_11447_));
 sky130_fd_sc_hd__buf_2 _19559_ (.A(_11447_),
    .X(_11448_));
 sky130_fd_sc_hd__a21o_1 _19560_ (.A1(net188),
    .A2(_11446_),
    .B1(_11448_),
    .X(_11449_));
 sky130_fd_sc_hd__mux4_2 _19561_ (.A0(net160),
    .A1(net156),
    .A2(net150),
    .A3(net144),
    .S0(net197),
    .S1(net191),
    .X(_11450_));
 sky130_fd_sc_hd__nor2_2 _19562_ (.A(net188),
    .B(_11448_),
    .Y(_11451_));
 sky130_fd_sc_hd__a32oi_4 _19563_ (.A1(_11443_),
    .A2(_11445_),
    .A3(_11449_),
    .B1(_11450_),
    .B2(_11451_),
    .Y(_11452_));
 sky130_fd_sc_hd__and2b_1 _19564_ (.A_N(\top0.cordic0.slte0.opB[4] ),
    .B(\top0.cordic0.slte0.opA[4] ),
    .X(_11453_));
 sky130_fd_sc_hd__a21bo_1 _19565_ (.A1(\top0.cordic0.slte0.opA[5] ),
    .A2(_11453_),
    .B1_N(\top0.cordic0.slte0.opB[5] ),
    .X(_11454_));
 sky130_fd_sc_hd__o21ai_1 _19566_ (.A1(\top0.cordic0.slte0.opA[5] ),
    .A2(_11453_),
    .B1(_11454_),
    .Y(_11455_));
 sky130_fd_sc_hd__or2b_1 _19567_ (.A(\top0.cordic0.slte0.opA[2] ),
    .B_N(\top0.cordic0.slte0.opB[2] ),
    .X(_11456_));
 sky130_fd_sc_hd__nand2_1 _19568_ (.A(\top0.cordic0.slte0.opA[3] ),
    .B(_11456_),
    .Y(_11457_));
 sky130_fd_sc_hd__nor2_1 _19569_ (.A(\top0.cordic0.slte0.opA[3] ),
    .B(_11456_),
    .Y(_11458_));
 sky130_fd_sc_hd__or2_1 _19570_ (.A(\top0.cordic0.slte0.opB[5] ),
    .B(\top0.cordic0.slte0.opA[5] ),
    .X(_11459_));
 sky130_fd_sc_hd__nand2_1 _19571_ (.A(\top0.cordic0.slte0.opB[5] ),
    .B(\top0.cordic0.slte0.opA[5] ),
    .Y(_11460_));
 sky130_fd_sc_hd__and2b_1 _19572_ (.A_N(\top0.cordic0.slte0.opA[4] ),
    .B(\top0.cordic0.slte0.opB[4] ),
    .X(_11461_));
 sky130_fd_sc_hd__a211o_1 _19573_ (.A1(_11459_),
    .A2(_11460_),
    .B1(_11453_),
    .C1(_11461_),
    .X(_11462_));
 sky130_fd_sc_hd__a211o_1 _19574_ (.A1(\top0.cordic0.slte0.opB[3] ),
    .A2(_11457_),
    .B1(_11458_),
    .C1(_11462_),
    .X(_11463_));
 sky130_fd_sc_hd__xor2_1 _19575_ (.A(\top0.cordic0.slte0.opB[13] ),
    .B(\top0.cordic0.slte0.opA[13] ),
    .X(_11464_));
 sky130_fd_sc_hd__nor2b_1 _19576_ (.A(\top0.cordic0.slte0.opB[12] ),
    .B_N(\top0.cordic0.slte0.opA[12] ),
    .Y(_11465_));
 sky130_fd_sc_hd__and2b_1 _19577_ (.A_N(\top0.cordic0.slte0.opA[12] ),
    .B(\top0.cordic0.slte0.opB[12] ),
    .X(_11466_));
 sky130_fd_sc_hd__and2b_1 _19578_ (.A_N(\top0.cordic0.slte0.opA[11] ),
    .B(\top0.cordic0.slte0.opB[11] ),
    .X(_11467_));
 sky130_fd_sc_hd__or4_1 _19579_ (.A(_11464_),
    .B(_11465_),
    .C(_11466_),
    .D(_11467_),
    .X(_11468_));
 sky130_fd_sc_hd__and2b_1 _19580_ (.A_N(\top0.cordic0.slte0.opB[14] ),
    .B(\top0.cordic0.slte0.opA[14] ),
    .X(_11469_));
 sky130_fd_sc_hd__and2b_1 _19581_ (.A_N(\top0.cordic0.slte0.opA[14] ),
    .B(\top0.cordic0.slte0.opB[14] ),
    .X(_11470_));
 sky130_fd_sc_hd__and2b_1 _19582_ (.A_N(\top0.cordic0.slte0.opB[15] ),
    .B(\top0.cordic0.slte0.opA[15] ),
    .X(_11471_));
 sky130_fd_sc_hd__and2b_1 _19583_ (.A_N(\top0.cordic0.slte0.opA[15] ),
    .B(\top0.cordic0.slte0.opB[15] ),
    .X(_11472_));
 sky130_fd_sc_hd__or4_1 _19584_ (.A(_11469_),
    .B(_11470_),
    .C(_11471_),
    .D(_11472_),
    .X(_11473_));
 sky130_fd_sc_hd__xor2_1 _19585_ (.A(\top0.cordic0.slte0.opA[10] ),
    .B(\top0.cordic0.slte0.opB[10] ),
    .X(_11474_));
 sky130_fd_sc_hd__and2b_1 _19586_ (.A_N(\top0.cordic0.slte0.opB[11] ),
    .B(\top0.cordic0.slte0.opA[11] ),
    .X(_11475_));
 sky130_fd_sc_hd__nor2_1 _19587_ (.A(\top0.cordic0.slte0.opA[16] ),
    .B(\top0.cordic0.slte0.opA[17] ),
    .Y(_11476_));
 sky130_fd_sc_hd__or3b_1 _19588_ (.A(_11474_),
    .B(_11475_),
    .C_N(_11476_),
    .X(_11477_));
 sky130_fd_sc_hd__xor2_1 _19589_ (.A(\top0.cordic0.slte0.opB[7] ),
    .B(\top0.cordic0.slte0.opA[7] ),
    .X(_11478_));
 sky130_fd_sc_hd__xor2_1 _19590_ (.A(\top0.cordic0.slte0.opB[8] ),
    .B(\top0.cordic0.slte0.opA[8] ),
    .X(_11479_));
 sky130_fd_sc_hd__xor2_1 _19591_ (.A(\top0.cordic0.slte0.opB[9] ),
    .B(\top0.cordic0.slte0.opA[9] ),
    .X(_11480_));
 sky130_fd_sc_hd__xor2_1 _19592_ (.A(\top0.cordic0.slte0.opA[6] ),
    .B(\top0.cordic0.slte0.opB[6] ),
    .X(_11481_));
 sky130_fd_sc_hd__or4_1 _19593_ (.A(_11478_),
    .B(_11479_),
    .C(_11480_),
    .D(_11481_),
    .X(_11482_));
 sky130_fd_sc_hd__or4_4 _19594_ (.A(_11468_),
    .B(_11473_),
    .C(_11477_),
    .D(_11482_),
    .X(_11483_));
 sky130_fd_sc_hd__a21o_4 _19595_ (.A1(_11455_),
    .A2(_11463_),
    .B1(_11483_),
    .X(_11484_));
 sky130_fd_sc_hd__inv_2 _19596_ (.A(\top0.cordic0.slte0.opB[8] ),
    .Y(_11485_));
 sky130_fd_sc_hd__or2_1 _19597_ (.A(_11485_),
    .B(\top0.cordic0.slte0.opA[8] ),
    .X(_11486_));
 sky130_fd_sc_hd__and2b_1 _19598_ (.A_N(\top0.cordic0.slte0.opB[6] ),
    .B(\top0.cordic0.slte0.opA[6] ),
    .X(_11487_));
 sky130_fd_sc_hd__a21bo_1 _19599_ (.A1(\top0.cordic0.slte0.opA[7] ),
    .A2(_11487_),
    .B1_N(\top0.cordic0.slte0.opB[7] ),
    .X(_11488_));
 sky130_fd_sc_hd__or2_1 _19600_ (.A(\top0.cordic0.slte0.opA[7] ),
    .B(_11487_),
    .X(_11489_));
 sky130_fd_sc_hd__a22o_1 _19601_ (.A1(_11485_),
    .A2(\top0.cordic0.slte0.opA[8] ),
    .B1(_11488_),
    .B2(_11489_),
    .X(_11490_));
 sky130_fd_sc_hd__a21oi_1 _19602_ (.A1(_11486_),
    .A2(_11490_),
    .B1(\top0.cordic0.slte0.opA[9] ),
    .Y(_11491_));
 sky130_fd_sc_hd__or3_1 _19603_ (.A(_11468_),
    .B(_11473_),
    .C(_11477_),
    .X(_11492_));
 sky130_fd_sc_hd__or2_1 _19604_ (.A(\top0.cordic0.slte0.opB[9] ),
    .B(_11492_),
    .X(_11493_));
 sky130_fd_sc_hd__inv_2 _19605_ (.A(\top0.cordic0.slte0.opA[9] ),
    .Y(_11494_));
 sky130_fd_sc_hd__or2_1 _19606_ (.A(_11494_),
    .B(_11492_),
    .X(_11495_));
 sky130_fd_sc_hd__nand2_1 _19607_ (.A(_11486_),
    .B(_11490_),
    .Y(_11496_));
 sky130_fd_sc_hd__a21boi_1 _19608_ (.A1(\top0.cordic0.slte0.opA[13] ),
    .A2(_11465_),
    .B1_N(\top0.cordic0.slte0.opB[13] ),
    .Y(_11497_));
 sky130_fd_sc_hd__nor2_1 _19609_ (.A(\top0.cordic0.slte0.opA[13] ),
    .B(_11465_),
    .Y(_11498_));
 sky130_fd_sc_hd__inv_2 _19610_ (.A(\top0.cordic0.slte0.opB[10] ),
    .Y(_11499_));
 sky130_fd_sc_hd__a21oi_1 _19611_ (.A1(\top0.cordic0.slte0.opA[10] ),
    .A2(_11499_),
    .B1(_11475_),
    .Y(_11500_));
 sky130_fd_sc_hd__o22a_1 _19612_ (.A1(_11497_),
    .A2(_11498_),
    .B1(_11500_),
    .B2(_11468_),
    .X(_11501_));
 sky130_fd_sc_hd__nor2_1 _19613_ (.A(_11469_),
    .B(_11471_),
    .Y(_11502_));
 sky130_fd_sc_hd__o221a_1 _19614_ (.A1(_11473_),
    .A2(_11501_),
    .B1(_11502_),
    .B2(_11472_),
    .C1(_11476_),
    .X(_11503_));
 sky130_fd_sc_hd__o221a_4 _19615_ (.A1(_11491_),
    .A2(_11493_),
    .B1(_11495_),
    .B2(_11496_),
    .C1(_11503_),
    .X(_11504_));
 sky130_fd_sc_hd__inv_2 _19616_ (.A(\top0.cordic0.slte0.opB[2] ),
    .Y(_11505_));
 sky130_fd_sc_hd__xor2_1 _19617_ (.A(\top0.cordic0.slte0.opB[3] ),
    .B(\top0.cordic0.slte0.opA[3] ),
    .X(_11506_));
 sky130_fd_sc_hd__or3b_1 _19618_ (.A(\top0.cordic0.slte0.opA[1] ),
    .B(\top0.cordic0.slte0.opA[0] ),
    .C_N(_11456_),
    .X(_11507_));
 sky130_fd_sc_hd__a2111o_1 _19619_ (.A1(\top0.cordic0.slte0.opA[2] ),
    .A2(_11505_),
    .B1(_11462_),
    .C1(_11506_),
    .D1(_11507_),
    .X(_11508_));
 sky130_fd_sc_hd__o21bai_4 _19620_ (.A1(_11483_),
    .A2(_11508_),
    .B1_N(\top0.cordic0.slte0.opA[17] ),
    .Y(_11509_));
 sky130_fd_sc_hd__a21oi_4 _19621_ (.A1(_11484_),
    .A2(_11504_),
    .B1(_11509_),
    .Y(_11510_));
 sky130_fd_sc_hd__buf_6 _19622_ (.A(_11510_),
    .X(_11511_));
 sky130_fd_sc_hd__buf_6 _19623_ (.A(_11511_),
    .X(_11512_));
 sky130_fd_sc_hd__clkbuf_4 _19624_ (.A(_11512_),
    .X(_11513_));
 sky130_fd_sc_hd__buf_2 _19625_ (.A(_11513_),
    .X(_11514_));
 sky130_fd_sc_hd__clkbuf_4 _19626_ (.A(_11514_),
    .X(_11515_));
 sky130_fd_sc_hd__nand2_1 _19627_ (.A(_11408_),
    .B(_11515_),
    .Y(_11516_));
 sky130_fd_sc_hd__a21o_1 _19628_ (.A1(_11484_),
    .A2(_11504_),
    .B1(_11509_),
    .X(_11517_));
 sky130_fd_sc_hd__clkbuf_4 _19629_ (.A(net1016),
    .X(_11518_));
 sky130_fd_sc_hd__buf_4 _19630_ (.A(_11518_),
    .X(_11519_));
 sky130_fd_sc_hd__nand2_1 _19631_ (.A(net306),
    .B(_11519_),
    .Y(_11520_));
 sky130_fd_sc_hd__and3_1 _19632_ (.A(_11424_),
    .B(_11516_),
    .C(_11520_),
    .X(_11521_));
 sky130_fd_sc_hd__xnor2_1 _19633_ (.A(_11452_),
    .B(_11521_),
    .Y(_11522_));
 sky130_fd_sc_hd__o21ai_1 _19634_ (.A1(net1014),
    .A2(_11522_),
    .B1(net174),
    .Y(_11523_));
 sky130_fd_sc_hd__and3_1 _19635_ (.A(net300),
    .B(_11435_),
    .C(_11522_),
    .X(_11524_));
 sky130_fd_sc_hd__a21oi_1 _19636_ (.A1(_11438_),
    .A2(_11523_),
    .B1(_11524_),
    .Y(_00343_));
 sky130_fd_sc_hd__inv_2 _19637_ (.A(net297),
    .Y(_11525_));
 sky130_fd_sc_hd__buf_4 _19638_ (.A(_11430_),
    .X(_11526_));
 sky130_fd_sc_hd__nor2_1 _19639_ (.A(net306),
    .B(net300),
    .Y(_11527_));
 sky130_fd_sc_hd__a32o_1 _19640_ (.A1(_11443_),
    .A2(_11445_),
    .A3(_11449_),
    .B1(_11450_),
    .B2(_11451_),
    .X(_11528_));
 sky130_fd_sc_hd__nand2_1 _19641_ (.A(_11438_),
    .B(_11528_),
    .Y(_11529_));
 sky130_fd_sc_hd__nor2_1 _19642_ (.A(_11424_),
    .B(_11529_),
    .Y(_11530_));
 sky130_fd_sc_hd__a21oi_1 _19643_ (.A1(_11424_),
    .A2(_11527_),
    .B1(_11530_),
    .Y(_11531_));
 sky130_fd_sc_hd__or3b_1 _19644_ (.A(net306),
    .B(_11452_),
    .C_N(_11424_),
    .X(_11532_));
 sky130_fd_sc_hd__a21o_1 _19645_ (.A1(_11529_),
    .A2(_11532_),
    .B1(_11511_),
    .X(_11533_));
 sky130_fd_sc_hd__o2111ai_4 _19646_ (.A1(_11408_),
    .A2(_11438_),
    .B1(_11424_),
    .C1(_11452_),
    .D1(_11511_),
    .Y(_11534_));
 sky130_fd_sc_hd__mux4_2 _19647_ (.A0(net98),
    .A1(net94),
    .A2(net88),
    .A3(net83),
    .S0(net199),
    .S1(net193),
    .X(_11535_));
 sky130_fd_sc_hd__mux4_1 _19648_ (.A0(net116),
    .A1(net111),
    .A2(net108),
    .A3(net103),
    .S0(net199),
    .S1(net193),
    .X(_11536_));
 sky130_fd_sc_hd__mux4_1 _19649_ (.A0(net133),
    .A1(net128),
    .A2(net123),
    .A3(net121),
    .S0(net199),
    .S1(net193),
    .X(_11537_));
 sky130_fd_sc_hd__mux4_1 _19650_ (.A0(net157),
    .A1(net150),
    .A2(net144),
    .A3(net140),
    .S0(net198),
    .S1(net191),
    .X(_11538_));
 sky130_fd_sc_hd__mux4_1 _19651_ (.A0(_11535_),
    .A1(_11536_),
    .A2(_11537_),
    .A3(_11538_),
    .S0(_11419_),
    .S1(_11420_),
    .X(_11539_));
 sky130_fd_sc_hd__mux2_2 _19652_ (.A0(net84),
    .A1(_11539_),
    .S(_11422_),
    .X(_11540_));
 sky130_fd_sc_hd__nor2_1 _19653_ (.A(_11424_),
    .B(_11528_),
    .Y(_11541_));
 sky130_fd_sc_hd__a211o_1 _19654_ (.A1(_11484_),
    .A2(_11504_),
    .B1(_11509_),
    .C1(_11541_),
    .X(_11542_));
 sky130_fd_sc_hd__xor2_2 _19655_ (.A(_11540_),
    .B(_11542_),
    .X(_11543_));
 sky130_fd_sc_hd__a31o_1 _19656_ (.A1(_11531_),
    .A2(_11533_),
    .A3(_11534_),
    .B1(_11543_),
    .X(_11544_));
 sky130_fd_sc_hd__nand4_1 _19657_ (.A(_11543_),
    .B(_11531_),
    .C(_11533_),
    .D(_11534_),
    .Y(_11545_));
 sky130_fd_sc_hd__and2_1 _19658_ (.A(_11544_),
    .B(_11545_),
    .X(_11546_));
 sky130_fd_sc_hd__or2_1 _19659_ (.A(_11526_),
    .B(_11546_),
    .X(_11547_));
 sky130_fd_sc_hd__clkbuf_2 _19660_ (.A(_11434_),
    .X(_11548_));
 sky130_fd_sc_hd__a21oi_1 _19661_ (.A1(net1013),
    .A2(_11546_),
    .B1(_11525_),
    .Y(_11549_));
 sky130_fd_sc_hd__a31o_1 _19662_ (.A1(net174),
    .A2(_11525_),
    .A3(_11547_),
    .B1(_11549_),
    .X(_00344_));
 sky130_fd_sc_hd__inv_2 _19663_ (.A(net291),
    .Y(_11550_));
 sky130_fd_sc_hd__a41o_1 _19664_ (.A1(_11543_),
    .A2(_11531_),
    .A3(_11533_),
    .A4(_11534_),
    .B1(net297),
    .X(_11551_));
 sky130_fd_sc_hd__nand2_1 _19665_ (.A(_11544_),
    .B(_11551_),
    .Y(_11552_));
 sky130_fd_sc_hd__mux2_1 _19666_ (.A0(net94),
    .A1(net88),
    .S(net200),
    .X(_11553_));
 sky130_fd_sc_hd__mux2_1 _19667_ (.A0(net111),
    .A1(net108),
    .S(net199),
    .X(_11554_));
 sky130_fd_sc_hd__and2b_1 _19668_ (.A_N(net199),
    .B(net84),
    .X(_11555_));
 sky130_fd_sc_hd__mux2_1 _19669_ (.A0(net103),
    .A1(net98),
    .S(net200),
    .X(_11556_));
 sky130_fd_sc_hd__mux4_1 _19670_ (.A0(_11553_),
    .A1(_11554_),
    .A2(_11555_),
    .A3(_11556_),
    .S0(_11419_),
    .S1(net193),
    .X(_11557_));
 sky130_fd_sc_hd__and3_1 _19671_ (.A(\top0.cordic0.gm0.iter[1] ),
    .B(net200),
    .C(net187),
    .X(_11558_));
 sky130_fd_sc_hd__a22o_1 _19672_ (.A1(_11422_),
    .A2(_11557_),
    .B1(_11558_),
    .B2(net84),
    .X(_11559_));
 sky130_fd_sc_hd__nor2_4 _19673_ (.A(net186),
    .B(net180),
    .Y(_11560_));
 sky130_fd_sc_hd__mux4_1 _19674_ (.A0(net150),
    .A1(net144),
    .A2(net138),
    .A3(net133),
    .S0(net199),
    .S1(net193),
    .X(_11561_));
 sky130_fd_sc_hd__mux4_1 _19675_ (.A0(net128),
    .A1(net123),
    .A2(net121),
    .A3(net116),
    .S0(net199),
    .S1(net193),
    .X(_11562_));
 sky130_fd_sc_hd__mux2_1 _19676_ (.A0(_11561_),
    .A1(_11562_),
    .S(net187),
    .X(_11563_));
 sky130_fd_sc_hd__a22o_1 _19677_ (.A1(net179),
    .A2(net84),
    .B1(_11560_),
    .B2(_11563_),
    .X(_11564_));
 sky130_fd_sc_hd__a21oi_2 _19678_ (.A1(net182),
    .A2(_11559_),
    .B1(_11564_),
    .Y(_11565_));
 sky130_fd_sc_hd__o31ai_2 _19679_ (.A1(_11424_),
    .A2(_11528_),
    .A3(_11540_),
    .B1(_11512_),
    .Y(_11566_));
 sky130_fd_sc_hd__xnor2_2 _19680_ (.A(_11565_),
    .B(_11566_),
    .Y(_11567_));
 sky130_fd_sc_hd__xnor2_1 _19681_ (.A(_11552_),
    .B(_11567_),
    .Y(_11568_));
 sky130_fd_sc_hd__o21ai_1 _19682_ (.A1(net1014),
    .A2(_11568_),
    .B1(net174),
    .Y(_11569_));
 sky130_fd_sc_hd__and3_1 _19683_ (.A(net291),
    .B(_11435_),
    .C(_11568_),
    .X(_11570_));
 sky130_fd_sc_hd__a21oi_1 _19684_ (.A1(_11550_),
    .A2(_11569_),
    .B1(_11570_),
    .Y(_00345_));
 sky130_fd_sc_hd__inv_2 _19685_ (.A(net286),
    .Y(_11571_));
 sky130_fd_sc_hd__clkbuf_4 _19686_ (.A(_11419_),
    .X(_11572_));
 sky130_fd_sc_hd__clkbuf_4 _19687_ (.A(_11572_),
    .X(_11573_));
 sky130_fd_sc_hd__nor2_1 _19688_ (.A(net194),
    .B(_11572_),
    .Y(_11574_));
 sky130_fd_sc_hd__mux2_1 _19689_ (.A0(net88),
    .A1(net83),
    .S(net203),
    .X(_11575_));
 sky130_fd_sc_hd__clkbuf_4 _19690_ (.A(_11420_),
    .X(_11576_));
 sky130_fd_sc_hd__a221o_1 _19691_ (.A1(_11573_),
    .A2(_11415_),
    .B1(_11574_),
    .B2(_11575_),
    .C1(_11576_),
    .X(_11577_));
 sky130_fd_sc_hd__mux2_1 _19692_ (.A0(_11416_),
    .A1(_11417_),
    .S(_11572_),
    .X(_11578_));
 sky130_fd_sc_hd__or2_1 _19693_ (.A(net182),
    .B(_11578_),
    .X(_11579_));
 sky130_fd_sc_hd__a31o_1 _19694_ (.A1(net193),
    .A2(net182),
    .A3(net187),
    .B1(net179),
    .X(_11580_));
 sky130_fd_sc_hd__a32o_2 _19695_ (.A1(_11425_),
    .A2(_11577_),
    .A3(_11579_),
    .B1(_11580_),
    .B2(net82),
    .X(_11581_));
 sky130_fd_sc_hd__or4b_2 _19696_ (.A(_11424_),
    .B(_11528_),
    .C(_11540_),
    .D_N(_11565_),
    .X(_11582_));
 sky130_fd_sc_hd__nand2_2 _19697_ (.A(_11511_),
    .B(_11582_),
    .Y(_11583_));
 sky130_fd_sc_hd__xor2_4 _19698_ (.A(_11581_),
    .B(_11583_),
    .X(_11584_));
 sky130_fd_sc_hd__inv_2 _19699_ (.A(_11584_),
    .Y(_11585_));
 sky130_fd_sc_hd__nor2_1 _19700_ (.A(net291),
    .B(_11567_),
    .Y(_11586_));
 sky130_fd_sc_hd__a22oi_2 _19701_ (.A1(_11544_),
    .A2(_11551_),
    .B1(_11567_),
    .B2(net292),
    .Y(_11587_));
 sky130_fd_sc_hd__nor2_1 _19702_ (.A(_11586_),
    .B(_11587_),
    .Y(_11588_));
 sky130_fd_sc_hd__xnor2_1 _19703_ (.A(_11585_),
    .B(_11588_),
    .Y(_11589_));
 sky130_fd_sc_hd__or2_1 _19704_ (.A(_11526_),
    .B(_11589_),
    .X(_11590_));
 sky130_fd_sc_hd__a21oi_1 _19705_ (.A1(net1013),
    .A2(_11589_),
    .B1(_11571_),
    .Y(_11591_));
 sky130_fd_sc_hd__a31o_1 _19706_ (.A1(net174),
    .A2(_11571_),
    .A3(_11590_),
    .B1(_11591_),
    .X(_00346_));
 sky130_fd_sc_hd__inv_2 _19707_ (.A(net277),
    .Y(_11592_));
 sky130_fd_sc_hd__clkbuf_4 _19708_ (.A(_11592_),
    .X(_11593_));
 sky130_fd_sc_hd__a31o_1 _19709_ (.A1(net182),
    .A2(net188),
    .A3(_11427_),
    .B1(net179),
    .X(_11594_));
 sky130_fd_sc_hd__nand2_1 _19710_ (.A(net188),
    .B(net82),
    .Y(_11595_));
 sky130_fd_sc_hd__o2bb2a_1 _19711_ (.A1_N(_11572_),
    .A2_N(_11440_),
    .B1(_11595_),
    .B2(_11427_),
    .X(_11596_));
 sky130_fd_sc_hd__nand2_1 _19712_ (.A(net188),
    .B(_11441_),
    .Y(_11597_));
 sky130_fd_sc_hd__mux2_1 _19713_ (.A0(_11596_),
    .A1(_11597_),
    .S(_11576_),
    .X(_11598_));
 sky130_fd_sc_hd__nor2_1 _19714_ (.A(net179),
    .B(_11598_),
    .Y(_11599_));
 sky130_fd_sc_hd__a221o_1 _19715_ (.A1(_11451_),
    .A2(_11446_),
    .B1(_11594_),
    .B2(net84),
    .C1(_11599_),
    .X(_11600_));
 sky130_fd_sc_hd__o21a_1 _19716_ (.A1(_11581_),
    .A2(_11582_),
    .B1(_11512_),
    .X(_11601_));
 sky130_fd_sc_hd__xnor2_2 _19717_ (.A(_11600_),
    .B(_11601_),
    .Y(_11602_));
 sky130_fd_sc_hd__o31a_1 _19718_ (.A1(_11585_),
    .A2(_11586_),
    .A3(_11587_),
    .B1(_11571_),
    .X(_11603_));
 sky130_fd_sc_hd__o21bai_2 _19719_ (.A1(_11584_),
    .A2(_11588_),
    .B1_N(_11603_),
    .Y(_11604_));
 sky130_fd_sc_hd__xnor2_1 _19720_ (.A(_11602_),
    .B(_11604_),
    .Y(_11605_));
 sky130_fd_sc_hd__or2_1 _19721_ (.A(_11430_),
    .B(_11605_),
    .X(_11606_));
 sky130_fd_sc_hd__a21oi_1 _19722_ (.A1(net1013),
    .A2(_11605_),
    .B1(_11593_),
    .Y(_11607_));
 sky130_fd_sc_hd__a31o_1 _19723_ (.A1(net175),
    .A2(_11593_),
    .A3(_11606_),
    .B1(_11607_),
    .X(_00347_));
 sky130_fd_sc_hd__inv_6 _19724_ (.A(net273),
    .Y(_11608_));
 sky130_fd_sc_hd__nor2_1 _19725_ (.A(net277),
    .B(_11602_),
    .Y(_11609_));
 sky130_fd_sc_hd__and2_1 _19726_ (.A(net277),
    .B(_11602_),
    .X(_11610_));
 sky130_fd_sc_hd__inv_2 _19727_ (.A(_11610_),
    .Y(_11611_));
 sky130_fd_sc_hd__clkbuf_4 _19728_ (.A(_11576_),
    .X(_11612_));
 sky130_fd_sc_hd__or2_1 _19729_ (.A(net188),
    .B(net179),
    .X(_11613_));
 sky130_fd_sc_hd__o22a_1 _19730_ (.A1(_11573_),
    .A2(net82),
    .B1(_11535_),
    .B2(_11613_),
    .X(_11614_));
 sky130_fd_sc_hd__mux2_1 _19731_ (.A0(_11536_),
    .A1(_11537_),
    .S(_11573_),
    .X(_11615_));
 sky130_fd_sc_hd__o221a_2 _19732_ (.A1(_11612_),
    .A2(_11614_),
    .B1(_11615_),
    .B2(_11448_),
    .C1(_11445_),
    .X(_11616_));
 sky130_fd_sc_hd__or3_1 _19733_ (.A(_11581_),
    .B(_11582_),
    .C(_11600_),
    .X(_11617_));
 sky130_fd_sc_hd__nand2_2 _19734_ (.A(_11512_),
    .B(_11617_),
    .Y(_11618_));
 sky130_fd_sc_hd__xor2_4 _19735_ (.A(_11616_),
    .B(_11618_),
    .X(_11619_));
 sky130_fd_sc_hd__inv_2 _19736_ (.A(_11619_),
    .Y(_11620_));
 sky130_fd_sc_hd__o211ai_4 _19737_ (.A1(_11604_),
    .A2(_11609_),
    .B1(_11611_),
    .C1(_11620_),
    .Y(_11621_));
 sky130_fd_sc_hd__nand2_1 _19738_ (.A(_11584_),
    .B(_11619_),
    .Y(_11622_));
 sky130_fd_sc_hd__nand2_1 _19739_ (.A(net286),
    .B(_11619_),
    .Y(_11623_));
 sky130_fd_sc_hd__a2111o_1 _19740_ (.A1(_11622_),
    .A2(_11623_),
    .B1(_11586_),
    .C1(_11587_),
    .D1(_11609_),
    .X(_11624_));
 sky130_fd_sc_hd__o2111a_1 _19741_ (.A1(net277),
    .A2(_11602_),
    .B1(_11619_),
    .C1(_11584_),
    .D1(net286),
    .X(_11625_));
 sky130_fd_sc_hd__a21oi_1 _19742_ (.A1(_11619_),
    .A2(_11610_),
    .B1(_11625_),
    .Y(_11626_));
 sky130_fd_sc_hd__a31o_1 _19743_ (.A1(_11621_),
    .A2(_11624_),
    .A3(_11626_),
    .B1(_11526_),
    .X(_11627_));
 sky130_fd_sc_hd__a41oi_1 _19744_ (.A1(_11435_),
    .A2(_11621_),
    .A3(_11624_),
    .A4(_11626_),
    .B1(_11608_),
    .Y(_11628_));
 sky130_fd_sc_hd__a31o_1 _19745_ (.A1(net174),
    .A2(_11608_),
    .A3(_11627_),
    .B1(_11628_),
    .X(_00348_));
 sky130_fd_sc_hd__nand2_1 _19746_ (.A(net194),
    .B(net203),
    .Y(_11629_));
 sky130_fd_sc_hd__a21oi_1 _19747_ (.A1(_11573_),
    .A2(_11629_),
    .B1(_11576_),
    .Y(_11630_));
 sky130_fd_sc_hd__or2_1 _19748_ (.A(net180),
    .B(_11630_),
    .X(_11631_));
 sky130_fd_sc_hd__clkbuf_4 _19749_ (.A(_11409_),
    .X(_11632_));
 sky130_fd_sc_hd__and2b_1 _19750_ (.A_N(net201),
    .B(net194),
    .X(_11633_));
 sky130_fd_sc_hd__a22oi_2 _19751_ (.A1(_11632_),
    .A2(_11553_),
    .B1(_11633_),
    .B2(net83),
    .Y(_11634_));
 sky130_fd_sc_hd__mux4_1 _19752_ (.A0(net120),
    .A1(net116),
    .A2(net103),
    .A3(net98),
    .S0(net200),
    .S1(net187),
    .X(_11635_));
 sky130_fd_sc_hd__mux4_1 _19753_ (.A0(net128),
    .A1(net123),
    .A2(net111),
    .A3(net107),
    .S0(net199),
    .S1(net187),
    .X(_11636_));
 sky130_fd_sc_hd__mux2_1 _19754_ (.A0(_11635_),
    .A1(_11636_),
    .S(_11632_),
    .X(_11637_));
 sky130_fd_sc_hd__nand2_1 _19755_ (.A(_11612_),
    .B(_11637_),
    .Y(_11638_));
 sky130_fd_sc_hd__o31a_1 _19756_ (.A1(_11612_),
    .A2(net187),
    .A3(_11634_),
    .B1(_11638_),
    .X(_11639_));
 sky130_fd_sc_hd__o2bb2a_1 _19757_ (.A1_N(net83),
    .A2_N(_11631_),
    .B1(_11639_),
    .B2(net180),
    .X(_11640_));
 sky130_fd_sc_hd__nor2_1 _19758_ (.A(_11616_),
    .B(_11617_),
    .Y(_11641_));
 sky130_fd_sc_hd__or2_1 _19759_ (.A(_11518_),
    .B(_11641_),
    .X(_11642_));
 sky130_fd_sc_hd__xnor2_2 _19760_ (.A(_11640_),
    .B(_11642_),
    .Y(_11643_));
 sky130_fd_sc_hd__nand2_1 _19761_ (.A(_11624_),
    .B(_11626_),
    .Y(_11644_));
 sky130_fd_sc_hd__a21oi_1 _19762_ (.A1(net272),
    .A2(_11621_),
    .B1(_11644_),
    .Y(_11645_));
 sky130_fd_sc_hd__xor2_1 _19763_ (.A(_11643_),
    .B(_11645_),
    .X(_11646_));
 sky130_fd_sc_hd__nand2_1 _19764_ (.A(net266),
    .B(_11435_),
    .Y(_11647_));
 sky130_fd_sc_hd__nand2_1 _19765_ (.A(net180),
    .B(_11413_),
    .Y(_11648_));
 sky130_fd_sc_hd__clkbuf_4 _19766_ (.A(_11648_),
    .X(_11649_));
 sky130_fd_sc_hd__buf_4 _19767_ (.A(_11649_),
    .X(_11650_));
 sky130_fd_sc_hd__buf_1 _19768_ (.A(_11433_),
    .X(_11651_));
 sky130_fd_sc_hd__a21oi_1 _19769_ (.A1(_11650_),
    .A2(_11646_),
    .B1(net1020),
    .Y(_11652_));
 sky130_fd_sc_hd__o22a_1 _19770_ (.A1(_11646_),
    .A2(_11647_),
    .B1(_11652_),
    .B2(net266),
    .X(_00349_));
 sky130_fd_sc_hd__inv_2 _19771_ (.A(net259),
    .Y(_11653_));
 sky130_fd_sc_hd__clkbuf_4 _19772_ (.A(_11573_),
    .X(_11654_));
 sky130_fd_sc_hd__mux2_1 _19773_ (.A0(_11415_),
    .A1(_11416_),
    .S(_11654_),
    .X(_11655_));
 sky130_fd_sc_hd__or2_1 _19774_ (.A(net194),
    .B(net190),
    .X(_11656_));
 sky130_fd_sc_hd__buf_2 _19775_ (.A(_11656_),
    .X(_11657_));
 sky130_fd_sc_hd__nor2_1 _19776_ (.A(net181),
    .B(_11657_),
    .Y(_11658_));
 sky130_fd_sc_hd__a22o_1 _19777_ (.A1(net82),
    .A2(_11657_),
    .B1(_11658_),
    .B2(_11575_),
    .X(_11659_));
 sky130_fd_sc_hd__a22o_1 _19778_ (.A1(net181),
    .A2(net82),
    .B1(_11659_),
    .B2(net182),
    .X(_11660_));
 sky130_fd_sc_hd__a21oi_2 _19779_ (.A1(_11655_),
    .A2(_11560_),
    .B1(_11660_),
    .Y(_11661_));
 sky130_fd_sc_hd__nand2_1 _19780_ (.A(_11640_),
    .B(_11641_),
    .Y(_11662_));
 sky130_fd_sc_hd__nand2_1 _19781_ (.A(_11513_),
    .B(_11662_),
    .Y(_11663_));
 sky130_fd_sc_hd__xnor2_2 _19782_ (.A(_11661_),
    .B(_11663_),
    .Y(_11664_));
 sky130_fd_sc_hd__or2_1 _19783_ (.A(net272),
    .B(_11644_),
    .X(_11665_));
 sky130_fd_sc_hd__or2_1 _19784_ (.A(net266),
    .B(_11643_),
    .X(_11666_));
 sky130_fd_sc_hd__and2_1 _19785_ (.A(net266),
    .B(_11643_),
    .X(_11667_));
 sky130_fd_sc_hd__a31o_1 _19786_ (.A1(_11621_),
    .A2(_11665_),
    .A3(_11666_),
    .B1(_11667_),
    .X(_11668_));
 sky130_fd_sc_hd__xor2_1 _19787_ (.A(_11664_),
    .B(_11668_),
    .X(_11669_));
 sky130_fd_sc_hd__o21ai_1 _19788_ (.A1(net1014),
    .A2(_11669_),
    .B1(net174),
    .Y(_11670_));
 sky130_fd_sc_hd__and3_1 _19789_ (.A(net260),
    .B(_11435_),
    .C(_11669_),
    .X(_11671_));
 sky130_fd_sc_hd__a21oi_1 _19790_ (.A1(_11653_),
    .A2(_11670_),
    .B1(_11671_),
    .Y(_00350_));
 sky130_fd_sc_hd__inv_2 _19791_ (.A(net253),
    .Y(_11672_));
 sky130_fd_sc_hd__buf_2 _19792_ (.A(_11672_),
    .X(_11673_));
 sky130_fd_sc_hd__buf_4 _19793_ (.A(_11444_),
    .X(_11674_));
 sky130_fd_sc_hd__nand2_1 _19794_ (.A(_11674_),
    .B(_11448_),
    .Y(_11675_));
 sky130_fd_sc_hd__o21a_1 _19795_ (.A1(_11448_),
    .A2(_11442_),
    .B1(_11675_),
    .X(_11676_));
 sky130_fd_sc_hd__nand2b_1 _19796_ (.A_N(_11662_),
    .B(_11661_),
    .Y(_11677_));
 sky130_fd_sc_hd__nand2_1 _19797_ (.A(_11513_),
    .B(_11677_),
    .Y(_11678_));
 sky130_fd_sc_hd__xor2_1 _19798_ (.A(_11676_),
    .B(_11678_),
    .X(_11679_));
 sky130_fd_sc_hd__inv_2 _19799_ (.A(_11679_),
    .Y(_11680_));
 sky130_fd_sc_hd__o2111a_1 _19800_ (.A1(net259),
    .A2(_11664_),
    .B1(_11665_),
    .C1(_11666_),
    .D1(_11621_),
    .X(_11681_));
 sky130_fd_sc_hd__o21a_1 _19801_ (.A1(net259),
    .A2(_11664_),
    .B1(_11667_),
    .X(_11682_));
 sky130_fd_sc_hd__a211oi_1 _19802_ (.A1(net260),
    .A2(_11664_),
    .B1(_11681_),
    .C1(_11682_),
    .Y(_11683_));
 sky130_fd_sc_hd__nor2_1 _19803_ (.A(_11680_),
    .B(_11683_),
    .Y(_11684_));
 sky130_fd_sc_hd__and2_1 _19804_ (.A(_11680_),
    .B(_11683_),
    .X(_11685_));
 sky130_fd_sc_hd__nor2_1 _19805_ (.A(_11684_),
    .B(_11685_),
    .Y(_11686_));
 sky130_fd_sc_hd__or2_1 _19806_ (.A(_11430_),
    .B(_11686_),
    .X(_11687_));
 sky130_fd_sc_hd__a21oi_1 _19807_ (.A1(net1013),
    .A2(_11686_),
    .B1(_11673_),
    .Y(_11688_));
 sky130_fd_sc_hd__a31o_1 _19808_ (.A1(net175),
    .A2(_11673_),
    .A3(_11687_),
    .B1(_11688_),
    .X(_00351_));
 sky130_fd_sc_hd__clkinv_4 _19809_ (.A(net250),
    .Y(_11689_));
 sky130_fd_sc_hd__a21oi_1 _19810_ (.A1(_11680_),
    .A2(_11683_),
    .B1(_11673_),
    .Y(_11690_));
 sky130_fd_sc_hd__mux2_1 _19811_ (.A0(_11535_),
    .A1(_11536_),
    .S(_11654_),
    .X(_11691_));
 sky130_fd_sc_hd__o21a_1 _19812_ (.A1(_11448_),
    .A2(_11691_),
    .B1(_11675_),
    .X(_11692_));
 sky130_fd_sc_hd__o21a_1 _19813_ (.A1(_11676_),
    .A2(_11677_),
    .B1(_11513_),
    .X(_11693_));
 sky130_fd_sc_hd__xnor2_1 _19814_ (.A(_11692_),
    .B(_11693_),
    .Y(_11694_));
 sky130_fd_sc_hd__o21a_1 _19815_ (.A1(_11684_),
    .A2(_11690_),
    .B1(_11694_),
    .X(_11695_));
 sky130_fd_sc_hd__or3_1 _19816_ (.A(_11684_),
    .B(_11690_),
    .C(_11694_),
    .X(_11696_));
 sky130_fd_sc_hd__and2b_1 _19817_ (.A_N(_11695_),
    .B(_11696_),
    .X(_11697_));
 sky130_fd_sc_hd__or2_1 _19818_ (.A(_11430_),
    .B(_11697_),
    .X(_11698_));
 sky130_fd_sc_hd__a21oi_1 _19819_ (.A1(net1013),
    .A2(_11697_),
    .B1(_11689_),
    .Y(_11699_));
 sky130_fd_sc_hd__a31o_1 _19820_ (.A1(net175),
    .A2(_11689_),
    .A3(_11698_),
    .B1(_11699_),
    .X(_00352_));
 sky130_fd_sc_hd__or3_1 _19821_ (.A(_11676_),
    .B(_11677_),
    .C(_11692_),
    .X(_11700_));
 sky130_fd_sc_hd__o21a_1 _19822_ (.A1(_11448_),
    .A2(_11558_),
    .B1(net82),
    .X(_11701_));
 sky130_fd_sc_hd__a21o_1 _19823_ (.A1(_11560_),
    .A2(_11557_),
    .B1(_11701_),
    .X(_11702_));
 sky130_fd_sc_hd__a21oi_1 _19824_ (.A1(_11514_),
    .A2(_11700_),
    .B1(_11702_),
    .Y(_11703_));
 sky130_fd_sc_hd__and3_1 _19825_ (.A(_11514_),
    .B(_11702_),
    .C(_11700_),
    .X(_11704_));
 sky130_fd_sc_hd__or2_1 _19826_ (.A(_11703_),
    .B(_11704_),
    .X(_11705_));
 sky130_fd_sc_hd__o21ai_1 _19827_ (.A1(net251),
    .A2(_11695_),
    .B1(_11696_),
    .Y(_11706_));
 sky130_fd_sc_hd__xnor2_1 _19828_ (.A(_11705_),
    .B(_11706_),
    .Y(_11707_));
 sky130_fd_sc_hd__o21a_1 _19829_ (.A1(_11430_),
    .A2(_11707_),
    .B1(net175),
    .X(_11708_));
 sky130_fd_sc_hd__nand2_1 _19830_ (.A(_11435_),
    .B(_11707_),
    .Y(_11709_));
 sky130_fd_sc_hd__mux2_1 _19831_ (.A0(_11708_),
    .A1(_11709_),
    .S(net248),
    .X(_11710_));
 sky130_fd_sc_hd__clkbuf_1 _19832_ (.A(_11710_),
    .X(_00353_));
 sky130_fd_sc_hd__nand2_1 _19833_ (.A(net244),
    .B(_11705_),
    .Y(_11711_));
 sky130_fd_sc_hd__nor2_1 _19834_ (.A(net244),
    .B(_11705_),
    .Y(_11712_));
 sky130_fd_sc_hd__a21o_1 _19835_ (.A1(_11706_),
    .A2(_11711_),
    .B1(_11712_),
    .X(_11713_));
 sky130_fd_sc_hd__nand2_1 _19836_ (.A(_11654_),
    .B(_11560_),
    .Y(_11714_));
 sky130_fd_sc_hd__nand2_1 _19837_ (.A(_11632_),
    .B(_11560_),
    .Y(_11715_));
 sky130_fd_sc_hd__o22a_1 _19838_ (.A1(_11632_),
    .A2(net83),
    .B1(_11575_),
    .B2(_11715_),
    .X(_11716_));
 sky130_fd_sc_hd__o221a_2 _19839_ (.A1(_11415_),
    .A2(_11714_),
    .B1(_11716_),
    .B2(_11654_),
    .C1(_11675_),
    .X(_11717_));
 sky130_fd_sc_hd__inv_2 _19840_ (.A(_11717_),
    .Y(_11718_));
 sky130_fd_sc_hd__or2_1 _19841_ (.A(_11702_),
    .B(_11700_),
    .X(_11719_));
 sky130_fd_sc_hd__and2_1 _19842_ (.A(_11514_),
    .B(_11719_),
    .X(_11720_));
 sky130_fd_sc_hd__xnor2_2 _19843_ (.A(_11718_),
    .B(_11720_),
    .Y(_11721_));
 sky130_fd_sc_hd__xor2_1 _19844_ (.A(_11713_),
    .B(_11721_),
    .X(_11722_));
 sky130_fd_sc_hd__o21a_1 _19845_ (.A1(_11430_),
    .A2(_11722_),
    .B1(net175),
    .X(_11723_));
 sky130_fd_sc_hd__nand2_1 _19846_ (.A(_11435_),
    .B(_11722_),
    .Y(_11724_));
 sky130_fd_sc_hd__mux2_1 _19847_ (.A0(_11723_),
    .A1(_11724_),
    .S(net241),
    .X(_11725_));
 sky130_fd_sc_hd__clkbuf_1 _19848_ (.A(_11725_),
    .X(_00354_));
 sky130_fd_sc_hd__inv_2 _19849_ (.A(net234),
    .Y(_11726_));
 sky130_fd_sc_hd__buf_4 _19850_ (.A(_11726_),
    .X(_11727_));
 sky130_fd_sc_hd__or2_1 _19851_ (.A(_11717_),
    .B(_11719_),
    .X(_11728_));
 sky130_fd_sc_hd__and2_1 _19852_ (.A(_11514_),
    .B(_11728_),
    .X(_11729_));
 sky130_fd_sc_hd__clkbuf_4 _19853_ (.A(_11451_),
    .X(_11730_));
 sky130_fd_sc_hd__mux2_1 _19854_ (.A0(net82),
    .A1(_11440_),
    .S(_11730_),
    .X(_11731_));
 sky130_fd_sc_hd__buf_2 _19855_ (.A(_11731_),
    .X(_11732_));
 sky130_fd_sc_hd__xor2_2 _19856_ (.A(_11729_),
    .B(_11732_),
    .X(_11733_));
 sky130_fd_sc_hd__o21ba_1 _19857_ (.A1(_11713_),
    .A2(_11721_),
    .B1_N(net241),
    .X(_11734_));
 sky130_fd_sc_hd__a21oi_1 _19858_ (.A1(_11713_),
    .A2(_11721_),
    .B1(_11734_),
    .Y(_11735_));
 sky130_fd_sc_hd__xnor2_1 _19859_ (.A(_11733_),
    .B(_11735_),
    .Y(_11736_));
 sky130_fd_sc_hd__or2_1 _19860_ (.A(_11430_),
    .B(_11736_),
    .X(_11737_));
 sky130_fd_sc_hd__a21oi_1 _19861_ (.A1(net1013),
    .A2(_11736_),
    .B1(_11727_),
    .Y(_11738_));
 sky130_fd_sc_hd__a31o_1 _19862_ (.A1(net175),
    .A2(_11727_),
    .A3(_11737_),
    .B1(_11738_),
    .X(_00355_));
 sky130_fd_sc_hd__clkinv_4 _19863_ (.A(net229),
    .Y(_11739_));
 sky130_fd_sc_hd__mux2_1 _19864_ (.A0(net82),
    .A1(_11535_),
    .S(_11730_),
    .X(_11740_));
 sky130_fd_sc_hd__o21ai_1 _19865_ (.A1(_11728_),
    .A2(_11732_),
    .B1(_11514_),
    .Y(_11741_));
 sky130_fd_sc_hd__xnor2_2 _19866_ (.A(_11740_),
    .B(_11741_),
    .Y(_11742_));
 sky130_fd_sc_hd__xnor2_1 _19867_ (.A(_11727_),
    .B(_11733_),
    .Y(_11743_));
 sky130_fd_sc_hd__xor2_1 _19868_ (.A(net241),
    .B(_11721_),
    .X(_11744_));
 sky130_fd_sc_hd__mux2_1 _19869_ (.A0(net237),
    .A1(_11514_),
    .S(_11717_),
    .X(_11745_));
 sky130_fd_sc_hd__o21ai_1 _19870_ (.A1(net243),
    .A2(_11729_),
    .B1(_11745_),
    .Y(_11746_));
 sky130_fd_sc_hd__a21o_1 _19871_ (.A1(_11719_),
    .A2(_11732_),
    .B1(net237),
    .X(_11747_));
 sky130_fd_sc_hd__o31ai_1 _19872_ (.A1(_11519_),
    .A2(_11719_),
    .A3(_11732_),
    .B1(_11747_),
    .Y(_11748_));
 sky130_fd_sc_hd__o31a_1 _19873_ (.A1(_11519_),
    .A2(_11718_),
    .A3(_11732_),
    .B1(net237),
    .X(_11749_));
 sky130_fd_sc_hd__nor2_1 _19874_ (.A(_11717_),
    .B(_11732_),
    .Y(_11750_));
 sky130_fd_sc_hd__a2bb2o_1 _19875_ (.A1_N(net243),
    .A2_N(_11749_),
    .B1(_11750_),
    .B2(_11720_),
    .X(_11751_));
 sky130_fd_sc_hd__a221o_1 _19876_ (.A1(_11732_),
    .A2(_11746_),
    .B1(_11748_),
    .B2(_11717_),
    .C1(_11751_),
    .X(_11752_));
 sky130_fd_sc_hd__o31a_1 _19877_ (.A1(_11713_),
    .A2(_11743_),
    .A3(_11744_),
    .B1(_11752_),
    .X(_11753_));
 sky130_fd_sc_hd__xor2_1 _19878_ (.A(_11742_),
    .B(_11753_),
    .X(_11754_));
 sky130_fd_sc_hd__o21ai_1 _19879_ (.A1(_11526_),
    .A2(_11754_),
    .B1(net175),
    .Y(_11755_));
 sky130_fd_sc_hd__and3_1 _19880_ (.A(net232),
    .B(_11435_),
    .C(_11754_),
    .X(_11756_));
 sky130_fd_sc_hd__a21oi_1 _19881_ (.A1(_11739_),
    .A2(_11755_),
    .B1(_11756_),
    .Y(_00356_));
 sky130_fd_sc_hd__inv_2 _19882_ (.A(net225),
    .Y(_11757_));
 sky130_fd_sc_hd__buf_4 _19883_ (.A(_11757_),
    .X(_11758_));
 sky130_fd_sc_hd__clkbuf_4 _19884_ (.A(_11758_),
    .X(_11759_));
 sky130_fd_sc_hd__nand2_1 _19885_ (.A(_11730_),
    .B(_11629_),
    .Y(_11760_));
 sky130_fd_sc_hd__a2bb2o_2 _19886_ (.A1_N(_11714_),
    .A2_N(_11634_),
    .B1(_11760_),
    .B2(net83),
    .X(_11761_));
 sky130_fd_sc_hd__or3_1 _19887_ (.A(_11728_),
    .B(_11732_),
    .C(_11740_),
    .X(_11762_));
 sky130_fd_sc_hd__nand2_1 _19888_ (.A(_11515_),
    .B(_11762_),
    .Y(_11763_));
 sky130_fd_sc_hd__xor2_2 _19889_ (.A(_11761_),
    .B(_11763_),
    .X(_11764_));
 sky130_fd_sc_hd__o21a_1 _19890_ (.A1(_11742_),
    .A2(_11753_),
    .B1(_11739_),
    .X(_11765_));
 sky130_fd_sc_hd__a21o_1 _19891_ (.A1(_11742_),
    .A2(_11753_),
    .B1(_11765_),
    .X(_11766_));
 sky130_fd_sc_hd__xnor2_1 _19892_ (.A(_11764_),
    .B(_11766_),
    .Y(_11767_));
 sky130_fd_sc_hd__o21ai_1 _19893_ (.A1(_11526_),
    .A2(_11767_),
    .B1(net175),
    .Y(_11768_));
 sky130_fd_sc_hd__and3_1 _19894_ (.A(net227),
    .B(_11435_),
    .C(_11767_),
    .X(_11769_));
 sky130_fd_sc_hd__a21oi_1 _19895_ (.A1(_11759_),
    .A2(_11768_),
    .B1(_11769_),
    .Y(_00357_));
 sky130_fd_sc_hd__nor2_1 _19896_ (.A(net228),
    .B(_11764_),
    .Y(_11770_));
 sky130_fd_sc_hd__a211o_1 _19897_ (.A1(_11742_),
    .A2(_11753_),
    .B1(_11765_),
    .C1(_11770_),
    .X(_11771_));
 sky130_fd_sc_hd__nand2_1 _19898_ (.A(net228),
    .B(_11764_),
    .Y(_11772_));
 sky130_fd_sc_hd__o21ai_1 _19899_ (.A1(_11761_),
    .A2(_11762_),
    .B1(_11515_),
    .Y(_11773_));
 sky130_fd_sc_hd__or2_1 _19900_ (.A(net194),
    .B(net184),
    .X(_11774_));
 sky130_fd_sc_hd__or2_2 _19901_ (.A(net190),
    .B(_11774_),
    .X(_11775_));
 sky130_fd_sc_hd__or2_1 _19902_ (.A(net181),
    .B(_11775_),
    .X(_11776_));
 sky130_fd_sc_hd__mux2_1 _19903_ (.A0(_11575_),
    .A1(net82),
    .S(_11776_),
    .X(_11777_));
 sky130_fd_sc_hd__xnor2_1 _19904_ (.A(_11773_),
    .B(_11777_),
    .Y(_11778_));
 sky130_fd_sc_hd__a21oi_1 _19905_ (.A1(_11771_),
    .A2(_11772_),
    .B1(_11778_),
    .Y(_11779_));
 sky130_fd_sc_hd__and3_1 _19906_ (.A(_11778_),
    .B(_11771_),
    .C(_11772_),
    .X(_11780_));
 sky130_fd_sc_hd__nor2_1 _19907_ (.A(_11779_),
    .B(_11780_),
    .Y(_11781_));
 sky130_fd_sc_hd__o21ai_1 _19908_ (.A1(_11431_),
    .A2(_11781_),
    .B1(net175),
    .Y(_11782_));
 sky130_fd_sc_hd__nand2_1 _19909_ (.A(net176),
    .B(_11648_),
    .Y(_11783_));
 sky130_fd_sc_hd__clkbuf_4 _19910_ (.A(_11783_),
    .X(_11784_));
 sky130_fd_sc_hd__clkbuf_4 _19911_ (.A(_11784_),
    .X(_11785_));
 sky130_fd_sc_hd__nor2_1 _19912_ (.A(net224),
    .B(_11785_),
    .Y(_11786_));
 sky130_fd_sc_hd__a22o_1 _19913_ (.A1(net224),
    .A2(_11782_),
    .B1(_11786_),
    .B2(_11781_),
    .X(_00358_));
 sky130_fd_sc_hd__inv_2 _19914_ (.A(net214),
    .Y(_11787_));
 sky130_fd_sc_hd__buf_6 _19915_ (.A(_11787_),
    .X(_11788_));
 sky130_fd_sc_hd__buf_4 _19916_ (.A(_11788_),
    .X(_11789_));
 sky130_fd_sc_hd__o31a_1 _19917_ (.A1(_11761_),
    .A2(_11762_),
    .A3(_11777_),
    .B1(_11515_),
    .X(_11790_));
 sky130_fd_sc_hd__xnor2_1 _19918_ (.A(net82),
    .B(_11790_),
    .Y(_11791_));
 sky130_fd_sc_hd__o21ba_1 _19919_ (.A1(net224),
    .A2(_11779_),
    .B1_N(_11780_),
    .X(_11792_));
 sky130_fd_sc_hd__xnor2_1 _19920_ (.A(_11791_),
    .B(_11792_),
    .Y(_11793_));
 sky130_fd_sc_hd__a21oi_1 _19921_ (.A1(_11650_),
    .A2(_11793_),
    .B1(net1020),
    .Y(_11794_));
 sky130_fd_sc_hd__or3_1 _19922_ (.A(net220),
    .B(_11784_),
    .C(_11793_),
    .X(_11795_));
 sky130_fd_sc_hd__o21ai_1 _19923_ (.A1(_11789_),
    .A2(_11794_),
    .B1(_11795_),
    .Y(_00359_));
 sky130_fd_sc_hd__or3_1 _19924_ (.A(_11632_),
    .B(net202),
    .C(net184),
    .X(_11796_));
 sky130_fd_sc_hd__nor2_1 _19925_ (.A(net194),
    .B(_11576_),
    .Y(_11797_));
 sky130_fd_sc_hd__o21ai_1 _19926_ (.A1(net190),
    .A2(_11797_),
    .B1(net201),
    .Y(_11798_));
 sky130_fd_sc_hd__a21oi_2 _19927_ (.A1(_11796_),
    .A2(_11798_),
    .B1(net181),
    .Y(_11799_));
 sky130_fd_sc_hd__o21ai_1 _19928_ (.A1(_11431_),
    .A2(_11799_),
    .B1(net177),
    .Y(_11800_));
 sky130_fd_sc_hd__nor2_1 _19929_ (.A(\top0.cordic0.slte0.opA[0] ),
    .B(_11785_),
    .Y(_11801_));
 sky130_fd_sc_hd__a22o_1 _19930_ (.A1(net901),
    .A2(_11800_),
    .B1(_11801_),
    .B2(_11799_),
    .X(_00360_));
 sky130_fd_sc_hd__and2_1 _19931_ (.A(\top0.cordic0.slte0.opA[0] ),
    .B(_11799_),
    .X(_11802_));
 sky130_fd_sc_hd__nor2_1 _19932_ (.A(_11576_),
    .B(_11427_),
    .Y(_11803_));
 sky130_fd_sc_hd__or3_1 _19933_ (.A(net201),
    .B(net184),
    .C(net190),
    .X(_11804_));
 sky130_fd_sc_hd__nor2_1 _19934_ (.A(_11632_),
    .B(_11804_),
    .Y(_11805_));
 sky130_fd_sc_hd__o22a_1 _19935_ (.A1(_11510_),
    .A2(_11803_),
    .B1(_11805_),
    .B2(_11797_),
    .X(_11806_));
 sky130_fd_sc_hd__nor2_2 _19936_ (.A(_11410_),
    .B(net1016),
    .Y(_11807_));
 sky130_fd_sc_hd__nor2_2 _19937_ (.A(net201),
    .B(_11510_),
    .Y(_11808_));
 sky130_fd_sc_hd__o21a_1 _19938_ (.A1(_11807_),
    .A2(_11808_),
    .B1(net195),
    .X(_11809_));
 sky130_fd_sc_hd__nor2_1 _19939_ (.A(net195),
    .B(_11410_),
    .Y(_11810_));
 sky130_fd_sc_hd__or2_1 _19940_ (.A(net183),
    .B(_11509_),
    .X(_11811_));
 sky130_fd_sc_hd__and2_1 _19941_ (.A(_11484_),
    .B(_11504_),
    .X(_11812_));
 sky130_fd_sc_hd__nand2_1 _19942_ (.A(net202),
    .B(net183),
    .Y(_11813_));
 sky130_fd_sc_hd__o221a_1 _19943_ (.A1(net183),
    .A2(_11810_),
    .B1(_11811_),
    .B2(_11812_),
    .C1(_11813_),
    .X(_11814_));
 sky130_fd_sc_hd__o21a_1 _19944_ (.A1(_11809_),
    .A2(_11814_),
    .B1(net189),
    .X(_11815_));
 sky130_fd_sc_hd__o21a_1 _19945_ (.A1(_11806_),
    .A2(_11815_),
    .B1(_11426_),
    .X(_11816_));
 sky130_fd_sc_hd__xor2_1 _19946_ (.A(_11802_),
    .B(_11816_),
    .X(_11817_));
 sky130_fd_sc_hd__o21ai_1 _19947_ (.A1(_11431_),
    .A2(_11817_),
    .B1(net177),
    .Y(_11818_));
 sky130_fd_sc_hd__nor2_1 _19948_ (.A(\top0.cordic0.slte0.opA[1] ),
    .B(_11785_),
    .Y(_11819_));
 sky130_fd_sc_hd__a22o_1 _19949_ (.A1(\top0.cordic0.slte0.opA[1] ),
    .A2(_11818_),
    .B1(_11819_),
    .B2(_11817_),
    .X(_00361_));
 sky130_fd_sc_hd__o211a_1 _19950_ (.A1(_11807_),
    .A2(_11808_),
    .B1(net195),
    .C1(net189),
    .X(_11820_));
 sky130_fd_sc_hd__a221o_1 _19951_ (.A1(\top0.cordic0.slte0.opA[1] ),
    .A2(_11802_),
    .B1(_11814_),
    .B2(net189),
    .C1(_11806_),
    .X(_11821_));
 sky130_fd_sc_hd__o221ai_4 _19952_ (.A1(\top0.cordic0.slte0.opA[1] ),
    .A2(_11802_),
    .B1(_11820_),
    .B2(_11821_),
    .C1(_11426_),
    .Y(_11822_));
 sky130_fd_sc_hd__nand2_1 _19953_ (.A(net195),
    .B(net183),
    .Y(_11823_));
 sky130_fd_sc_hd__nor2_1 _19954_ (.A(_11410_),
    .B(net185),
    .Y(_11824_));
 sky130_fd_sc_hd__and4b_1 _19955_ (.A_N(_11824_),
    .B(net189),
    .C(net195),
    .D(net1016),
    .X(_11825_));
 sky130_fd_sc_hd__a31o_1 _19956_ (.A1(net189),
    .A2(_11823_),
    .A3(_11807_),
    .B1(_11825_),
    .X(_11826_));
 sky130_fd_sc_hd__a21oi_1 _19957_ (.A1(net185),
    .A2(_11510_),
    .B1(_11657_),
    .Y(_11827_));
 sky130_fd_sc_hd__a31o_1 _19958_ (.A1(_11654_),
    .A2(_11510_),
    .A3(_11633_),
    .B1(_11827_),
    .X(_11828_));
 sky130_fd_sc_hd__a2111o_1 _19959_ (.A1(net183),
    .A2(_11808_),
    .B1(_11826_),
    .C1(_11828_),
    .D1(net181),
    .X(_11829_));
 sky130_fd_sc_hd__xor2_1 _19960_ (.A(_11822_),
    .B(_11829_),
    .X(_11830_));
 sky130_fd_sc_hd__o21ai_1 _19961_ (.A1(_11431_),
    .A2(_11830_),
    .B1(net177),
    .Y(_11831_));
 sky130_fd_sc_hd__nor2_1 _19962_ (.A(\top0.cordic0.slte0.opA[2] ),
    .B(_11785_),
    .Y(_11832_));
 sky130_fd_sc_hd__a22o_1 _19963_ (.A1(net992),
    .A2(_11831_),
    .B1(_11832_),
    .B2(_11830_),
    .X(_00362_));
 sky130_fd_sc_hd__or2_1 _19964_ (.A(_11612_),
    .B(_11574_),
    .X(_11833_));
 sky130_fd_sc_hd__a31o_1 _19965_ (.A1(net195),
    .A2(net185),
    .A3(net189),
    .B1(net201),
    .X(_11834_));
 sky130_fd_sc_hd__a21o_1 _19966_ (.A1(_11517_),
    .A2(_11834_),
    .B1(net181),
    .X(_11835_));
 sky130_fd_sc_hd__a311o_2 _19967_ (.A1(_11410_),
    .A2(_11511_),
    .A3(_11833_),
    .B1(_11835_),
    .C1(_11827_),
    .X(_11836_));
 sky130_fd_sc_hd__nor2_1 _19968_ (.A(_11822_),
    .B(_11829_),
    .Y(_11837_));
 sky130_fd_sc_hd__a21boi_1 _19969_ (.A1(_11822_),
    .A2(_11829_),
    .B1_N(\top0.cordic0.slte0.opA[2] ),
    .Y(_11838_));
 sky130_fd_sc_hd__nor2_1 _19970_ (.A(_11837_),
    .B(_11838_),
    .Y(_11839_));
 sky130_fd_sc_hd__xor2_1 _19971_ (.A(_11836_),
    .B(_11839_),
    .X(_11840_));
 sky130_fd_sc_hd__o21ai_1 _19972_ (.A1(_11431_),
    .A2(_11840_),
    .B1(net177),
    .Y(_11841_));
 sky130_fd_sc_hd__nor2_1 _19973_ (.A(\top0.cordic0.slte0.opA[3] ),
    .B(_11785_),
    .Y(_11842_));
 sky130_fd_sc_hd__a22o_1 _19974_ (.A1(\top0.cordic0.slte0.opA[3] ),
    .A2(_11841_),
    .B1(_11842_),
    .B2(_11840_),
    .X(_00363_));
 sky130_fd_sc_hd__a2111o_1 _19975_ (.A1(_11484_),
    .A2(_11504_),
    .B1(_11509_),
    .C1(net189),
    .D1(_11410_),
    .X(_11843_));
 sky130_fd_sc_hd__o21ai_1 _19976_ (.A1(_11573_),
    .A2(_11510_),
    .B1(_11843_),
    .Y(_11844_));
 sky130_fd_sc_hd__nor2_1 _19977_ (.A(_11632_),
    .B(net183),
    .Y(_11845_));
 sky130_fd_sc_hd__a21o_1 _19978_ (.A1(_11509_),
    .A2(_11845_),
    .B1(_11413_),
    .X(_11846_));
 sky130_fd_sc_hd__or4b_1 _19979_ (.A(net183),
    .B(_11573_),
    .C(_11509_),
    .D_N(_11810_),
    .X(_11847_));
 sky130_fd_sc_hd__a21oi_1 _19980_ (.A1(_11484_),
    .A2(_11504_),
    .B1(_11847_),
    .Y(_11848_));
 sky130_fd_sc_hd__a211o_1 _19981_ (.A1(_11812_),
    .A2(_11845_),
    .B1(_11846_),
    .C1(_11848_),
    .X(_11849_));
 sky130_fd_sc_hd__a2111oi_1 _19982_ (.A1(net184),
    .A2(_11844_),
    .B1(_11849_),
    .C1(net181),
    .D1(_11808_),
    .Y(_11850_));
 sky130_fd_sc_hd__inv_2 _19983_ (.A(\top0.cordic0.slte0.opA[3] ),
    .Y(_11851_));
 sky130_fd_sc_hd__nand2_1 _19984_ (.A(_11851_),
    .B(_11836_),
    .Y(_11852_));
 sky130_fd_sc_hd__nor2_1 _19985_ (.A(_11851_),
    .B(_11836_),
    .Y(_11853_));
 sky130_fd_sc_hd__or3_1 _19986_ (.A(_11837_),
    .B(_11838_),
    .C(_11853_),
    .X(_11854_));
 sky130_fd_sc_hd__nand2_1 _19987_ (.A(_11852_),
    .B(_11854_),
    .Y(_11855_));
 sky130_fd_sc_hd__xnor2_1 _19988_ (.A(net10),
    .B(_11855_),
    .Y(_11856_));
 sky130_fd_sc_hd__buf_4 _19989_ (.A(_11783_),
    .X(_11857_));
 sky130_fd_sc_hd__nor2_1 _19990_ (.A(\top0.cordic0.slte0.opA[4] ),
    .B(_11857_),
    .Y(_11858_));
 sky130_fd_sc_hd__o21ai_1 _19991_ (.A1(_11431_),
    .A2(_11856_),
    .B1(net177),
    .Y(_11859_));
 sky130_fd_sc_hd__a22o_1 _19992_ (.A1(_11856_),
    .A2(_11858_),
    .B1(_11859_),
    .B2(net981),
    .X(_00364_));
 sky130_fd_sc_hd__inv_2 _19993_ (.A(_11807_),
    .Y(_11860_));
 sky130_fd_sc_hd__nand2_1 _19994_ (.A(net189),
    .B(_11511_),
    .Y(_11861_));
 sky130_fd_sc_hd__or3_1 _19995_ (.A(net202),
    .B(net190),
    .C(_11510_),
    .X(_11862_));
 sky130_fd_sc_hd__o311a_1 _19996_ (.A1(net202),
    .A2(_11573_),
    .A3(_11510_),
    .B1(_11612_),
    .C1(_11632_),
    .X(_11863_));
 sky130_fd_sc_hd__a31o_1 _19997_ (.A1(_11774_),
    .A2(_11861_),
    .A3(_11862_),
    .B1(_11863_),
    .X(_11864_));
 sky130_fd_sc_hd__a21oi_2 _19998_ (.A1(_11860_),
    .A2(_11864_),
    .B1(\top0.cordic0.gm0.iter[4] ),
    .Y(_11865_));
 sky130_fd_sc_hd__and2_1 _19999_ (.A(\top0.cordic0.slte0.opA[4] ),
    .B(net10),
    .X(_11866_));
 sky130_fd_sc_hd__a21o_1 _20000_ (.A1(_11852_),
    .A2(_11854_),
    .B1(_11866_),
    .X(_11867_));
 sky130_fd_sc_hd__or2_1 _20001_ (.A(\top0.cordic0.slte0.opA[4] ),
    .B(net1012),
    .X(_11868_));
 sky130_fd_sc_hd__nand2_1 _20002_ (.A(_11867_),
    .B(_11868_),
    .Y(_11869_));
 sky130_fd_sc_hd__xnor2_1 _20003_ (.A(_11865_),
    .B(_11869_),
    .Y(_11870_));
 sky130_fd_sc_hd__o21ai_1 _20004_ (.A1(_11431_),
    .A2(_11870_),
    .B1(net177),
    .Y(_11871_));
 sky130_fd_sc_hd__nor2_1 _20005_ (.A(\top0.cordic0.slte0.opA[5] ),
    .B(_11785_),
    .Y(_11872_));
 sky130_fd_sc_hd__a22o_1 _20006_ (.A1(\top0.cordic0.slte0.opA[5] ),
    .A2(_11871_),
    .B1(_11872_),
    .B2(_11870_),
    .X(_00365_));
 sky130_fd_sc_hd__nor2_1 _20007_ (.A(net189),
    .B(_11824_),
    .Y(_11873_));
 sky130_fd_sc_hd__o221a_1 _20008_ (.A1(net201),
    .A2(_11411_),
    .B1(_11873_),
    .B2(net194),
    .C1(_11823_),
    .X(_11874_));
 sky130_fd_sc_hd__nand2_1 _20009_ (.A(_11512_),
    .B(_11874_),
    .Y(_11875_));
 sky130_fd_sc_hd__nor2_1 _20010_ (.A(_11612_),
    .B(net190),
    .Y(_11876_));
 sky130_fd_sc_hd__a21oi_1 _20011_ (.A1(_11410_),
    .A2(\top0.cordic0.gm0.iter[2] ),
    .B1(net183),
    .Y(_11877_));
 sky130_fd_sc_hd__a221o_1 _20012_ (.A1(_11876_),
    .A2(_11810_),
    .B1(_11877_),
    .B2(net195),
    .C1(_11512_),
    .X(_11878_));
 sky130_fd_sc_hd__and3_1 _20013_ (.A(_11426_),
    .B(_11875_),
    .C(_11878_),
    .X(_11879_));
 sky130_fd_sc_hd__inv_2 _20014_ (.A(_11879_),
    .Y(_11880_));
 sky130_fd_sc_hd__and3_1 _20015_ (.A(_11852_),
    .B(_11865_),
    .C(_11868_),
    .X(_11881_));
 sky130_fd_sc_hd__and3_1 _20016_ (.A(\top0.cordic0.slte0.opA[5] ),
    .B(_11852_),
    .C(_11868_),
    .X(_11882_));
 sky130_fd_sc_hd__o32a_1 _20017_ (.A1(_11837_),
    .A2(_11838_),
    .A3(_11853_),
    .B1(_11881_),
    .B2(_11882_),
    .X(_11883_));
 sky130_fd_sc_hd__o21a_1 _20018_ (.A1(\top0.cordic0.slte0.opA[5] ),
    .A2(_11866_),
    .B1(_11865_),
    .X(_11884_));
 sky130_fd_sc_hd__a21o_1 _20019_ (.A1(\top0.cordic0.slte0.opA[5] ),
    .A2(_11866_),
    .B1(_11884_),
    .X(_11885_));
 sky130_fd_sc_hd__nor2_1 _20020_ (.A(_11883_),
    .B(_11885_),
    .Y(_11886_));
 sky130_fd_sc_hd__xnor2_1 _20021_ (.A(_11880_),
    .B(_11886_),
    .Y(_11887_));
 sky130_fd_sc_hd__a21o_1 _20022_ (.A1(_11650_),
    .A2(_11887_),
    .B1(net1020),
    .X(_11888_));
 sky130_fd_sc_hd__or3_1 _20023_ (.A(\top0.cordic0.slte0.opA[6] ),
    .B(_11784_),
    .C(_11887_),
    .X(_11889_));
 sky130_fd_sc_hd__a21bo_1 _20024_ (.A1(\top0.cordic0.slte0.opA[6] ),
    .A2(_11888_),
    .B1_N(_11889_),
    .X(_00366_));
 sky130_fd_sc_hd__o21a_1 _20025_ (.A1(net201),
    .A2(net185),
    .B1(net195),
    .X(_11890_));
 sky130_fd_sc_hd__a211o_1 _20026_ (.A1(net201),
    .A2(net185),
    .B1(_11574_),
    .C1(_11890_),
    .X(_11891_));
 sky130_fd_sc_hd__nor2_1 _20027_ (.A(net201),
    .B(_11612_),
    .Y(_11892_));
 sky130_fd_sc_hd__nor2_1 _20028_ (.A(_11892_),
    .B(_11824_),
    .Y(_11893_));
 sky130_fd_sc_hd__o211ai_1 _20029_ (.A1(_11657_),
    .A2(_11893_),
    .B1(_11796_),
    .C1(_11518_),
    .Y(_11894_));
 sky130_fd_sc_hd__o211a_1 _20030_ (.A1(_11518_),
    .A2(_11891_),
    .B1(_11894_),
    .C1(_11426_),
    .X(_11895_));
 sky130_fd_sc_hd__o31ai_1 _20031_ (.A1(_11879_),
    .A2(_11883_),
    .A3(_11885_),
    .B1(\top0.cordic0.slte0.opA[6] ),
    .Y(_11896_));
 sky130_fd_sc_hd__o21ai_1 _20032_ (.A1(_11880_),
    .A2(_11886_),
    .B1(_11896_),
    .Y(_11897_));
 sky130_fd_sc_hd__xor2_1 _20033_ (.A(_11895_),
    .B(_11897_),
    .X(_11898_));
 sky130_fd_sc_hd__o21ai_1 _20034_ (.A1(_11431_),
    .A2(_11898_),
    .B1(net178),
    .Y(_11899_));
 sky130_fd_sc_hd__nor2_1 _20035_ (.A(\top0.cordic0.slte0.opA[7] ),
    .B(_11785_),
    .Y(_11900_));
 sky130_fd_sc_hd__a22o_1 _20036_ (.A1(\top0.cordic0.slte0.opA[7] ),
    .A2(_11899_),
    .B1(_11900_),
    .B2(_11898_),
    .X(_00367_));
 sky130_fd_sc_hd__nor2_1 _20037_ (.A(_11632_),
    .B(\top0.cordic0.gm0.iter[2] ),
    .Y(_11901_));
 sky130_fd_sc_hd__nand2_1 _20038_ (.A(_11612_),
    .B(_11518_),
    .Y(_11902_));
 sky130_fd_sc_hd__or2_1 _20039_ (.A(_11518_),
    .B(_11877_),
    .X(_11903_));
 sky130_fd_sc_hd__nor2_1 _20040_ (.A(net202),
    .B(_11902_),
    .Y(_11904_));
 sky130_fd_sc_hd__o21ai_1 _20041_ (.A1(_11807_),
    .A2(_11904_),
    .B1(_11901_),
    .Y(_11905_));
 sky130_fd_sc_hd__o311a_1 _20042_ (.A1(_11410_),
    .A2(_11901_),
    .A3(_11902_),
    .B1(_11903_),
    .C1(_11905_),
    .X(_11906_));
 sky130_fd_sc_hd__nor2_1 _20043_ (.A(net181),
    .B(_11906_),
    .Y(_11907_));
 sky130_fd_sc_hd__nor2_1 _20044_ (.A(\top0.cordic0.slte0.opA[7] ),
    .B(_11895_),
    .Y(_11908_));
 sky130_fd_sc_hd__or2_1 _20045_ (.A(_11880_),
    .B(_11908_),
    .X(_11909_));
 sky130_fd_sc_hd__nand2_1 _20046_ (.A(\top0.cordic0.slte0.opA[7] ),
    .B(_11895_),
    .Y(_11910_));
 sky130_fd_sc_hd__o221a_1 _20047_ (.A1(_11896_),
    .A2(_11908_),
    .B1(_11909_),
    .B2(_11886_),
    .C1(_11910_),
    .X(_11911_));
 sky130_fd_sc_hd__xor2_1 _20048_ (.A(_11907_),
    .B(_11911_),
    .X(_11912_));
 sky130_fd_sc_hd__a21o_1 _20049_ (.A1(_11650_),
    .A2(_11912_),
    .B1(net1020),
    .X(_11913_));
 sky130_fd_sc_hd__or3_1 _20050_ (.A(\top0.cordic0.slte0.opA[8] ),
    .B(_11784_),
    .C(_11912_),
    .X(_11914_));
 sky130_fd_sc_hd__a21bo_1 _20051_ (.A1(net932),
    .A2(_11913_),
    .B1_N(_11914_),
    .X(_00368_));
 sky130_fd_sc_hd__a22o_1 _20052_ (.A1(net183),
    .A2(_11513_),
    .B1(_11657_),
    .B2(_11904_),
    .X(_11915_));
 sky130_fd_sc_hd__mux2_1 _20053_ (.A0(_11902_),
    .A1(_11518_),
    .S(_11657_),
    .X(_11916_));
 sky130_fd_sc_hd__nor2_1 _20054_ (.A(_11410_),
    .B(_11916_),
    .Y(_11917_));
 sky130_fd_sc_hd__o21a_1 _20055_ (.A1(_11915_),
    .A2(_11917_),
    .B1(_11426_),
    .X(_11918_));
 sky130_fd_sc_hd__o21ba_1 _20056_ (.A1(\top0.cordic0.slte0.opA[8] ),
    .A2(_11907_),
    .B1_N(_11911_),
    .X(_11919_));
 sky130_fd_sc_hd__a21oi_1 _20057_ (.A1(\top0.cordic0.slte0.opA[8] ),
    .A2(_11907_),
    .B1(_11919_),
    .Y(_11920_));
 sky130_fd_sc_hd__xnor2_1 _20058_ (.A(_11918_),
    .B(_11920_),
    .Y(_11921_));
 sky130_fd_sc_hd__o21a_1 _20059_ (.A1(_11526_),
    .A2(_11921_),
    .B1(net178),
    .X(_11922_));
 sky130_fd_sc_hd__nor2_1 _20060_ (.A(_11494_),
    .B(_11922_),
    .Y(_11923_));
 sky130_fd_sc_hd__a31o_1 _20061_ (.A1(_11494_),
    .A2(net1013),
    .A3(_11921_),
    .B1(_11923_),
    .X(_00369_));
 sky130_fd_sc_hd__and2_1 _20062_ (.A(\top0.cordic0.slte0.opA[9] ),
    .B(_11918_),
    .X(_11924_));
 sky130_fd_sc_hd__o21ba_1 _20063_ (.A1(\top0.cordic0.slte0.opA[9] ),
    .A2(_11918_),
    .B1_N(_11920_),
    .X(_11925_));
 sky130_fd_sc_hd__o21ai_1 _20064_ (.A1(net190),
    .A2(_11902_),
    .B1(_11861_),
    .Y(_11926_));
 sky130_fd_sc_hd__and3_1 _20065_ (.A(_11612_),
    .B(net190),
    .C(_11518_),
    .X(_11927_));
 sky130_fd_sc_hd__a21o_1 _20066_ (.A1(_11654_),
    .A2(_11513_),
    .B1(_11927_),
    .X(_11928_));
 sky130_fd_sc_hd__a22oi_1 _20067_ (.A1(net195),
    .A2(_11926_),
    .B1(_11928_),
    .B2(_11810_),
    .Y(_11929_));
 sky130_fd_sc_hd__a21oi_1 _20068_ (.A1(_11903_),
    .A2(_11929_),
    .B1(net181),
    .Y(_11930_));
 sky130_fd_sc_hd__o21a_1 _20069_ (.A1(_11924_),
    .A2(_11925_),
    .B1(_11930_),
    .X(_11931_));
 sky130_fd_sc_hd__or3_1 _20070_ (.A(_11930_),
    .B(_11924_),
    .C(_11925_),
    .X(_11932_));
 sky130_fd_sc_hd__and2b_1 _20071_ (.A_N(_11931_),
    .B(_11932_),
    .X(_11933_));
 sky130_fd_sc_hd__o21ai_1 _20072_ (.A1(net1014),
    .A2(_11933_),
    .B1(net177),
    .Y(_11934_));
 sky130_fd_sc_hd__nor2_1 _20073_ (.A(\top0.cordic0.slte0.opA[10] ),
    .B(_11785_),
    .Y(_11935_));
 sky130_fd_sc_hd__a22o_1 _20074_ (.A1(net913),
    .A2(_11934_),
    .B1(_11935_),
    .B2(_11933_),
    .X(_00370_));
 sky130_fd_sc_hd__nor2_2 _20075_ (.A(net181),
    .B(_11519_),
    .Y(_11936_));
 sky130_fd_sc_hd__nand2_1 _20076_ (.A(_11428_),
    .B(_11936_),
    .Y(_11937_));
 sky130_fd_sc_hd__xnor2_1 _20077_ (.A(net203),
    .B(net187),
    .Y(_11938_));
 sky130_fd_sc_hd__nor2_1 _20078_ (.A(_11715_),
    .B(_11938_),
    .Y(_11939_));
 sky130_fd_sc_hd__xnor2_2 _20079_ (.A(_11937_),
    .B(_11939_),
    .Y(_11940_));
 sky130_fd_sc_hd__a21o_1 _20080_ (.A1(\top0.cordic0.slte0.opA[10] ),
    .A2(_11932_),
    .B1(_11931_),
    .X(_11941_));
 sky130_fd_sc_hd__nor2_1 _20081_ (.A(_11940_),
    .B(_11941_),
    .Y(_11942_));
 sky130_fd_sc_hd__and2_1 _20082_ (.A(_11940_),
    .B(_11941_),
    .X(_11943_));
 sky130_fd_sc_hd__nor2_1 _20083_ (.A(_11942_),
    .B(_11943_),
    .Y(_11944_));
 sky130_fd_sc_hd__o21ai_1 _20084_ (.A1(net1014),
    .A2(_11944_),
    .B1(net177),
    .Y(_11945_));
 sky130_fd_sc_hd__nor2_1 _20085_ (.A(\top0.cordic0.slte0.opA[11] ),
    .B(_11785_),
    .Y(_11946_));
 sky130_fd_sc_hd__a22o_1 _20086_ (.A1(\top0.cordic0.slte0.opA[11] ),
    .A2(_11945_),
    .B1(_11946_),
    .B2(_11944_),
    .X(_00371_));
 sky130_fd_sc_hd__nand2_1 _20087_ (.A(_11426_),
    .B(_11514_),
    .Y(_11947_));
 sky130_fd_sc_hd__o211a_1 _20088_ (.A1(_11714_),
    .A2(_11629_),
    .B1(_11936_),
    .C1(_11428_),
    .X(_11948_));
 sky130_fd_sc_hd__a41o_1 _20089_ (.A1(net194),
    .A2(net203),
    .A3(_11730_),
    .A4(_11947_),
    .B1(_11948_),
    .X(_11949_));
 sky130_fd_sc_hd__a21oi_1 _20090_ (.A1(_11940_),
    .A2(_11941_),
    .B1(\top0.cordic0.slte0.opA[11] ),
    .Y(_11950_));
 sky130_fd_sc_hd__nor2_1 _20091_ (.A(_11942_),
    .B(_11950_),
    .Y(_11951_));
 sky130_fd_sc_hd__xnor2_1 _20092_ (.A(_11949_),
    .B(_11951_),
    .Y(_11952_));
 sky130_fd_sc_hd__nor2_1 _20093_ (.A(_11857_),
    .B(_11952_),
    .Y(_11953_));
 sky130_fd_sc_hd__buf_4 _20094_ (.A(_11433_),
    .X(_11954_));
 sky130_fd_sc_hd__a21o_1 _20095_ (.A1(_11649_),
    .A2(_11952_),
    .B1(_11954_),
    .X(_11955_));
 sky130_fd_sc_hd__mux2_1 _20096_ (.A0(_11953_),
    .A1(_11955_),
    .S(\top0.cordic0.slte0.opA[12] ),
    .X(_11956_));
 sky130_fd_sc_hd__clkbuf_1 _20097_ (.A(_11956_),
    .X(_00372_));
 sky130_fd_sc_hd__a32o_1 _20098_ (.A1(net194),
    .A2(_11730_),
    .A3(_11808_),
    .B1(_11936_),
    .B2(_11804_),
    .X(_11957_));
 sky130_fd_sc_hd__nor2_1 _20099_ (.A(\top0.cordic0.slte0.opA[12] ),
    .B(_11949_),
    .Y(_11958_));
 sky130_fd_sc_hd__nand2_1 _20100_ (.A(\top0.cordic0.slte0.opA[12] ),
    .B(_11949_),
    .Y(_11959_));
 sky130_fd_sc_hd__o31a_1 _20101_ (.A1(_11942_),
    .A2(_11950_),
    .A3(_11958_),
    .B1(_11959_),
    .X(_11960_));
 sky130_fd_sc_hd__xor2_1 _20102_ (.A(_11957_),
    .B(_11960_),
    .X(_11961_));
 sky130_fd_sc_hd__nor2_1 _20103_ (.A(_11857_),
    .B(_11961_),
    .Y(_11962_));
 sky130_fd_sc_hd__a21o_1 _20104_ (.A1(_11649_),
    .A2(_11961_),
    .B1(_11954_),
    .X(_11963_));
 sky130_fd_sc_hd__mux2_1 _20105_ (.A0(_11962_),
    .A1(_11963_),
    .S(\top0.cordic0.slte0.opA[13] ),
    .X(_11964_));
 sky130_fd_sc_hd__clkbuf_1 _20106_ (.A(_11964_),
    .X(_00373_));
 sky130_fd_sc_hd__o21ba_1 _20107_ (.A1(\top0.cordic0.slte0.opA[13] ),
    .A2(_11957_),
    .B1_N(_11960_),
    .X(_11965_));
 sky130_fd_sc_hd__and2_1 _20108_ (.A(\top0.cordic0.slte0.opA[13] ),
    .B(_11957_),
    .X(_11966_));
 sky130_fd_sc_hd__or2_1 _20109_ (.A(_11965_),
    .B(_11966_),
    .X(_11967_));
 sky130_fd_sc_hd__and2_1 _20110_ (.A(_11426_),
    .B(_11775_),
    .X(_11968_));
 sky130_fd_sc_hd__and3_1 _20111_ (.A(_11730_),
    .B(_11519_),
    .C(_11810_),
    .X(_11969_));
 sky130_fd_sc_hd__a21o_1 _20112_ (.A1(_11515_),
    .A2(_11968_),
    .B1(_11969_),
    .X(_11970_));
 sky130_fd_sc_hd__xor2_1 _20113_ (.A(_11967_),
    .B(_11970_),
    .X(_11971_));
 sky130_fd_sc_hd__o21ai_1 _20114_ (.A1(net1014),
    .A2(_11971_),
    .B1(net177),
    .Y(_11972_));
 sky130_fd_sc_hd__nor2_1 _20115_ (.A(\top0.cordic0.slte0.opA[14] ),
    .B(_11857_),
    .Y(_11973_));
 sky130_fd_sc_hd__a22o_1 _20116_ (.A1(\top0.cordic0.slte0.opA[14] ),
    .A2(_11972_),
    .B1(_11973_),
    .B2(_11971_),
    .X(_00374_));
 sky130_fd_sc_hd__nor2_1 _20117_ (.A(_11413_),
    .B(_11515_),
    .Y(_11974_));
 sky130_fd_sc_hd__nor2_1 _20118_ (.A(\top0.cordic0.gm0.iter[4] ),
    .B(_11974_),
    .Y(_11975_));
 sky130_fd_sc_hd__nand2_1 _20119_ (.A(net177),
    .B(\top0.cordic0.slte0.opA[15] ),
    .Y(_11976_));
 sky130_fd_sc_hd__a211o_1 _20120_ (.A1(\top0.cordic0.slte0.opA[14] ),
    .A2(_11970_),
    .B1(_11966_),
    .C1(_11965_),
    .X(_11977_));
 sky130_fd_sc_hd__o21a_2 _20121_ (.A1(\top0.cordic0.slte0.opA[14] ),
    .A2(_11970_),
    .B1(_11977_),
    .X(_11978_));
 sky130_fd_sc_hd__mux2_1 _20122_ (.A0(net212),
    .A1(_11976_),
    .S(_11978_),
    .X(_11979_));
 sky130_fd_sc_hd__a211o_1 _20123_ (.A1(_11428_),
    .A2(_11947_),
    .B1(_11978_),
    .C1(_11976_),
    .X(_11980_));
 sky130_fd_sc_hd__nand2_1 _20124_ (.A(_11936_),
    .B(_11978_),
    .Y(_11981_));
 sky130_fd_sc_hd__a21o_1 _20125_ (.A1(net176),
    .A2(_11981_),
    .B1(net212),
    .X(_11982_));
 sky130_fd_sc_hd__o211a_1 _20126_ (.A1(_11975_),
    .A2(_11979_),
    .B1(_11980_),
    .C1(_11982_),
    .X(_00375_));
 sky130_fd_sc_hd__inv_2 _20127_ (.A(\top0.cordic0.slte0.opA[16] ),
    .Y(_11983_));
 sky130_fd_sc_hd__inv_2 _20128_ (.A(_11978_),
    .Y(_11984_));
 sky130_fd_sc_hd__nand2_1 _20129_ (.A(net212),
    .B(_11947_),
    .Y(_11985_));
 sky130_fd_sc_hd__nor2_1 _20130_ (.A(\top0.cordic0.slte0.opA[14] ),
    .B(_11775_),
    .Y(_11986_));
 sky130_fd_sc_hd__a21oi_1 _20131_ (.A1(\top0.cordic0.slte0.opA[14] ),
    .A2(_11775_),
    .B1(_11967_),
    .Y(_11987_));
 sky130_fd_sc_hd__o21ai_1 _20132_ (.A1(_11986_),
    .A2(_11987_),
    .B1(_11936_),
    .Y(_11988_));
 sky130_fd_sc_hd__or2_1 _20133_ (.A(_11426_),
    .B(net212),
    .X(_11989_));
 sky130_fd_sc_hd__a21o_1 _20134_ (.A1(_11985_),
    .A2(_11989_),
    .B1(_11428_),
    .X(_11990_));
 sky130_fd_sc_hd__o221a_1 _20135_ (.A1(_11984_),
    .A2(_11985_),
    .B1(_11988_),
    .B2(net212),
    .C1(_11990_),
    .X(_11991_));
 sky130_fd_sc_hd__a41o_1 _20136_ (.A1(net212),
    .A2(_11434_),
    .A3(_11947_),
    .A4(_11978_),
    .B1(\top0.cordic0.slte0.opA[16] ),
    .X(_11992_));
 sky130_fd_sc_hd__and3_1 _20137_ (.A(net212),
    .B(_11413_),
    .C(_11519_),
    .X(_11993_));
 sky130_fd_sc_hd__or2_1 _20138_ (.A(_11967_),
    .B(_11968_),
    .X(_11994_));
 sky130_fd_sc_hd__a21o_1 _20139_ (.A1(_11967_),
    .A2(_11968_),
    .B1(\top0.cordic0.slte0.opA[14] ),
    .X(_11995_));
 sky130_fd_sc_hd__a211oi_1 _20140_ (.A1(_11994_),
    .A2(_11995_),
    .B1(net212),
    .C1(_11519_),
    .Y(_11996_));
 sky130_fd_sc_hd__nor2_1 _20141_ (.A(_11433_),
    .B(net180),
    .Y(_11997_));
 sky130_fd_sc_hd__o21a_1 _20142_ (.A1(_11993_),
    .A2(_11996_),
    .B1(_11997_),
    .X(_11998_));
 sky130_fd_sc_hd__o32a_1 _20143_ (.A1(net1020),
    .A2(_11983_),
    .A3(_11991_),
    .B1(_11992_),
    .B2(_11998_),
    .X(_00376_));
 sky130_fd_sc_hd__a32o_1 _20144_ (.A1(_11983_),
    .A2(_11515_),
    .A3(_11997_),
    .B1(\top0.cordic0.slte0.opA[17] ),
    .B2(_11649_),
    .X(_11999_));
 sky130_fd_sc_hd__or3b_1 _20145_ (.A(net180),
    .B(_11974_),
    .C_N(net212),
    .X(_12000_));
 sky130_fd_sc_hd__o21ai_1 _20146_ (.A1(net212),
    .A2(_11936_),
    .B1(_11978_),
    .Y(_12001_));
 sky130_fd_sc_hd__a21o_1 _20147_ (.A1(_11983_),
    .A2(_11649_),
    .B1(_11954_),
    .X(_12002_));
 sky130_fd_sc_hd__a32o_1 _20148_ (.A1(_11999_),
    .A2(_12000_),
    .A3(_12001_),
    .B1(_12002_),
    .B2(\top0.cordic0.slte0.opA[17] ),
    .X(_00377_));
 sky130_fd_sc_hd__nand2_4 _20149_ (.A(_11433_),
    .B(\top0.cordic0.in_valid ),
    .Y(_12003_));
 sky130_fd_sc_hd__clkbuf_4 _20150_ (.A(_12003_),
    .X(_12004_));
 sky130_fd_sc_hd__mux2_1 _20151_ (.A0(\spi0.data_packed[14] ),
    .A1(\top0.cordic0.domain[0] ),
    .S(_12004_),
    .X(_12005_));
 sky130_fd_sc_hd__clkbuf_1 _20152_ (.A(_12005_),
    .X(_00378_));
 sky130_fd_sc_hd__clkbuf_4 _20153_ (.A(_12003_),
    .X(_12006_));
 sky130_fd_sc_hd__mux2_1 _20154_ (.A0(\spi0.data_packed[15] ),
    .A1(net211),
    .S(_12006_),
    .X(_12007_));
 sky130_fd_sc_hd__clkbuf_1 _20155_ (.A(_12007_),
    .X(_00379_));
 sky130_fd_sc_hd__a21oi_1 _20156_ (.A1(net207),
    .A2(net206),
    .B1(net209),
    .Y(_12008_));
 sky130_fd_sc_hd__inv_2 _20157_ (.A(net207),
    .Y(_12009_));
 sky130_fd_sc_hd__or2_1 _20158_ (.A(_12009_),
    .B(net208),
    .X(_12010_));
 sky130_fd_sc_hd__mux2_1 _20159_ (.A0(_05437_),
    .A1(\top0.svm0.out_valid ),
    .S(net206),
    .X(_12011_));
 sky130_fd_sc_hd__nand2_1 _20160_ (.A(net209),
    .B(net206),
    .Y(_12012_));
 sky130_fd_sc_hd__or2_1 _20161_ (.A(\top0.state[1] ),
    .B(_12012_),
    .X(_12013_));
 sky130_fd_sc_hd__buf_2 _20162_ (.A(_12013_),
    .X(_12014_));
 sky130_fd_sc_hd__and2b_1 _20163_ (.A_N(net205),
    .B(net208),
    .X(_12015_));
 sky130_fd_sc_hd__nand2_1 _20164_ (.A(net207),
    .B(_12015_),
    .Y(_12016_));
 sky130_fd_sc_hd__or2_2 _20165_ (.A(net205),
    .B(_05425_),
    .X(_12017_));
 sky130_fd_sc_hd__inv_2 _20166_ (.A(_12017_),
    .Y(_12018_));
 sky130_fd_sc_hd__or2_2 _20167_ (.A(net207),
    .B(net208),
    .X(_12019_));
 sky130_fd_sc_hd__a21o_1 _20168_ (.A1(net205),
    .A2(_05437_),
    .B1(_12019_),
    .X(_12020_));
 sky130_fd_sc_hd__a21o_1 _20169_ (.A1(\top0.clarke_done ),
    .A2(\top0.cordic0.out_valid ),
    .B1(_05437_),
    .X(_12021_));
 sky130_fd_sc_hd__or2_1 _20170_ (.A(\top0.cordic0.out_valid ),
    .B(\top0.cordic_done ),
    .X(_12022_));
 sky130_fd_sc_hd__a21oi_1 _20171_ (.A1(_12021_),
    .A2(_12022_),
    .B1(net207),
    .Y(_12023_));
 sky130_fd_sc_hd__nand2_1 _20172_ (.A(_12015_),
    .B(_12023_),
    .Y(_12024_));
 sky130_fd_sc_hd__o221a_1 _20173_ (.A1(\top0.pid_d.out_valid ),
    .A2(_12016_),
    .B1(_12018_),
    .B2(_12020_),
    .C1(_12024_),
    .X(_12025_));
 sky130_fd_sc_hd__o221a_2 _20174_ (.A1(_12010_),
    .A2(_12011_),
    .B1(_12014_),
    .B2(_05439_),
    .C1(_12025_),
    .X(_12026_));
 sky130_fd_sc_hd__mux2_1 _20175_ (.A0(net209),
    .A1(_12008_),
    .S(_12026_),
    .X(_12027_));
 sky130_fd_sc_hd__clkbuf_1 _20176_ (.A(_12027_),
    .X(_00380_));
 sky130_fd_sc_hd__or2_1 _20177_ (.A(net209),
    .B(net206),
    .X(_12028_));
 sky130_fd_sc_hd__a21oi_1 _20178_ (.A1(_12026_),
    .A2(_12028_),
    .B1(_12009_),
    .Y(_12029_));
 sky130_fd_sc_hd__a31o_1 _20179_ (.A1(_12009_),
    .A2(net208),
    .A3(_12026_),
    .B1(_12029_),
    .X(_00381_));
 sky130_fd_sc_hd__nand2b_2 _20180_ (.A_N(net205),
    .B(net208),
    .Y(_12030_));
 sky130_fd_sc_hd__nor2_2 _20181_ (.A(_12009_),
    .B(_12030_),
    .Y(_12031_));
 sky130_fd_sc_hd__clkbuf_4 _20182_ (.A(_12031_),
    .X(_12032_));
 sky130_fd_sc_hd__nand2_1 _20183_ (.A(\top0.state[1] ),
    .B(_12026_),
    .Y(_12033_));
 sky130_fd_sc_hd__a22o_1 _20184_ (.A1(_12032_),
    .A2(_12026_),
    .B1(_12033_),
    .B2(net206),
    .X(_00382_));
 sky130_fd_sc_hd__buf_6 _20185_ (.A(_12004_),
    .X(_12034_));
 sky130_fd_sc_hd__nand2_2 _20186_ (.A(net176),
    .B(_11429_),
    .Y(_12035_));
 sky130_fd_sc_hd__buf_6 _20187_ (.A(_12035_),
    .X(_12036_));
 sky130_fd_sc_hd__buf_6 _20188_ (.A(_12036_),
    .X(_12037_));
 sky130_fd_sc_hd__xnor2_2 _20189_ (.A(net245),
    .B(net237),
    .Y(_12038_));
 sky130_fd_sc_hd__nor2b_2 _20190_ (.A(net259),
    .B_N(net255),
    .Y(_12039_));
 sky130_fd_sc_hd__xnor2_4 _20191_ (.A(net252),
    .B(_12039_),
    .Y(_12040_));
 sky130_fd_sc_hd__xor2_1 _20192_ (.A(_12038_),
    .B(_12040_),
    .X(_12041_));
 sky130_fd_sc_hd__xnor2_4 _20193_ (.A(net252),
    .B(net240),
    .Y(_12042_));
 sky130_fd_sc_hd__or2_1 _20194_ (.A(net258),
    .B(net253),
    .X(_12043_));
 sky130_fd_sc_hd__a21boi_1 _20195_ (.A1(net253),
    .A2(_12042_),
    .B1_N(_12043_),
    .Y(_12044_));
 sky130_fd_sc_hd__and2_1 _20196_ (.A(net262),
    .B(net257),
    .X(_12045_));
 sky130_fd_sc_hd__o21bai_2 _20197_ (.A1(_12042_),
    .A2(_12045_),
    .B1_N(net267),
    .Y(_12046_));
 sky130_fd_sc_hd__nand2_2 _20198_ (.A(net299),
    .B(net296),
    .Y(_12047_));
 sky130_fd_sc_hd__or2b_1 _20199_ (.A(net269),
    .B_N(net283),
    .X(_12048_));
 sky130_fd_sc_hd__and2b_2 _20200_ (.A_N(net283),
    .B(net276),
    .X(_12049_));
 sky130_fd_sc_hd__nor2_1 _20201_ (.A(net276),
    .B(net269),
    .Y(_12050_));
 sky130_fd_sc_hd__a221o_1 _20202_ (.A1(_12047_),
    .A2(_12048_),
    .B1(_12049_),
    .B2(net269),
    .C1(_12050_),
    .X(_12051_));
 sky130_fd_sc_hd__and3_1 _20203_ (.A(_12044_),
    .B(_12046_),
    .C(_12051_),
    .X(_12052_));
 sky130_fd_sc_hd__a21oi_1 _20204_ (.A1(_12044_),
    .A2(_12046_),
    .B1(_12051_),
    .Y(_12053_));
 sky130_fd_sc_hd__or3_1 _20205_ (.A(_12041_),
    .B(_12052_),
    .C(_12053_),
    .X(_12054_));
 sky130_fd_sc_hd__o21ai_1 _20206_ (.A1(_12052_),
    .A2(_12053_),
    .B1(_12041_),
    .Y(_12055_));
 sky130_fd_sc_hd__xnor2_4 _20207_ (.A(net269),
    .B(_12049_),
    .Y(_12056_));
 sky130_fd_sc_hd__nand2b_2 _20208_ (.A_N(net296),
    .B(net289),
    .Y(_12057_));
 sky130_fd_sc_hd__xnor2_1 _20209_ (.A(net299),
    .B(_12056_),
    .Y(_12058_));
 sky130_fd_sc_hd__nor2b_2 _20210_ (.A(net290),
    .B_N(net296),
    .Y(_12059_));
 sky130_fd_sc_hd__a2bb2o_1 _20211_ (.A1_N(_12056_),
    .A2_N(_12057_),
    .B1(_12058_),
    .B2(_12059_),
    .X(_12060_));
 sky130_fd_sc_hd__xnor2_1 _20212_ (.A(net304),
    .B(net281),
    .Y(_12061_));
 sky130_fd_sc_hd__nor2_1 _20213_ (.A(_11550_),
    .B(_12061_),
    .Y(_12062_));
 sky130_fd_sc_hd__nand2_1 _20214_ (.A(_11550_),
    .B(_12061_),
    .Y(_12063_));
 sky130_fd_sc_hd__and2b_1 _20215_ (.A_N(_12062_),
    .B(_12063_),
    .X(_12064_));
 sky130_fd_sc_hd__nand2_4 _20216_ (.A(net297),
    .B(net290),
    .Y(_12065_));
 sky130_fd_sc_hd__and2b_2 _20217_ (.A_N(net279),
    .B(net269),
    .X(_12066_));
 sky130_fd_sc_hd__xnor2_4 _20218_ (.A(net264),
    .B(_12066_),
    .Y(_12067_));
 sky130_fd_sc_hd__xnor2_2 _20219_ (.A(_12065_),
    .B(_12067_),
    .Y(_12068_));
 sky130_fd_sc_hd__xnor2_2 _20220_ (.A(_12064_),
    .B(_12068_),
    .Y(_12069_));
 sky130_fd_sc_hd__a31o_1 _20221_ (.A1(_12054_),
    .A2(_12055_),
    .A3(_12060_),
    .B1(_12069_),
    .X(_12070_));
 sky130_fd_sc_hd__a21o_1 _20222_ (.A1(_12054_),
    .A2(_12055_),
    .B1(_12060_),
    .X(_12071_));
 sky130_fd_sc_hd__clkinv_4 _20223_ (.A(net221),
    .Y(_12072_));
 sky130_fd_sc_hd__nand2_1 _20224_ (.A(net247),
    .B(net234),
    .Y(_12073_));
 sky130_fd_sc_hd__xnor2_2 _20225_ (.A(_12072_),
    .B(_12073_),
    .Y(_12074_));
 sky130_fd_sc_hd__nand2_2 _20226_ (.A(net252),
    .B(net240),
    .Y(_12075_));
 sky130_fd_sc_hd__nor3_1 _20227_ (.A(_11758_),
    .B(_12074_),
    .C(_12075_),
    .Y(_12076_));
 sky130_fd_sc_hd__o21ai_2 _20228_ (.A1(_11758_),
    .A2(_12075_),
    .B1(_12074_),
    .Y(_12077_));
 sky130_fd_sc_hd__or2b_1 _20229_ (.A(_12076_),
    .B_N(_12077_),
    .X(_12078_));
 sky130_fd_sc_hd__a21bo_1 _20230_ (.A1(_12044_),
    .A2(_12046_),
    .B1_N(_12051_),
    .X(_12079_));
 sky130_fd_sc_hd__nand2_1 _20231_ (.A(net253),
    .B(_12042_),
    .Y(_12080_));
 sky130_fd_sc_hd__and4b_1 _20232_ (.A_N(_12051_),
    .B(_12046_),
    .C(_12080_),
    .D(_12043_),
    .X(_12081_));
 sky130_fd_sc_hd__a21o_1 _20233_ (.A1(_12041_),
    .A2(_12079_),
    .B1(_12081_),
    .X(_12082_));
 sky130_fd_sc_hd__xnor2_2 _20234_ (.A(_12078_),
    .B(_12082_),
    .Y(_12083_));
 sky130_fd_sc_hd__a21oi_2 _20235_ (.A1(_12070_),
    .A2(_12071_),
    .B1(_12083_),
    .Y(_12084_));
 sky130_fd_sc_hd__nor2_1 _20236_ (.A(net253),
    .B(net249),
    .Y(_12085_));
 sky130_fd_sc_hd__a21oi_1 _20237_ (.A1(net249),
    .A2(_12038_),
    .B1(_12085_),
    .Y(_12086_));
 sky130_fd_sc_hd__and2_1 _20238_ (.A(net253),
    .B(net249),
    .X(_12087_));
 sky130_fd_sc_hd__o21ai_1 _20239_ (.A1(_12087_),
    .A2(_12038_),
    .B1(_11653_),
    .Y(_12088_));
 sky130_fd_sc_hd__or2b_1 _20240_ (.A(net264),
    .B_N(net279),
    .X(_12089_));
 sky130_fd_sc_hd__nor2_1 _20241_ (.A(net270),
    .B(net264),
    .Y(_12090_));
 sky130_fd_sc_hd__a221o_2 _20242_ (.A1(net264),
    .A2(_12066_),
    .B1(_12089_),
    .B2(_12065_),
    .C1(_12090_),
    .X(_12091_));
 sky130_fd_sc_hd__nand3_1 _20243_ (.A(_12086_),
    .B(_12088_),
    .C(_12091_),
    .Y(_12092_));
 sky130_fd_sc_hd__a21o_1 _20244_ (.A1(_12086_),
    .A2(_12088_),
    .B1(_12091_),
    .X(_12093_));
 sky130_fd_sc_hd__nor2b_2 _20245_ (.A(net255),
    .B_N(net250),
    .Y(_12094_));
 sky130_fd_sc_hd__xnor2_4 _20246_ (.A(net244),
    .B(_12094_),
    .Y(_12095_));
 sky130_fd_sc_hd__xnor2_4 _20247_ (.A(net240),
    .B(net230),
    .Y(_12096_));
 sky130_fd_sc_hd__xnor2_2 _20248_ (.A(_12095_),
    .B(_12096_),
    .Y(_12097_));
 sky130_fd_sc_hd__a21bo_1 _20249_ (.A1(_12092_),
    .A2(_12093_),
    .B1_N(_12097_),
    .X(_12098_));
 sky130_fd_sc_hd__nand3b_1 _20250_ (.A_N(_12097_),
    .B(_12092_),
    .C(_12093_),
    .Y(_12099_));
 sky130_fd_sc_hd__xnor2_4 _20251_ (.A(net301),
    .B(net276),
    .Y(_12100_));
 sky130_fd_sc_hd__nor2b_2 _20252_ (.A(net271),
    .B_N(net265),
    .Y(_12101_));
 sky130_fd_sc_hd__xnor2_4 _20253_ (.A(net258),
    .B(_12101_),
    .Y(_12102_));
 sky130_fd_sc_hd__xnor2_2 _20254_ (.A(_12100_),
    .B(_12102_),
    .Y(_12103_));
 sky130_fd_sc_hd__inv_2 _20255_ (.A(_12103_),
    .Y(_12104_));
 sky130_fd_sc_hd__a21o_1 _20256_ (.A1(_12098_),
    .A2(_12099_),
    .B1(_12104_),
    .X(_12105_));
 sky130_fd_sc_hd__nand3_1 _20257_ (.A(_12098_),
    .B(_12099_),
    .C(_12104_),
    .Y(_12106_));
 sky130_fd_sc_hd__nand2_1 _20258_ (.A(net305),
    .B(net290),
    .Y(_12107_));
 sky130_fd_sc_hd__nor2b_4 _20259_ (.A(net290),
    .B_N(net284),
    .Y(_12108_));
 sky130_fd_sc_hd__and2_1 _20260_ (.A(net305),
    .B(net290),
    .X(_12109_));
 sky130_fd_sc_hd__a32oi_1 _20261_ (.A1(_11408_),
    .A2(_12067_),
    .A3(_12108_),
    .B1(_12109_),
    .B2(_11571_),
    .Y(_12110_));
 sky130_fd_sc_hd__a211o_1 _20262_ (.A1(_11408_),
    .A2(_11550_),
    .B1(net282),
    .C1(_12068_),
    .X(_12111_));
 sky130_fd_sc_hd__o211a_1 _20263_ (.A1(_12068_),
    .A2(_12107_),
    .B1(_12110_),
    .C1(_12111_),
    .X(_12112_));
 sky130_fd_sc_hd__a21oi_1 _20264_ (.A1(_12105_),
    .A2(_12106_),
    .B1(_12112_),
    .Y(_12113_));
 sky130_fd_sc_hd__and3_1 _20265_ (.A(_12112_),
    .B(_12105_),
    .C(_12106_),
    .X(_12114_));
 sky130_fd_sc_hd__nor2_2 _20266_ (.A(_12113_),
    .B(_12114_),
    .Y(_12115_));
 sky130_fd_sc_hd__and3_1 _20267_ (.A(_12083_),
    .B(_12070_),
    .C(_12071_),
    .X(_12116_));
 sky130_fd_sc_hd__nor2_1 _20268_ (.A(_12115_),
    .B(_12116_),
    .Y(_12117_));
 sky130_fd_sc_hd__nand2_1 _20269_ (.A(net289),
    .B(_11571_),
    .Y(_12118_));
 sky130_fd_sc_hd__o21a_1 _20270_ (.A1(net289),
    .A2(_12102_),
    .B1(_12118_),
    .X(_12119_));
 sky130_fd_sc_hd__o2bb2a_1 _20271_ (.A1_N(_12108_),
    .A2_N(_12100_),
    .B1(_12102_),
    .B2(_12118_),
    .X(_12120_));
 sky130_fd_sc_hd__o21ai_1 _20272_ (.A1(_12100_),
    .A2(_12119_),
    .B1(_12120_),
    .Y(_12121_));
 sky130_fd_sc_hd__xnor2_1 _20273_ (.A(net289),
    .B(_12102_),
    .Y(_12122_));
 sky130_fd_sc_hd__nor3_1 _20274_ (.A(net283),
    .B(_12100_),
    .C(_12102_),
    .Y(_12123_));
 sky130_fd_sc_hd__a31o_1 _20275_ (.A1(net283),
    .A2(_12100_),
    .A3(_12122_),
    .B1(_12123_),
    .X(_12124_));
 sky130_fd_sc_hd__a21o_1 _20276_ (.A1(net304),
    .A2(_12121_),
    .B1(_12124_),
    .X(_12125_));
 sky130_fd_sc_hd__nand2b_4 _20277_ (.A_N(net267),
    .B(\top0.cordic0.vec[0][8] ),
    .Y(_12126_));
 sky130_fd_sc_hd__xnor2_4 _20278_ (.A(_11672_),
    .B(_12126_),
    .Y(_12127_));
 sky130_fd_sc_hd__or2b_1 _20279_ (.A(net276),
    .B_N(net283),
    .X(_12128_));
 sky130_fd_sc_hd__or3b_1 _20280_ (.A(net299),
    .B(net283),
    .C_N(net276),
    .X(_12129_));
 sky130_fd_sc_hd__o21a_1 _20281_ (.A1(_11437_),
    .A2(_12128_),
    .B1(_12129_),
    .X(_12130_));
 sky130_fd_sc_hd__xnor2_2 _20282_ (.A(net296),
    .B(net269),
    .Y(_12131_));
 sky130_fd_sc_hd__xnor2_1 _20283_ (.A(_12130_),
    .B(_12131_),
    .Y(_12132_));
 sky130_fd_sc_hd__xnor2_2 _20284_ (.A(_12127_),
    .B(_12132_),
    .Y(_12133_));
 sky130_fd_sc_hd__nor2b_2 _20285_ (.A(net252),
    .B_N(net246),
    .Y(_12134_));
 sky130_fd_sc_hd__xnor2_4 _20286_ (.A(net238),
    .B(_12134_),
    .Y(_12135_));
 sky130_fd_sc_hd__xnor2_2 _20287_ (.A(net234),
    .B(net226),
    .Y(_12136_));
 sky130_fd_sc_hd__xnor2_2 _20288_ (.A(_12135_),
    .B(_12136_),
    .Y(_12137_));
 sky130_fd_sc_hd__nor2_1 _20289_ (.A(net250),
    .B(net244),
    .Y(_12138_));
 sky130_fd_sc_hd__a21oi_2 _20290_ (.A1(net245),
    .A2(_12096_),
    .B1(_12138_),
    .Y(_12139_));
 sky130_fd_sc_hd__and2_1 _20291_ (.A(net252),
    .B(net246),
    .X(_12140_));
 sky130_fd_sc_hd__o21ai_1 _20292_ (.A1(_12096_),
    .A2(_12140_),
    .B1(_11672_),
    .Y(_12141_));
 sky130_fd_sc_hd__nand2_2 _20293_ (.A(net290),
    .B(net282),
    .Y(_12142_));
 sky130_fd_sc_hd__or2b_1 _20294_ (.A(net261),
    .B_N(net269),
    .X(_12143_));
 sky130_fd_sc_hd__nor2_1 _20295_ (.A(net264),
    .B(net261),
    .Y(_12144_));
 sky130_fd_sc_hd__a221o_1 _20296_ (.A1(net258),
    .A2(_12101_),
    .B1(_12142_),
    .B2(_12143_),
    .C1(_12144_),
    .X(_12145_));
 sky130_fd_sc_hd__a21o_1 _20297_ (.A1(_12139_),
    .A2(_12141_),
    .B1(_12145_),
    .X(_12146_));
 sky130_fd_sc_hd__nand3_1 _20298_ (.A(_12139_),
    .B(_12141_),
    .C(_12145_),
    .Y(_12147_));
 sky130_fd_sc_hd__nand3_2 _20299_ (.A(_12137_),
    .B(_12146_),
    .C(_12147_),
    .Y(_12148_));
 sky130_fd_sc_hd__a21o_1 _20300_ (.A1(_12146_),
    .A2(_12147_),
    .B1(_12137_),
    .X(_12149_));
 sky130_fd_sc_hd__nand3_2 _20301_ (.A(_12133_),
    .B(_12148_),
    .C(_12149_),
    .Y(_12150_));
 sky130_fd_sc_hd__a21o_1 _20302_ (.A1(_12148_),
    .A2(_12149_),
    .B1(_12133_),
    .X(_12151_));
 sky130_fd_sc_hd__nand2_1 _20303_ (.A(_12150_),
    .B(_12151_),
    .Y(_12152_));
 sky130_fd_sc_hd__xnor2_1 _20304_ (.A(_12125_),
    .B(_12152_),
    .Y(_12153_));
 sky130_fd_sc_hd__nand2_1 _20305_ (.A(_12098_),
    .B(_12099_),
    .Y(_12154_));
 sky130_fd_sc_hd__or3b_1 _20306_ (.A(_12062_),
    .B(_12068_),
    .C_N(_12063_),
    .X(_12155_));
 sky130_fd_sc_hd__nand2b_2 _20307_ (.A_N(net289),
    .B(net282),
    .Y(_12156_));
 sky130_fd_sc_hd__o22a_1 _20308_ (.A1(net304),
    .A2(_12156_),
    .B1(_12107_),
    .B2(net280),
    .X(_12157_));
 sky130_fd_sc_hd__xnor2_1 _20309_ (.A(_12103_),
    .B(_12157_),
    .Y(_12158_));
 sky130_fd_sc_hd__nor2_1 _20310_ (.A(_12155_),
    .B(_12158_),
    .Y(_12159_));
 sky130_fd_sc_hd__nand2_1 _20311_ (.A(_12155_),
    .B(_12158_),
    .Y(_12160_));
 sky130_fd_sc_hd__o21a_4 _20312_ (.A1(_12154_),
    .A2(_12159_),
    .B1(_12160_),
    .X(_12161_));
 sky130_fd_sc_hd__o2bb2a_1 _20313_ (.A1_N(_12086_),
    .A2_N(_12088_),
    .B1(_12091_),
    .B2(_12097_),
    .X(_12162_));
 sky130_fd_sc_hd__a21oi_4 _20314_ (.A1(_12097_),
    .A2(_12091_),
    .B1(_12162_),
    .Y(_12163_));
 sky130_fd_sc_hd__nor2_1 _20315_ (.A(_12072_),
    .B(_12073_),
    .Y(_12164_));
 sky130_fd_sc_hd__nand2_2 _20316_ (.A(net239),
    .B(net230),
    .Y(_12165_));
 sky130_fd_sc_hd__xnor2_2 _20317_ (.A(net214),
    .B(_12165_),
    .Y(_12166_));
 sky130_fd_sc_hd__xnor2_1 _20318_ (.A(_12164_),
    .B(_12166_),
    .Y(_12167_));
 sky130_fd_sc_hd__xnor2_1 _20319_ (.A(_12163_),
    .B(_12167_),
    .Y(_12168_));
 sky130_fd_sc_hd__xnor2_1 _20320_ (.A(_12161_),
    .B(_12168_),
    .Y(_12169_));
 sky130_fd_sc_hd__xnor2_2 _20321_ (.A(_12153_),
    .B(_12169_),
    .Y(_12170_));
 sky130_fd_sc_hd__a21oi_2 _20322_ (.A1(_12077_),
    .A2(_12082_),
    .B1(_12076_),
    .Y(_12171_));
 sky130_fd_sc_hd__o22a_1 _20323_ (.A1(_12084_),
    .A2(_12117_),
    .B1(_12170_),
    .B2(_12171_),
    .X(_12172_));
 sky130_fd_sc_hd__and2_1 _20324_ (.A(_12170_),
    .B(_12171_),
    .X(_12173_));
 sky130_fd_sc_hd__inv_2 _20325_ (.A(_12163_),
    .Y(_12174_));
 sky130_fd_sc_hd__a21oi_2 _20326_ (.A1(net304),
    .A2(_12121_),
    .B1(_12124_),
    .Y(_12175_));
 sky130_fd_sc_hd__a211o_1 _20327_ (.A1(_12150_),
    .A2(_12151_),
    .B1(_12166_),
    .C1(_12175_),
    .X(_12176_));
 sky130_fd_sc_hd__xnor2_1 _20328_ (.A(_11787_),
    .B(_12165_),
    .Y(_12177_));
 sky130_fd_sc_hd__nand4_2 _20329_ (.A(_12175_),
    .B(_12150_),
    .C(_12151_),
    .D(_12177_),
    .Y(_12178_));
 sky130_fd_sc_hd__nand2_1 _20330_ (.A(_12176_),
    .B(_12178_),
    .Y(_12179_));
 sky130_fd_sc_hd__buf_6 _20331_ (.A(_12072_),
    .X(_12180_));
 sky130_fd_sc_hd__or2_1 _20332_ (.A(_12180_),
    .B(_12073_),
    .X(_12181_));
 sky130_fd_sc_hd__a211o_1 _20333_ (.A1(_12150_),
    .A2(_12151_),
    .B1(_12177_),
    .C1(_12125_),
    .X(_12182_));
 sky130_fd_sc_hd__nand4_2 _20334_ (.A(_12125_),
    .B(_12150_),
    .C(_12151_),
    .D(_12166_),
    .Y(_12183_));
 sky130_fd_sc_hd__and3_1 _20335_ (.A(_12181_),
    .B(_12182_),
    .C(_12183_),
    .X(_12184_));
 sky130_fd_sc_hd__a21o_1 _20336_ (.A1(_12182_),
    .A2(_12183_),
    .B1(_12181_),
    .X(_12185_));
 sky130_fd_sc_hd__o311a_1 _20337_ (.A1(_12174_),
    .A2(_12179_),
    .A3(_12184_),
    .B1(_12185_),
    .C1(_12161_),
    .X(_12186_));
 sky130_fd_sc_hd__nand2_2 _20338_ (.A(_12182_),
    .B(_12183_),
    .Y(_12187_));
 sky130_fd_sc_hd__and3_1 _20339_ (.A(_12164_),
    .B(_12176_),
    .C(_12178_),
    .X(_12188_));
 sky130_fd_sc_hd__a21o_1 _20340_ (.A1(_12176_),
    .A2(_12178_),
    .B1(_12164_),
    .X(_12189_));
 sky130_fd_sc_hd__inv_2 _20341_ (.A(_12161_),
    .Y(_12190_));
 sky130_fd_sc_hd__o311a_1 _20342_ (.A1(_12163_),
    .A2(_12187_),
    .A3(_12188_),
    .B1(_12189_),
    .C1(_12190_),
    .X(_12191_));
 sky130_fd_sc_hd__nor2_1 _20343_ (.A(_12174_),
    .B(_12181_),
    .Y(_12192_));
 sky130_fd_sc_hd__nand2_1 _20344_ (.A(_12187_),
    .B(_12192_),
    .Y(_12193_));
 sky130_fd_sc_hd__or2_2 _20345_ (.A(_12163_),
    .B(_12164_),
    .X(_12194_));
 sky130_fd_sc_hd__a21o_1 _20346_ (.A1(_12176_),
    .A2(_12178_),
    .B1(_12194_),
    .X(_12195_));
 sky130_fd_sc_hd__o211ai_1 _20347_ (.A1(_12186_),
    .A2(_12191_),
    .B1(_12193_),
    .C1(_12195_),
    .Y(_12196_));
 sky130_fd_sc_hd__nor2_1 _20348_ (.A(net246),
    .B(net238),
    .Y(_12197_));
 sky130_fd_sc_hd__a21oi_1 _20349_ (.A1(net238),
    .A2(_12136_),
    .B1(_12197_),
    .Y(_12198_));
 sky130_fd_sc_hd__and2_1 _20350_ (.A(net247),
    .B(net238),
    .X(_12199_));
 sky130_fd_sc_hd__o21ai_1 _20351_ (.A1(_12136_),
    .A2(_12199_),
    .B1(_11689_),
    .Y(_12200_));
 sky130_fd_sc_hd__and2_1 _20352_ (.A(net283),
    .B(net276),
    .X(_12201_));
 sky130_fd_sc_hd__and2b_1 _20353_ (.A_N(net253),
    .B(net267),
    .X(_12202_));
 sky130_fd_sc_hd__o221a_1 _20354_ (.A1(_11672_),
    .A2(_12126_),
    .B1(_12201_),
    .B2(_12202_),
    .C1(_12043_),
    .X(_12203_));
 sky130_fd_sc_hd__a21o_1 _20355_ (.A1(_12198_),
    .A2(_12200_),
    .B1(_12203_),
    .X(_12204_));
 sky130_fd_sc_hd__nand3_1 _20356_ (.A(_12198_),
    .B(_12200_),
    .C(_12203_),
    .Y(_12205_));
 sky130_fd_sc_hd__xor2_2 _20357_ (.A(net229),
    .B(net221),
    .X(_12206_));
 sky130_fd_sc_hd__nor2b_2 _20358_ (.A(net246),
    .B_N(net239),
    .Y(_12207_));
 sky130_fd_sc_hd__xnor2_4 _20359_ (.A(net234),
    .B(_12207_),
    .Y(_12208_));
 sky130_fd_sc_hd__xnor2_2 _20360_ (.A(_12206_),
    .B(_12208_),
    .Y(_12209_));
 sky130_fd_sc_hd__a21oi_1 _20361_ (.A1(_12204_),
    .A2(_12205_),
    .B1(_12209_),
    .Y(_12210_));
 sky130_fd_sc_hd__and3_1 _20362_ (.A(_12209_),
    .B(_12204_),
    .C(_12205_),
    .X(_12211_));
 sky130_fd_sc_hd__or2b_1 _20363_ (.A(net271),
    .B_N(net277),
    .X(_12212_));
 sky130_fd_sc_hd__or3b_1 _20364_ (.A(net296),
    .B(net277),
    .C_N(net269),
    .X(_12213_));
 sky130_fd_sc_hd__o21a_1 _20365_ (.A1(_11525_),
    .A2(_12212_),
    .B1(_12213_),
    .X(_12214_));
 sky130_fd_sc_hd__xnor2_2 _20366_ (.A(net291),
    .B(net265),
    .Y(_12215_));
 sky130_fd_sc_hd__xnor2_1 _20367_ (.A(_12214_),
    .B(_12215_),
    .Y(_12216_));
 sky130_fd_sc_hd__xnor2_2 _20368_ (.A(_12040_),
    .B(_12216_),
    .Y(_12217_));
 sky130_fd_sc_hd__or3b_1 _20369_ (.A(_12210_),
    .B(_12211_),
    .C_N(_12217_),
    .X(_12218_));
 sky130_fd_sc_hd__o21bai_1 _20370_ (.A1(_12210_),
    .A2(_12211_),
    .B1_N(_12217_),
    .Y(_12219_));
 sky130_fd_sc_hd__o2bb2a_1 _20371_ (.A1_N(_12049_),
    .A2_N(_12131_),
    .B1(_12127_),
    .B2(_12128_),
    .X(_12220_));
 sky130_fd_sc_hd__or2_1 _20372_ (.A(_11437_),
    .B(_12131_),
    .X(_12221_));
 sky130_fd_sc_hd__o21a_1 _20373_ (.A1(net283),
    .A2(_12127_),
    .B1(_12128_),
    .X(_12222_));
 sky130_fd_sc_hd__o22a_1 _20374_ (.A1(_11438_),
    .A2(_12220_),
    .B1(_12221_),
    .B2(_12222_),
    .X(_12223_));
 sky130_fd_sc_hd__xnor2_1 _20375_ (.A(net283),
    .B(_12127_),
    .Y(_12224_));
 sky130_fd_sc_hd__nor3_1 _20376_ (.A(net276),
    .B(_12127_),
    .C(_12131_),
    .Y(_12225_));
 sky130_fd_sc_hd__a31oi_2 _20377_ (.A1(net276),
    .A2(_12131_),
    .A3(_12224_),
    .B1(_12225_),
    .Y(_12226_));
 sky130_fd_sc_hd__and2_1 _20378_ (.A(_12223_),
    .B(_12226_),
    .X(_12227_));
 sky130_fd_sc_hd__a21o_1 _20379_ (.A1(_12218_),
    .A2(_12219_),
    .B1(_12227_),
    .X(_12228_));
 sky130_fd_sc_hd__nand3_1 _20380_ (.A(_12227_),
    .B(_12218_),
    .C(_12219_),
    .Y(_12229_));
 sky130_fd_sc_hd__and2_1 _20381_ (.A(_12228_),
    .B(_12229_),
    .X(_12230_));
 sky130_fd_sc_hd__and3b_1 _20382_ (.A_N(_12133_),
    .B(_12148_),
    .C(_12149_),
    .X(_12231_));
 sky130_fd_sc_hd__a21bo_1 _20383_ (.A1(_12148_),
    .A2(_12149_),
    .B1_N(_12133_),
    .X(_12232_));
 sky130_fd_sc_hd__o21a_1 _20384_ (.A1(_12125_),
    .A2(_12231_),
    .B1(_12232_),
    .X(_12233_));
 sky130_fd_sc_hd__nand2_1 _20385_ (.A(_12139_),
    .B(_12141_),
    .Y(_12234_));
 sky130_fd_sc_hd__o21a_1 _20386_ (.A1(_12137_),
    .A2(_12234_),
    .B1(_12145_),
    .X(_12235_));
 sky130_fd_sc_hd__a21o_1 _20387_ (.A1(_12137_),
    .A2(_12234_),
    .B1(_12235_),
    .X(_12236_));
 sky130_fd_sc_hd__nand2_1 _20388_ (.A(net214),
    .B(_12165_),
    .Y(_12237_));
 sky130_fd_sc_hd__nand2_2 _20389_ (.A(net235),
    .B(net226),
    .Y(_12238_));
 sky130_fd_sc_hd__xor2_1 _20390_ (.A(_12237_),
    .B(_12238_),
    .X(_12239_));
 sky130_fd_sc_hd__xnor2_2 _20391_ (.A(_12236_),
    .B(_12239_),
    .Y(_12240_));
 sky130_fd_sc_hd__xor2_1 _20392_ (.A(_12233_),
    .B(_12240_),
    .X(_12241_));
 sky130_fd_sc_hd__xnor2_2 _20393_ (.A(_12230_),
    .B(_12241_),
    .Y(_12242_));
 sky130_fd_sc_hd__xnor2_1 _20394_ (.A(_12196_),
    .B(_12242_),
    .Y(_12243_));
 sky130_fd_sc_hd__o21ai_1 _20395_ (.A1(_12172_),
    .A2(_12173_),
    .B1(_12243_),
    .Y(_12244_));
 sky130_fd_sc_hd__and3_1 _20396_ (.A(net264),
    .B(net253),
    .C(net240),
    .X(_12245_));
 sky130_fd_sc_hd__nand2_1 _20397_ (.A(net262),
    .B(net252),
    .Y(_12246_));
 sky130_fd_sc_hd__xnor2_2 _20398_ (.A(_11727_),
    .B(_12246_),
    .Y(_12247_));
 sky130_fd_sc_hd__inv_2 _20399_ (.A(_12247_),
    .Y(_12248_));
 sky130_fd_sc_hd__nor2_1 _20400_ (.A(net289),
    .B(_12047_),
    .Y(_12249_));
 sky130_fd_sc_hd__xnor2_2 _20401_ (.A(net261),
    .B(net249),
    .Y(_12250_));
 sky130_fd_sc_hd__xnor2_2 _20402_ (.A(_12067_),
    .B(_12250_),
    .Y(_12251_));
 sky130_fd_sc_hd__and2b_1 _20403_ (.A_N(_12249_),
    .B(_12251_),
    .X(_12252_));
 sky130_fd_sc_hd__xor2_2 _20404_ (.A(net265),
    .B(net254),
    .X(_12253_));
 sky130_fd_sc_hd__inv_2 _20405_ (.A(_12253_),
    .Y(_12254_));
 sky130_fd_sc_hd__nand2_1 _20406_ (.A(net277),
    .B(net271),
    .Y(_12255_));
 sky130_fd_sc_hd__nand2_1 _20407_ (.A(_12253_),
    .B(_12255_),
    .Y(_12256_));
 sky130_fd_sc_hd__a221o_2 _20408_ (.A1(net269),
    .A2(_12254_),
    .B1(_12256_),
    .B2(_11571_),
    .C1(_12050_),
    .X(_12257_));
 sky130_fd_sc_hd__o31a_1 _20409_ (.A1(net289),
    .A2(_12047_),
    .A3(_12251_),
    .B1(_12257_),
    .X(_12258_));
 sky130_fd_sc_hd__nor2_1 _20410_ (.A(_12252_),
    .B(_12258_),
    .Y(_12259_));
 sky130_fd_sc_hd__a21o_1 _20411_ (.A1(_12245_),
    .A2(_12248_),
    .B1(_12259_),
    .X(_12260_));
 sky130_fd_sc_hd__o21a_1 _20412_ (.A1(_12245_),
    .A2(_12248_),
    .B1(_12260_),
    .X(_12261_));
 sky130_fd_sc_hd__xnor2_4 _20413_ (.A(net275),
    .B(_12108_),
    .Y(_12262_));
 sky130_fd_sc_hd__xnor2_1 _20414_ (.A(net302),
    .B(_12262_),
    .Y(_12263_));
 sky130_fd_sc_hd__nor2b_2 _20415_ (.A(net295),
    .B_N(net298),
    .Y(_12264_));
 sky130_fd_sc_hd__or2b_1 _20416_ (.A(net298),
    .B_N(net294),
    .X(_12265_));
 sky130_fd_sc_hd__o2bb2a_4 _20417_ (.A1_N(_12263_),
    .A2_N(_12264_),
    .B1(_12265_),
    .B2(_12262_),
    .X(_12266_));
 sky130_fd_sc_hd__xor2_2 _20418_ (.A(net256),
    .B(net245),
    .X(_12267_));
 sky130_fd_sc_hd__o21bai_1 _20419_ (.A1(_11653_),
    .A2(_12267_),
    .B1_N(_12144_),
    .Y(_12268_));
 sky130_fd_sc_hd__nand2_2 _20420_ (.A(net267),
    .B(net262),
    .Y(_12269_));
 sky130_fd_sc_hd__a21oi_1 _20421_ (.A1(_12267_),
    .A2(_12269_),
    .B1(net269),
    .Y(_12270_));
 sky130_fd_sc_hd__or2_1 _20422_ (.A(_12268_),
    .B(_12270_),
    .X(_12271_));
 sky130_fd_sc_hd__nand2_1 _20423_ (.A(net304),
    .B(net299),
    .Y(_12272_));
 sky130_fd_sc_hd__or2b_1 _20424_ (.A(net275),
    .B_N(net289),
    .X(_12273_));
 sky130_fd_sc_hd__nor2_1 _20425_ (.A(net281),
    .B(net274),
    .Y(_12274_));
 sky130_fd_sc_hd__a221o_2 _20426_ (.A1(net276),
    .A2(_12108_),
    .B1(_12272_),
    .B2(_12273_),
    .C1(_12274_),
    .X(_12275_));
 sky130_fd_sc_hd__xnor2_2 _20427_ (.A(_12271_),
    .B(_12275_),
    .Y(_12276_));
 sky130_fd_sc_hd__nor2b_2 _20428_ (.A(net300),
    .B_N(net297),
    .Y(_12277_));
 sky130_fd_sc_hd__xnor2_4 _20429_ (.A(net291),
    .B(_12277_),
    .Y(_12278_));
 sky130_fd_sc_hd__xnor2_4 _20430_ (.A(_12056_),
    .B(_12278_),
    .Y(_12279_));
 sky130_fd_sc_hd__xnor2_4 _20431_ (.A(_12042_),
    .B(_12127_),
    .Y(_12280_));
 sky130_fd_sc_hd__xnor2_1 _20432_ (.A(_12279_),
    .B(_12280_),
    .Y(_12281_));
 sky130_fd_sc_hd__xnor2_2 _20433_ (.A(_12276_),
    .B(_12281_),
    .Y(_12282_));
 sky130_fd_sc_hd__xor2_4 _20434_ (.A(_12266_),
    .B(_12282_),
    .X(_12283_));
 sky130_fd_sc_hd__nor2_2 _20435_ (.A(net302),
    .B(_11437_),
    .Y(_12284_));
 sky130_fd_sc_hd__nor2_1 _20436_ (.A(_11407_),
    .B(net299),
    .Y(_12285_));
 sky130_fd_sc_hd__mux2_1 _20437_ (.A0(_12284_),
    .A1(_12285_),
    .S(net274),
    .X(_12286_));
 sky130_fd_sc_hd__and2b_2 _20438_ (.A_N(net294),
    .B(net287),
    .X(_12287_));
 sky130_fd_sc_hd__a22o_1 _20439_ (.A1(_11571_),
    .A2(_12287_),
    .B1(_12108_),
    .B2(net296),
    .X(_12288_));
 sky130_fd_sc_hd__or3_1 _20440_ (.A(_11407_),
    .B(net301),
    .C(net275),
    .X(_12289_));
 sky130_fd_sc_hd__a21bo_1 _20441_ (.A1(net275),
    .A2(_12284_),
    .B1_N(_12289_),
    .X(_12290_));
 sky130_fd_sc_hd__and4b_1 _20442_ (.A_N(_12059_),
    .B(net281),
    .C(_12057_),
    .D(_12290_),
    .X(_12291_));
 sky130_fd_sc_hd__a21oi_1 _20443_ (.A1(_12286_),
    .A2(_12288_),
    .B1(_12291_),
    .Y(_12292_));
 sky130_fd_sc_hd__nand2_1 _20444_ (.A(net271),
    .B(net265),
    .Y(_12293_));
 sky130_fd_sc_hd__or2b_1 _20445_ (.A(_12250_),
    .B_N(_12293_),
    .X(_12294_));
 sky130_fd_sc_hd__a221o_1 _20446_ (.A1(net264),
    .A2(_12250_),
    .B1(_12294_),
    .B2(_11593_),
    .C1(_12090_),
    .X(_12295_));
 sky130_fd_sc_hd__xnor2_2 _20447_ (.A(_12102_),
    .B(_12267_),
    .Y(_12296_));
 sky130_fd_sc_hd__nor2_1 _20448_ (.A(net283),
    .B(_12065_),
    .Y(_12297_));
 sky130_fd_sc_hd__xnor2_1 _20449_ (.A(_12296_),
    .B(_12297_),
    .Y(_12298_));
 sky130_fd_sc_hd__xnor2_2 _20450_ (.A(_12295_),
    .B(_12298_),
    .Y(_12299_));
 sky130_fd_sc_hd__mux2_1 _20451_ (.A0(net302),
    .A1(_12284_),
    .S(net275),
    .X(_12300_));
 sky130_fd_sc_hd__or2b_1 _20452_ (.A(net274),
    .B_N(net294),
    .X(_12301_));
 sky130_fd_sc_hd__or2b_1 _20453_ (.A(net294),
    .B_N(net274),
    .X(_12302_));
 sky130_fd_sc_hd__nand2_1 _20454_ (.A(_12301_),
    .B(_12302_),
    .Y(_12303_));
 sky130_fd_sc_hd__mux2_1 _20455_ (.A0(net287),
    .A1(_12108_),
    .S(_12303_),
    .X(_12304_));
 sky130_fd_sc_hd__nor2_1 _20456_ (.A(_12284_),
    .B(_12285_),
    .Y(_12305_));
 sky130_fd_sc_hd__a32o_1 _20457_ (.A1(net280),
    .A2(_12287_),
    .A3(_12300_),
    .B1(_12304_),
    .B2(_12305_),
    .X(_12306_));
 sky130_fd_sc_hd__or2_1 _20458_ (.A(net287),
    .B(_12302_),
    .X(_12307_));
 sky130_fd_sc_hd__or2_1 _20459_ (.A(net295),
    .B(net275),
    .X(_12308_));
 sky130_fd_sc_hd__nand2_1 _20460_ (.A(net295),
    .B(net278),
    .Y(_12309_));
 sky130_fd_sc_hd__o211a_1 _20461_ (.A1(net288),
    .A2(_12308_),
    .B1(_12309_),
    .C1(net303),
    .X(_12310_));
 sky130_fd_sc_hd__a31o_1 _20462_ (.A1(_11527_),
    .A2(_12308_),
    .A3(_12309_),
    .B1(_12310_),
    .X(_12311_));
 sky130_fd_sc_hd__a311o_1 _20463_ (.A1(_12284_),
    .A2(_12301_),
    .A3(_12307_),
    .B1(_12311_),
    .C1(net280),
    .X(_12312_));
 sky130_fd_sc_hd__or2b_1 _20464_ (.A(_12306_),
    .B_N(_12312_),
    .X(_12313_));
 sky130_fd_sc_hd__a21oi_2 _20465_ (.A1(_12292_),
    .A2(_12299_),
    .B1(_12313_),
    .Y(_12314_));
 sky130_fd_sc_hd__o21ba_1 _20466_ (.A1(_12296_),
    .A2(_12297_),
    .B1_N(_12295_),
    .X(_12315_));
 sky130_fd_sc_hd__a21o_1 _20467_ (.A1(_12296_),
    .A2(_12297_),
    .B1(_12315_),
    .X(_12316_));
 sky130_fd_sc_hd__nand2_1 _20468_ (.A(net257),
    .B(net248),
    .Y(_12317_));
 sky130_fd_sc_hd__xnor2_1 _20469_ (.A(_11739_),
    .B(_12317_),
    .Y(_12318_));
 sky130_fd_sc_hd__nor3_1 _20470_ (.A(_11726_),
    .B(_12246_),
    .C(_12318_),
    .Y(_12319_));
 sky130_fd_sc_hd__o21ai_1 _20471_ (.A1(_11726_),
    .A2(_12246_),
    .B1(_12318_),
    .Y(_12320_));
 sky130_fd_sc_hd__or2b_1 _20472_ (.A(_12319_),
    .B_N(_12320_),
    .X(_12321_));
 sky130_fd_sc_hd__xnor2_2 _20473_ (.A(_12316_),
    .B(_12321_),
    .Y(_12322_));
 sky130_fd_sc_hd__xnor2_2 _20474_ (.A(_12314_),
    .B(_12322_),
    .Y(_12323_));
 sky130_fd_sc_hd__xnor2_4 _20475_ (.A(_12283_),
    .B(_12323_),
    .Y(_12324_));
 sky130_fd_sc_hd__nand2_1 _20476_ (.A(_12261_),
    .B(_12324_),
    .Y(_12325_));
 sky130_fd_sc_hd__nor2_1 _20477_ (.A(net298),
    .B(net282),
    .Y(_12326_));
 sky130_fd_sc_hd__xnor2_1 _20478_ (.A(net300),
    .B(net297),
    .Y(_12327_));
 sky130_fd_sc_hd__mux2_1 _20479_ (.A0(_12264_),
    .A1(_12327_),
    .S(net280),
    .X(_12328_));
 sky130_fd_sc_hd__a22o_1 _20480_ (.A1(_12059_),
    .A2(_12326_),
    .B1(_12328_),
    .B2(net287),
    .X(_12329_));
 sky130_fd_sc_hd__nand2_1 _20481_ (.A(net304),
    .B(_12329_),
    .Y(_12330_));
 sky130_fd_sc_hd__xor2_1 _20482_ (.A(_12251_),
    .B(_12249_),
    .X(_12331_));
 sky130_fd_sc_hd__xnor2_2 _20483_ (.A(_12257_),
    .B(_12331_),
    .Y(_12332_));
 sky130_fd_sc_hd__and3b_1 _20484_ (.A_N(_12059_),
    .B(net302),
    .C(_12057_),
    .X(_12333_));
 sky130_fd_sc_hd__nor2_1 _20485_ (.A(net304),
    .B(_12057_),
    .Y(_12334_));
 sky130_fd_sc_hd__o21ai_1 _20486_ (.A1(_12333_),
    .A2(_12334_),
    .B1(net280),
    .Y(_12335_));
 sky130_fd_sc_hd__or3_1 _20487_ (.A(net304),
    .B(net281),
    .C(_12287_),
    .X(_12336_));
 sky130_fd_sc_hd__nand2_2 _20488_ (.A(net294),
    .B(net280),
    .Y(_12337_));
 sky130_fd_sc_hd__o21a_1 _20489_ (.A1(net280),
    .A2(_12057_),
    .B1(_12337_),
    .X(_12338_));
 sky130_fd_sc_hd__o221a_1 _20490_ (.A1(net289),
    .A2(_12061_),
    .B1(_12338_),
    .B2(net304),
    .C1(net301),
    .X(_12339_));
 sky130_fd_sc_hd__a31oi_2 _20491_ (.A1(_11438_),
    .A2(_12335_),
    .A3(_12336_),
    .B1(_12339_),
    .Y(_12340_));
 sky130_fd_sc_hd__a21oi_1 _20492_ (.A1(_12330_),
    .A2(_12332_),
    .B1(_12340_),
    .Y(_12341_));
 sky130_fd_sc_hd__xor2_2 _20493_ (.A(_12245_),
    .B(_12247_),
    .X(_12342_));
 sky130_fd_sc_hd__xnor2_1 _20494_ (.A(_12259_),
    .B(_12342_),
    .Y(_12343_));
 sky130_fd_sc_hd__and2b_1 _20495_ (.A_N(net282),
    .B(net288),
    .X(_12344_));
 sky130_fd_sc_hd__or3_1 _20496_ (.A(_11437_),
    .B(_12059_),
    .C(_12344_),
    .X(_12345_));
 sky130_fd_sc_hd__o221a_1 _20497_ (.A1(net298),
    .A2(_12065_),
    .B1(_12156_),
    .B2(net295),
    .C1(_12345_),
    .X(_12346_));
 sky130_fd_sc_hd__or2_2 _20498_ (.A(net295),
    .B(net287),
    .X(_12347_));
 sky130_fd_sc_hd__and2b_1 _20499_ (.A_N(net282),
    .B(net295),
    .X(_12348_));
 sky130_fd_sc_hd__a31o_1 _20500_ (.A1(_11438_),
    .A2(_12142_),
    .A3(_12347_),
    .B1(_12348_),
    .X(_12349_));
 sky130_fd_sc_hd__nand2_1 _20501_ (.A(net302),
    .B(_12349_),
    .Y(_12350_));
 sky130_fd_sc_hd__o22a_1 _20502_ (.A1(_11407_),
    .A2(_12065_),
    .B1(_12156_),
    .B2(net296),
    .X(_12351_));
 sky130_fd_sc_hd__o2bb2a_1 _20503_ (.A1_N(net294),
    .A2_N(_12326_),
    .B1(_12351_),
    .B2(_11438_),
    .X(_12352_));
 sky130_fd_sc_hd__o211a_1 _20504_ (.A1(net303),
    .A2(_12346_),
    .B1(_12350_),
    .C1(_12352_),
    .X(_12353_));
 sky130_fd_sc_hd__xnor2_1 _20505_ (.A(net274),
    .B(_12353_),
    .Y(_12354_));
 sky130_fd_sc_hd__xnor2_1 _20506_ (.A(_12299_),
    .B(_12354_),
    .Y(_12355_));
 sky130_fd_sc_hd__o21a_1 _20507_ (.A1(_12341_),
    .A2(_12343_),
    .B1(_12355_),
    .X(_12356_));
 sky130_fd_sc_hd__a21oi_2 _20508_ (.A1(_12341_),
    .A2(_12343_),
    .B1(_12356_),
    .Y(_12357_));
 sky130_fd_sc_hd__nor2_1 _20509_ (.A(_12261_),
    .B(_12324_),
    .Y(_12358_));
 sky130_fd_sc_hd__a21o_1 _20510_ (.A1(_12325_),
    .A2(_12357_),
    .B1(_12358_),
    .X(_12359_));
 sky130_fd_sc_hd__or3_2 _20511_ (.A(_12268_),
    .B(_12270_),
    .C(_12275_),
    .X(_12360_));
 sky130_fd_sc_hd__o21a_1 _20512_ (.A1(_12268_),
    .A2(_12270_),
    .B1(_12275_),
    .X(_12361_));
 sky130_fd_sc_hd__a21o_1 _20513_ (.A1(_12280_),
    .A2(_12360_),
    .B1(_12361_),
    .X(_12362_));
 sky130_fd_sc_hd__or2_1 _20514_ (.A(_12280_),
    .B(_12360_),
    .X(_12363_));
 sky130_fd_sc_hd__o21a_1 _20515_ (.A1(_12266_),
    .A2(_12362_),
    .B1(_12363_),
    .X(_12364_));
 sky130_fd_sc_hd__nand2_1 _20516_ (.A(_12280_),
    .B(_12361_),
    .Y(_12365_));
 sky130_fd_sc_hd__a21bo_1 _20517_ (.A1(_12266_),
    .A2(_12362_),
    .B1_N(_12365_),
    .X(_12366_));
 sky130_fd_sc_hd__nand2_1 _20518_ (.A(_12279_),
    .B(_12366_),
    .Y(_12367_));
 sky130_fd_sc_hd__mux2_1 _20519_ (.A0(_12363_),
    .A1(_12365_),
    .S(_12266_),
    .X(_12368_));
 sky130_fd_sc_hd__o211a_1 _20520_ (.A1(_12279_),
    .A2(_12364_),
    .B1(_12367_),
    .C1(_12368_),
    .X(_12369_));
 sky130_fd_sc_hd__nor2_2 _20521_ (.A(_11739_),
    .B(_12317_),
    .Y(_12370_));
 sky130_fd_sc_hd__xnor2_4 _20522_ (.A(_11758_),
    .B(_12075_),
    .Y(_12371_));
 sky130_fd_sc_hd__xor2_4 _20523_ (.A(_12370_),
    .B(_12371_),
    .X(_12372_));
 sky130_fd_sc_hd__nand2_1 _20524_ (.A(_12054_),
    .B(_12055_),
    .Y(_12373_));
 sky130_fd_sc_hd__xor2_1 _20525_ (.A(_12069_),
    .B(_12060_),
    .X(_12374_));
 sky130_fd_sc_hd__xnor2_1 _20526_ (.A(_12373_),
    .B(_12374_),
    .Y(_12375_));
 sky130_fd_sc_hd__xnor2_1 _20527_ (.A(_12372_),
    .B(_12375_),
    .Y(_12376_));
 sky130_fd_sc_hd__xnor2_2 _20528_ (.A(_12369_),
    .B(_12376_),
    .Y(_12377_));
 sky130_fd_sc_hd__a21o_1 _20529_ (.A1(_12283_),
    .A2(_12314_),
    .B1(_12322_),
    .X(_12378_));
 sky130_fd_sc_hd__or2_1 _20530_ (.A(_12283_),
    .B(_12314_),
    .X(_12379_));
 sky130_fd_sc_hd__a21o_1 _20531_ (.A1(_12316_),
    .A2(_12320_),
    .B1(_12319_),
    .X(_12380_));
 sky130_fd_sc_hd__a21oi_1 _20532_ (.A1(_12378_),
    .A2(_12379_),
    .B1(_12380_),
    .Y(_12381_));
 sky130_fd_sc_hd__and3_1 _20533_ (.A(_12378_),
    .B(_12379_),
    .C(_12380_),
    .X(_12382_));
 sky130_fd_sc_hd__or2_1 _20534_ (.A(_12381_),
    .B(_12382_),
    .X(_12383_));
 sky130_fd_sc_hd__xnor2_2 _20535_ (.A(_12377_),
    .B(_12383_),
    .Y(_12384_));
 sky130_fd_sc_hd__nand2_1 _20536_ (.A(_12359_),
    .B(_12384_),
    .Y(_12385_));
 sky130_fd_sc_hd__nor2_1 _20537_ (.A(_12279_),
    .B(_12266_),
    .Y(_12386_));
 sky130_fd_sc_hd__a21oi_1 _20538_ (.A1(_12280_),
    .A2(_12360_),
    .B1(_12361_),
    .Y(_12387_));
 sky130_fd_sc_hd__mux2_1 _20539_ (.A0(_12361_),
    .A1(_12387_),
    .S(_12372_),
    .X(_12388_));
 sky130_fd_sc_hd__or2_1 _20540_ (.A(_12372_),
    .B(_12276_),
    .X(_12389_));
 sky130_fd_sc_hd__nand2_1 _20541_ (.A(_12271_),
    .B(_12275_),
    .Y(_12390_));
 sky130_fd_sc_hd__mux2_1 _20542_ (.A0(_12360_),
    .A1(_12390_),
    .S(_12372_),
    .X(_12391_));
 sky130_fd_sc_hd__mux2_1 _20543_ (.A0(_12389_),
    .A1(_12391_),
    .S(_12280_),
    .X(_12392_));
 sky130_fd_sc_hd__mux2_1 _20544_ (.A0(_12360_),
    .A1(_12387_),
    .S(_12372_),
    .X(_12393_));
 sky130_fd_sc_hd__nand2_1 _20545_ (.A(_12279_),
    .B(_12266_),
    .Y(_12394_));
 sky130_fd_sc_hd__o221a_1 _20546_ (.A1(_12386_),
    .A2(_12392_),
    .B1(_12393_),
    .B2(_12394_),
    .C1(_12375_),
    .X(_12395_));
 sky130_fd_sc_hd__mux2_1 _20547_ (.A0(_12390_),
    .A1(_12276_),
    .S(_12280_),
    .X(_12396_));
 sky130_fd_sc_hd__mux2_1 _20548_ (.A0(_12396_),
    .A1(_12363_),
    .S(_12372_),
    .X(_12397_));
 sky130_fd_sc_hd__a21oi_1 _20549_ (.A1(_12279_),
    .A2(_12266_),
    .B1(_12397_),
    .Y(_12398_));
 sky130_fd_sc_hd__a211oi_2 _20550_ (.A1(_12386_),
    .A2(_12388_),
    .B1(_12395_),
    .C1(_12398_),
    .Y(_12399_));
 sky130_fd_sc_hd__o21ba_1 _20551_ (.A1(_12377_),
    .A2(_12381_),
    .B1_N(_12382_),
    .X(_12400_));
 sky130_fd_sc_hd__and2_1 _20552_ (.A(_12399_),
    .B(_12400_),
    .X(_12401_));
 sky130_fd_sc_hd__nor2_1 _20553_ (.A(_12399_),
    .B(_12400_),
    .Y(_12402_));
 sky130_fd_sc_hd__or3b_1 _20554_ (.A(_12116_),
    .B(_12171_),
    .C_N(_12084_),
    .X(_12403_));
 sky130_fd_sc_hd__a21o_1 _20555_ (.A1(_12077_),
    .A2(_12082_),
    .B1(_12076_),
    .X(_12404_));
 sky130_fd_sc_hd__nand4_1 _20556_ (.A(_12083_),
    .B(_12070_),
    .C(_12071_),
    .D(_12171_),
    .Y(_12405_));
 sky130_fd_sc_hd__o41a_1 _20557_ (.A1(_12113_),
    .A2(_12114_),
    .A3(_12084_),
    .A4(_12404_),
    .B1(_12405_),
    .X(_12406_));
 sky130_fd_sc_hd__o311a_1 _20558_ (.A1(_12115_),
    .A2(_12116_),
    .A3(_12171_),
    .B1(_12403_),
    .C1(_12406_),
    .X(_12407_));
 sky130_fd_sc_hd__xnor2_2 _20559_ (.A(_12170_),
    .B(_12407_),
    .Y(_12408_));
 sky130_fd_sc_hd__mux2_1 _20560_ (.A0(_12401_),
    .A1(_12402_),
    .S(_12408_),
    .X(_12409_));
 sky130_fd_sc_hd__or2_1 _20561_ (.A(_12084_),
    .B(_12116_),
    .X(_12410_));
 sky130_fd_sc_hd__xnor2_2 _20562_ (.A(_12115_),
    .B(_12410_),
    .Y(_12411_));
 sky130_fd_sc_hd__inv_2 _20563_ (.A(_12371_),
    .Y(_12412_));
 sky130_fd_sc_hd__a21oi_1 _20564_ (.A1(_12370_),
    .A2(_12412_),
    .B1(_12387_),
    .Y(_12413_));
 sky130_fd_sc_hd__o21ba_1 _20565_ (.A1(_12370_),
    .A2(_12412_),
    .B1_N(_12413_),
    .X(_12414_));
 sky130_fd_sc_hd__xor2_1 _20566_ (.A(_12411_),
    .B(_12414_),
    .X(_12415_));
 sky130_fd_sc_hd__or2_1 _20567_ (.A(_12411_),
    .B(_12414_),
    .X(_12416_));
 sky130_fd_sc_hd__nand2_1 _20568_ (.A(_12411_),
    .B(_12414_),
    .Y(_12417_));
 sky130_fd_sc_hd__mux2_1 _20569_ (.A0(_12416_),
    .A1(_12417_),
    .S(_12408_),
    .X(_12418_));
 sky130_fd_sc_hd__a2111oi_1 _20570_ (.A1(_12359_),
    .A2(_12384_),
    .B1(_12401_),
    .C1(_12402_),
    .D1(_12418_),
    .Y(_12419_));
 sky130_fd_sc_hd__a31o_1 _20571_ (.A1(_12385_),
    .A2(_12409_),
    .A3(_12415_),
    .B1(_12419_),
    .X(_12420_));
 sky130_fd_sc_hd__inv_2 _20572_ (.A(_12340_),
    .Y(_12421_));
 sky130_fd_sc_hd__a21oi_1 _20573_ (.A1(net304),
    .A2(_12329_),
    .B1(_12249_),
    .Y(_12422_));
 sky130_fd_sc_hd__or4_1 _20574_ (.A(_12251_),
    .B(_12257_),
    .C(_12340_),
    .D(_12422_),
    .X(_12423_));
 sky130_fd_sc_hd__nand3_1 _20575_ (.A(_12251_),
    .B(_12257_),
    .C(_12422_),
    .Y(_12424_));
 sky130_fd_sc_hd__o211a_1 _20576_ (.A1(_12259_),
    .A2(_12421_),
    .B1(_12423_),
    .C1(_12424_),
    .X(_12425_));
 sky130_fd_sc_hd__xnor2_1 _20577_ (.A(_12355_),
    .B(_12425_),
    .Y(_12426_));
 sky130_fd_sc_hd__xnor2_2 _20578_ (.A(_12342_),
    .B(_12426_),
    .Y(_12427_));
 sky130_fd_sc_hd__xnor2_2 _20579_ (.A(_12056_),
    .B(_12254_),
    .Y(_12428_));
 sky130_fd_sc_hd__xnor2_2 _20580_ (.A(net270),
    .B(net258),
    .Y(_12429_));
 sky130_fd_sc_hd__a21o_1 _20581_ (.A1(net275),
    .A2(_12429_),
    .B1(_12274_),
    .X(_12430_));
 sky130_fd_sc_hd__o21a_1 _20582_ (.A1(_12201_),
    .A2(_12429_),
    .B1(_11550_),
    .X(_12431_));
 sky130_fd_sc_hd__nand2_1 _20583_ (.A(net302),
    .B(_12264_),
    .Y(_12432_));
 sky130_fd_sc_hd__or3_1 _20584_ (.A(_12430_),
    .B(_12431_),
    .C(_12432_),
    .X(_12433_));
 sky130_fd_sc_hd__o21a_1 _20585_ (.A1(_12430_),
    .A2(_12431_),
    .B1(_12432_),
    .X(_12434_));
 sky130_fd_sc_hd__a21oi_1 _20586_ (.A1(_12428_),
    .A2(_12433_),
    .B1(_12434_),
    .Y(_12435_));
 sky130_fd_sc_hd__and3_1 _20587_ (.A(net270),
    .B(net258),
    .C(net245),
    .X(_12436_));
 sky130_fd_sc_hd__nand2_1 _20588_ (.A(net264),
    .B(net253),
    .Y(_12437_));
 sky130_fd_sc_hd__xnor2_2 _20589_ (.A(net240),
    .B(_12437_),
    .Y(_12438_));
 sky130_fd_sc_hd__xor2_1 _20590_ (.A(_12436_),
    .B(_12438_),
    .X(_12439_));
 sky130_fd_sc_hd__xnor2_1 _20591_ (.A(_12435_),
    .B(_12439_),
    .Y(_12440_));
 sky130_fd_sc_hd__nor2_1 _20592_ (.A(_12059_),
    .B(_12264_),
    .Y(_12441_));
 sky130_fd_sc_hd__nor2_1 _20593_ (.A(net298),
    .B(_12057_),
    .Y(_12442_));
 sky130_fd_sc_hd__a221o_1 _20594_ (.A1(_12057_),
    .A2(_12284_),
    .B1(_12441_),
    .B2(net302),
    .C1(_12442_),
    .X(_12443_));
 sky130_fd_sc_hd__xnor2_1 _20595_ (.A(net281),
    .B(_12443_),
    .Y(_12444_));
 sky130_fd_sc_hd__xnor2_2 _20596_ (.A(_12332_),
    .B(_12444_),
    .Y(_12445_));
 sky130_fd_sc_hd__or2_1 _20597_ (.A(_12440_),
    .B(_12445_),
    .X(_12446_));
 sky130_fd_sc_hd__or2_1 _20598_ (.A(_12272_),
    .B(_12347_),
    .X(_12447_));
 sky130_fd_sc_hd__a21oi_1 _20599_ (.A1(_11408_),
    .A2(_12059_),
    .B1(_12333_),
    .Y(_12448_));
 sky130_fd_sc_hd__mux2_1 _20600_ (.A0(net287),
    .A1(_12059_),
    .S(net302),
    .X(_12449_));
 sky130_fd_sc_hd__nand2_1 _20601_ (.A(net298),
    .B(_12449_),
    .Y(_12450_));
 sky130_fd_sc_hd__o221a_1 _20602_ (.A1(net302),
    .A2(_12057_),
    .B1(_12448_),
    .B2(net298),
    .C1(_12450_),
    .X(_12451_));
 sky130_fd_sc_hd__nor2_1 _20603_ (.A(_12430_),
    .B(_12431_),
    .Y(_12452_));
 sky130_fd_sc_hd__xnor2_2 _20604_ (.A(_12428_),
    .B(_12452_),
    .Y(_12453_));
 sky130_fd_sc_hd__mux2_1 _20605_ (.A0(_12447_),
    .A1(_12451_),
    .S(_12453_),
    .X(_12454_));
 sky130_fd_sc_hd__a21o_1 _20606_ (.A1(_12440_),
    .A2(_12445_),
    .B1(_12454_),
    .X(_12455_));
 sky130_fd_sc_hd__a21o_1 _20607_ (.A1(_12436_),
    .A2(_12438_),
    .B1(_12435_),
    .X(_12456_));
 sky130_fd_sc_hd__o21ai_2 _20608_ (.A1(_12436_),
    .A2(_12438_),
    .B1(_12456_),
    .Y(_12457_));
 sky130_fd_sc_hd__a21o_1 _20609_ (.A1(_12446_),
    .A2(_12455_),
    .B1(_12457_),
    .X(_12458_));
 sky130_fd_sc_hd__nand3_1 _20610_ (.A(_12457_),
    .B(_12446_),
    .C(_12455_),
    .Y(_12459_));
 sky130_fd_sc_hd__nand3_2 _20611_ (.A(_12427_),
    .B(_12458_),
    .C(_12459_),
    .Y(_12460_));
 sky130_fd_sc_hd__a21o_1 _20612_ (.A1(_12458_),
    .A2(_12459_),
    .B1(_12427_),
    .X(_12461_));
 sky130_fd_sc_hd__xor2_1 _20613_ (.A(_12440_),
    .B(_12454_),
    .X(_12462_));
 sky130_fd_sc_hd__xnor2_2 _20614_ (.A(_12445_),
    .B(_12462_),
    .Y(_12463_));
 sky130_fd_sc_hd__and3_1 _20615_ (.A(net274),
    .B(net263),
    .C(net249),
    .X(_12464_));
 sky130_fd_sc_hd__xor2_2 _20616_ (.A(net275),
    .B(net263),
    .X(_12465_));
 sky130_fd_sc_hd__inv_2 _20617_ (.A(_12465_),
    .Y(_12466_));
 sky130_fd_sc_hd__nand2_1 _20618_ (.A(_12142_),
    .B(_12465_),
    .Y(_12467_));
 sky130_fd_sc_hd__nor2_1 _20619_ (.A(net288),
    .B(net282),
    .Y(_12468_));
 sky130_fd_sc_hd__a221o_2 _20620_ (.A1(net282),
    .A2(_12466_),
    .B1(_12467_),
    .B2(_11525_),
    .C1(_12468_),
    .X(_12469_));
 sky130_fd_sc_hd__xnor2_2 _20621_ (.A(_12262_),
    .B(_12429_),
    .Y(_12470_));
 sky130_fd_sc_hd__nor2_2 _20622_ (.A(_12469_),
    .B(_12470_),
    .Y(_12471_));
 sky130_fd_sc_hd__nand2_1 _20623_ (.A(net270),
    .B(net258),
    .Y(_12472_));
 sky130_fd_sc_hd__xor2_1 _20624_ (.A(net245),
    .B(_12472_),
    .X(_12473_));
 sky130_fd_sc_hd__a21bo_1 _20625_ (.A1(_12464_),
    .A2(_12471_),
    .B1_N(_12473_),
    .X(_12474_));
 sky130_fd_sc_hd__o21a_1 _20626_ (.A1(_12464_),
    .A2(_12471_),
    .B1(_12474_),
    .X(_12475_));
 sky130_fd_sc_hd__nand2_1 _20627_ (.A(_12463_),
    .B(_12475_),
    .Y(_12476_));
 sky130_fd_sc_hd__xnor2_1 _20628_ (.A(_12473_),
    .B(_12464_),
    .Y(_12477_));
 sky130_fd_sc_hd__mux2_1 _20629_ (.A0(_12277_),
    .A1(_12327_),
    .S(net306),
    .X(_12478_));
 sky130_fd_sc_hd__xnor2_1 _20630_ (.A(net287),
    .B(_12478_),
    .Y(_12479_));
 sky130_fd_sc_hd__xnor2_2 _20631_ (.A(_12453_),
    .B(_12479_),
    .Y(_12480_));
 sky130_fd_sc_hd__xnor2_1 _20632_ (.A(net294),
    .B(_12284_),
    .Y(_12481_));
 sky130_fd_sc_hd__a21oi_2 _20633_ (.A1(_12469_),
    .A2(_12470_),
    .B1(_12481_),
    .Y(_12482_));
 sky130_fd_sc_hd__or2_1 _20634_ (.A(_12471_),
    .B(_12482_),
    .X(_12483_));
 sky130_fd_sc_hd__a21oi_1 _20635_ (.A1(_12480_),
    .A2(_12483_),
    .B1(_12477_),
    .Y(_12484_));
 sky130_fd_sc_hd__nor2_1 _20636_ (.A(_12480_),
    .B(_12482_),
    .Y(_12485_));
 sky130_fd_sc_hd__a211o_1 _20637_ (.A1(_12471_),
    .A2(_12477_),
    .B1(_12484_),
    .C1(_12485_),
    .X(_12486_));
 sky130_fd_sc_hd__a31o_1 _20638_ (.A1(_12460_),
    .A2(_12461_),
    .A3(_12476_),
    .B1(_12486_),
    .X(_12487_));
 sky130_fd_sc_hd__nor2_1 _20639_ (.A(_12463_),
    .B(_12475_),
    .Y(_12488_));
 sky130_fd_sc_hd__a21o_1 _20640_ (.A1(_12460_),
    .A2(_12461_),
    .B1(_12488_),
    .X(_12489_));
 sky130_fd_sc_hd__xnor2_2 _20641_ (.A(net280),
    .B(_12287_),
    .Y(_12490_));
 sky130_fd_sc_hd__xor2_4 _20642_ (.A(net285),
    .B(net273),
    .X(_12491_));
 sky130_fd_sc_hd__a21o_1 _20643_ (.A1(_12065_),
    .A2(_12491_),
    .B1(net298),
    .X(_12492_));
 sky130_fd_sc_hd__o211a_1 _20644_ (.A1(_11550_),
    .A2(_12491_),
    .B1(_12492_),
    .C1(_12347_),
    .X(_12493_));
 sky130_fd_sc_hd__mux2_1 _20645_ (.A0(net263),
    .A1(_12490_),
    .S(_12493_),
    .X(_12494_));
 sky130_fd_sc_hd__nor2_1 _20646_ (.A(net274),
    .B(net263),
    .Y(_12495_));
 sky130_fd_sc_hd__mux2_1 _20647_ (.A0(_12495_),
    .A1(net263),
    .S(_12490_),
    .X(_12496_));
 sky130_fd_sc_hd__a22o_1 _20648_ (.A1(net274),
    .A2(_12494_),
    .B1(_12496_),
    .B2(_12493_),
    .X(_12497_));
 sky130_fd_sc_hd__and3_1 _20649_ (.A(net280),
    .B(net270),
    .C(net253),
    .X(_12498_));
 sky130_fd_sc_hd__clkbuf_2 _20650_ (.A(_12498_),
    .X(_12499_));
 sky130_fd_sc_hd__xnor2_1 _20651_ (.A(net249),
    .B(_12499_),
    .Y(_12500_));
 sky130_fd_sc_hd__xnor2_2 _20652_ (.A(_12497_),
    .B(_12500_),
    .Y(_12501_));
 sky130_fd_sc_hd__xnor2_1 _20653_ (.A(_12470_),
    .B(_12481_),
    .Y(_12502_));
 sky130_fd_sc_hd__xnor2_2 _20654_ (.A(_12469_),
    .B(_12502_),
    .Y(_12503_));
 sky130_fd_sc_hd__mux2_1 _20655_ (.A0(net270),
    .A1(net280),
    .S(net287),
    .X(_12504_));
 sky130_fd_sc_hd__or2_1 _20656_ (.A(net298),
    .B(_12504_),
    .X(_12505_));
 sky130_fd_sc_hd__or2b_1 _20657_ (.A(net270),
    .B_N(net287),
    .X(_12506_));
 sky130_fd_sc_hd__a21o_1 _20658_ (.A1(_12156_),
    .A2(_12506_),
    .B1(_11438_),
    .X(_12507_));
 sky130_fd_sc_hd__a21oi_1 _20659_ (.A1(_12156_),
    .A2(_12506_),
    .B1(net294),
    .Y(_12508_));
 sky130_fd_sc_hd__a31o_1 _20660_ (.A1(net294),
    .A2(_12505_),
    .A3(_12507_),
    .B1(_12508_),
    .X(_12509_));
 sky130_fd_sc_hd__nor2_1 _20661_ (.A(_12465_),
    .B(_12509_),
    .Y(_12510_));
 sky130_fd_sc_hd__nand2_1 _20662_ (.A(_12465_),
    .B(_12509_),
    .Y(_12511_));
 sky130_fd_sc_hd__or3b_2 _20663_ (.A(_12305_),
    .B(_12510_),
    .C_N(_12511_),
    .X(_12512_));
 sky130_fd_sc_hd__nand2_1 _20664_ (.A(_12503_),
    .B(_12512_),
    .Y(_12513_));
 sky130_fd_sc_hd__nor2_1 _20665_ (.A(_12503_),
    .B(_12512_),
    .Y(_12514_));
 sky130_fd_sc_hd__a21oi_2 _20666_ (.A1(_12501_),
    .A2(_12513_),
    .B1(_12514_),
    .Y(_12515_));
 sky130_fd_sc_hd__inv_2 _20667_ (.A(_12515_),
    .Y(_12516_));
 sky130_fd_sc_hd__or3b_1 _20668_ (.A(_12471_),
    .B(_12482_),
    .C_N(_12477_),
    .X(_12517_));
 sky130_fd_sc_hd__o21bai_1 _20669_ (.A1(_12471_),
    .A2(_12482_),
    .B1_N(_12477_),
    .Y(_12518_));
 sky130_fd_sc_hd__a21bo_1 _20670_ (.A1(_12517_),
    .A2(_12518_),
    .B1_N(_12480_),
    .X(_12519_));
 sky130_fd_sc_hd__nand3b_1 _20671_ (.A_N(_12480_),
    .B(_12517_),
    .C(_12518_),
    .Y(_12520_));
 sky130_fd_sc_hd__o21a_1 _20672_ (.A1(net249),
    .A2(_12499_),
    .B1(_12490_),
    .X(_12521_));
 sky130_fd_sc_hd__o21ba_1 _20673_ (.A1(_11689_),
    .A2(_12499_),
    .B1_N(_12490_),
    .X(_12522_));
 sky130_fd_sc_hd__mux2_1 _20674_ (.A0(_12521_),
    .A1(_12522_),
    .S(net263),
    .X(_12523_));
 sky130_fd_sc_hd__a32o_1 _20675_ (.A1(net263),
    .A2(_11689_),
    .A3(_12499_),
    .B1(_12523_),
    .B2(_12493_),
    .X(_12524_));
 sky130_fd_sc_hd__nand2_1 _20676_ (.A(net249),
    .B(_12499_),
    .Y(_12525_));
 sky130_fd_sc_hd__xnor2_1 _20677_ (.A(net263),
    .B(_12490_),
    .Y(_12526_));
 sky130_fd_sc_hd__o211ai_1 _20678_ (.A1(net249),
    .A2(_12499_),
    .B1(_12526_),
    .C1(_12493_),
    .Y(_12527_));
 sky130_fd_sc_hd__a21oi_1 _20679_ (.A1(_12525_),
    .A2(_12527_),
    .B1(net274),
    .Y(_12528_));
 sky130_fd_sc_hd__nor2_1 _20680_ (.A(net263),
    .B(_12525_),
    .Y(_12529_));
 sky130_fd_sc_hd__a211o_1 _20681_ (.A1(net274),
    .A2(_12524_),
    .B1(_12528_),
    .C1(_12529_),
    .X(_12530_));
 sky130_fd_sc_hd__a21o_1 _20682_ (.A1(_12519_),
    .A2(_12520_),
    .B1(_12530_),
    .X(_12531_));
 sky130_fd_sc_hd__nand3_2 _20683_ (.A(_12530_),
    .B(_12519_),
    .C(_12520_),
    .Y(_12532_));
 sky130_fd_sc_hd__a21boi_1 _20684_ (.A1(_12516_),
    .A2(_12531_),
    .B1_N(_12532_),
    .Y(_12533_));
 sky130_fd_sc_hd__xnor2_2 _20685_ (.A(_12261_),
    .B(_12357_),
    .Y(_12534_));
 sky130_fd_sc_hd__xnor2_4 _20686_ (.A(_12324_),
    .B(_12534_),
    .Y(_12535_));
 sky130_fd_sc_hd__a211o_1 _20687_ (.A1(_12487_),
    .A2(_12489_),
    .B1(_12533_),
    .C1(_12535_),
    .X(_12536_));
 sky130_fd_sc_hd__or2_1 _20688_ (.A(_12427_),
    .B(_12457_),
    .X(_12537_));
 sky130_fd_sc_hd__and2_1 _20689_ (.A(_12427_),
    .B(_12457_),
    .X(_12538_));
 sky130_fd_sc_hd__a31o_1 _20690_ (.A1(_12446_),
    .A2(_12455_),
    .A3(_12537_),
    .B1(_12538_),
    .X(_12539_));
 sky130_fd_sc_hd__a21o_1 _20691_ (.A1(_12476_),
    .A2(_12486_),
    .B1(_12488_),
    .X(_12540_));
 sky130_fd_sc_hd__a21o_1 _20692_ (.A1(_12460_),
    .A2(_12461_),
    .B1(_12540_),
    .X(_12541_));
 sky130_fd_sc_hd__a21o_1 _20693_ (.A1(_12539_),
    .A2(_12541_),
    .B1(_12535_),
    .X(_12542_));
 sky130_fd_sc_hd__o211ai_2 _20694_ (.A1(_12359_),
    .A2(_12384_),
    .B1(_12536_),
    .C1(_12542_),
    .Y(_12543_));
 sky130_fd_sc_hd__a21oi_1 _20695_ (.A1(_12531_),
    .A2(_12532_),
    .B1(_12515_),
    .Y(_12544_));
 sky130_fd_sc_hd__and3_1 _20696_ (.A(_12515_),
    .B(_12531_),
    .C(_12532_),
    .X(_12545_));
 sky130_fd_sc_hd__nor2_2 _20697_ (.A(_12544_),
    .B(_12545_),
    .Y(_12546_));
 sky130_fd_sc_hd__nand2_1 _20698_ (.A(_12347_),
    .B(_12309_),
    .Y(_12547_));
 sky130_fd_sc_hd__xnor2_1 _20699_ (.A(net300),
    .B(_12491_),
    .Y(_12548_));
 sky130_fd_sc_hd__xnor2_1 _20700_ (.A(_12547_),
    .B(_12548_),
    .Y(_12549_));
 sky130_fd_sc_hd__o21ai_1 _20701_ (.A1(net285),
    .A2(net273),
    .B1(_12278_),
    .Y(_12550_));
 sky130_fd_sc_hd__xor2_2 _20702_ (.A(net289),
    .B(net278),
    .X(_12551_));
 sky130_fd_sc_hd__a21o_1 _20703_ (.A1(_12047_),
    .A2(_12551_),
    .B1(net305),
    .X(_12552_));
 sky130_fd_sc_hd__xnor2_4 _20704_ (.A(net292),
    .B(net278),
    .Y(_12553_));
 sky130_fd_sc_hd__nor2_1 _20705_ (.A(net301),
    .B(net296),
    .Y(_12554_));
 sky130_fd_sc_hd__a21oi_1 _20706_ (.A1(net296),
    .A2(_12553_),
    .B1(_12554_),
    .Y(_12555_));
 sky130_fd_sc_hd__nor2_1 _20707_ (.A(net285),
    .B(_11608_),
    .Y(_12556_));
 sky130_fd_sc_hd__a311o_1 _20708_ (.A1(net285),
    .A2(_12552_),
    .A3(_12555_),
    .B1(_12278_),
    .C1(_12556_),
    .X(_12557_));
 sky130_fd_sc_hd__and3_1 _20709_ (.A(net292),
    .B(net278),
    .C(net261),
    .X(_12558_));
 sky130_fd_sc_hd__buf_6 _20710_ (.A(_12558_),
    .X(_12559_));
 sky130_fd_sc_hd__o2bb2a_1 _20711_ (.A1_N(_12552_),
    .A2_N(_12555_),
    .B1(_11571_),
    .B2(_11608_),
    .X(_12560_));
 sky130_fd_sc_hd__a211o_1 _20712_ (.A1(_12550_),
    .A2(_12557_),
    .B1(_12559_),
    .C1(_12560_),
    .X(_12561_));
 sky130_fd_sc_hd__o311a_1 _20713_ (.A1(net285),
    .A2(net273),
    .A3(_12277_),
    .B1(_12552_),
    .C1(_12555_),
    .X(_12562_));
 sky130_fd_sc_hd__o21ai_1 _20714_ (.A1(_12560_),
    .A2(_12562_),
    .B1(_12559_),
    .Y(_12563_));
 sky130_fd_sc_hd__a21oi_1 _20715_ (.A1(_12561_),
    .A2(_12563_),
    .B1(_11673_),
    .Y(_12564_));
 sky130_fd_sc_hd__and3_1 _20716_ (.A(_11673_),
    .B(_12561_),
    .C(_12563_),
    .X(_12565_));
 sky130_fd_sc_hd__or2_1 _20717_ (.A(_12564_),
    .B(_12565_),
    .X(_12566_));
 sky130_fd_sc_hd__nor2_1 _20718_ (.A(_12265_),
    .B(_12504_),
    .Y(_12567_));
 sky130_fd_sc_hd__and3_1 _20719_ (.A(_12156_),
    .B(_12327_),
    .C(_12506_),
    .X(_12568_));
 sky130_fd_sc_hd__a211o_1 _20720_ (.A1(net298),
    .A2(_12508_),
    .B1(_12567_),
    .C1(_12568_),
    .X(_12569_));
 sky130_fd_sc_hd__xnor2_1 _20721_ (.A(_11593_),
    .B(_12569_),
    .Y(_12570_));
 sky130_fd_sc_hd__xnor2_1 _20722_ (.A(net268),
    .B(_12570_),
    .Y(_12571_));
 sky130_fd_sc_hd__and2_1 _20723_ (.A(net306),
    .B(_12549_),
    .X(_12572_));
 sky130_fd_sc_hd__or3_1 _20724_ (.A(_12572_),
    .B(_12564_),
    .C(_12565_),
    .X(_12573_));
 sky130_fd_sc_hd__nor2_1 _20725_ (.A(net306),
    .B(_12571_),
    .Y(_12574_));
 sky130_fd_sc_hd__a221o_2 _20726_ (.A1(_12549_),
    .A2(_12566_),
    .B1(_12571_),
    .B2(_12573_),
    .C1(_12574_),
    .X(_12575_));
 sky130_fd_sc_hd__xnor2_1 _20727_ (.A(_12503_),
    .B(_12512_),
    .Y(_12576_));
 sky130_fd_sc_hd__xnor2_2 _20728_ (.A(_12501_),
    .B(_12576_),
    .Y(_12577_));
 sky130_fd_sc_hd__inv_2 _20729_ (.A(_12577_),
    .Y(_12578_));
 sky130_fd_sc_hd__or2_1 _20730_ (.A(_12575_),
    .B(_12578_),
    .X(_12579_));
 sky130_fd_sc_hd__nand2_1 _20731_ (.A(_12561_),
    .B(_12563_),
    .Y(_12580_));
 sky130_fd_sc_hd__xnor2_1 _20732_ (.A(_12253_),
    .B(_12572_),
    .Y(_12581_));
 sky130_fd_sc_hd__xnor2_1 _20733_ (.A(_12570_),
    .B(_12581_),
    .Y(_12582_));
 sky130_fd_sc_hd__xnor2_2 _20734_ (.A(_12580_),
    .B(_12582_),
    .Y(_12583_));
 sky130_fd_sc_hd__and2b_1 _20735_ (.A_N(net295),
    .B(net282),
    .X(_12584_));
 sky130_fd_sc_hd__mux2_1 _20736_ (.A0(_12348_),
    .A1(_12584_),
    .S(_12553_),
    .X(_12585_));
 sky130_fd_sc_hd__mux2_1 _20737_ (.A0(_12348_),
    .A1(_12584_),
    .S(_12551_),
    .X(_12586_));
 sky130_fd_sc_hd__a22o_1 _20738_ (.A1(_12284_),
    .A2(_12585_),
    .B1(_12586_),
    .B2(_12285_),
    .X(_12587_));
 sky130_fd_sc_hd__and3_1 _20739_ (.A(net294),
    .B(net282),
    .C(net264),
    .X(_12588_));
 sky130_fd_sc_hd__or2_1 _20740_ (.A(_12587_),
    .B(_12588_),
    .X(_12589_));
 sky130_fd_sc_hd__or3_1 _20741_ (.A(net301),
    .B(_11525_),
    .C(_12551_),
    .X(_12590_));
 sky130_fd_sc_hd__a21o_1 _20742_ (.A1(net295),
    .A2(_12553_),
    .B1(_11437_),
    .X(_12591_));
 sky130_fd_sc_hd__nand2_1 _20743_ (.A(net305),
    .B(_12491_),
    .Y(_12592_));
 sky130_fd_sc_hd__a21oi_1 _20744_ (.A1(_12590_),
    .A2(_12591_),
    .B1(_12592_),
    .Y(_12593_));
 sky130_fd_sc_hd__and4bb_1 _20745_ (.A_N(_11407_),
    .B_N(_12491_),
    .C(_12590_),
    .D(_12591_),
    .X(_12594_));
 sky130_fd_sc_hd__nand2_1 _20746_ (.A(_12264_),
    .B(_12551_),
    .Y(_12595_));
 sky130_fd_sc_hd__a211oi_1 _20747_ (.A1(_12590_),
    .A2(_12595_),
    .B1(net303),
    .C1(_12491_),
    .Y(_12596_));
 sky130_fd_sc_hd__and4_1 _20748_ (.A(_11408_),
    .B(_12491_),
    .C(_12590_),
    .D(_12595_),
    .X(_12597_));
 sky130_fd_sc_hd__or4_4 _20749_ (.A(_12593_),
    .B(_12594_),
    .C(_12596_),
    .D(_12597_),
    .X(_12598_));
 sky130_fd_sc_hd__o21a_1 _20750_ (.A1(_12589_),
    .A2(_12598_),
    .B1(net258),
    .X(_12599_));
 sky130_fd_sc_hd__a211o_1 _20751_ (.A1(_12589_),
    .A2(_12598_),
    .B1(_12599_),
    .C1(net288),
    .X(_12600_));
 sky130_fd_sc_hd__a21oi_1 _20752_ (.A1(_11593_),
    .A2(net258),
    .B1(_12589_),
    .Y(_12601_));
 sky130_fd_sc_hd__nor2_1 _20753_ (.A(_12587_),
    .B(_12588_),
    .Y(_12602_));
 sky130_fd_sc_hd__a211o_1 _20754_ (.A1(_12602_),
    .A2(_12598_),
    .B1(_11593_),
    .C1(net258),
    .X(_12603_));
 sky130_fd_sc_hd__o211ai_1 _20755_ (.A1(_12598_),
    .A2(_12601_),
    .B1(_12603_),
    .C1(net287),
    .Y(_12604_));
 sky130_fd_sc_hd__a32o_1 _20756_ (.A1(_11593_),
    .A2(net258),
    .A3(_12589_),
    .B1(_12600_),
    .B2(_12604_),
    .X(_12605_));
 sky130_fd_sc_hd__nor2_1 _20757_ (.A(_12583_),
    .B(_12605_),
    .Y(_12606_));
 sky130_fd_sc_hd__a211o_1 _20758_ (.A1(net300),
    .A2(net285),
    .B1(_12554_),
    .C1(net302),
    .X(_12607_));
 sky130_fd_sc_hd__o31a_2 _20759_ (.A1(_11408_),
    .A2(_12264_),
    .A3(_12326_),
    .B1(_12607_),
    .X(_12608_));
 sky130_fd_sc_hd__xnor2_4 _20760_ (.A(_12553_),
    .B(_12608_),
    .Y(_12609_));
 sky130_fd_sc_hd__xor2_4 _20761_ (.A(net263),
    .B(_12337_),
    .X(_12610_));
 sky130_fd_sc_hd__nand2_1 _20762_ (.A(net300),
    .B(net292),
    .Y(_12611_));
 sky130_fd_sc_hd__nor2_1 _20763_ (.A(net300),
    .B(_11550_),
    .Y(_12612_));
 sky130_fd_sc_hd__nor2_1 _20764_ (.A(_11438_),
    .B(net292),
    .Y(_12613_));
 sky130_fd_sc_hd__or2_2 _20765_ (.A(_12348_),
    .B(_12584_),
    .X(_12614_));
 sky130_fd_sc_hd__mux2_1 _20766_ (.A0(_12612_),
    .A1(_12613_),
    .S(_12614_),
    .X(_12615_));
 sky130_fd_sc_hd__a2bb2o_1 _20767_ (.A1_N(_11608_),
    .A2_N(_12611_),
    .B1(_12615_),
    .B2(net306),
    .X(_12616_));
 sky130_fd_sc_hd__o21ba_1 _20768_ (.A1(_12609_),
    .A2(_12610_),
    .B1_N(_12616_),
    .X(_12617_));
 sky130_fd_sc_hd__a21oi_2 _20769_ (.A1(_12609_),
    .A2(_12610_),
    .B1(_12617_),
    .Y(_12618_));
 sky130_fd_sc_hd__xnor2_1 _20770_ (.A(_12609_),
    .B(_12616_),
    .Y(_12619_));
 sky130_fd_sc_hd__xnor2_2 _20771_ (.A(_12610_),
    .B(_12619_),
    .Y(_12620_));
 sky130_fd_sc_hd__nor2_1 _20772_ (.A(_11527_),
    .B(_12109_),
    .Y(_12621_));
 sky130_fd_sc_hd__xor2_2 _20773_ (.A(_12614_),
    .B(_12621_),
    .X(_12622_));
 sky130_fd_sc_hd__and2_1 _20774_ (.A(net295),
    .B(net278),
    .X(_12623_));
 sky130_fd_sc_hd__nand2_1 _20775_ (.A(net303),
    .B(_12623_),
    .Y(_12624_));
 sky130_fd_sc_hd__xnor2_1 _20776_ (.A(_11608_),
    .B(_12611_),
    .Y(_12625_));
 sky130_fd_sc_hd__nand2_1 _20777_ (.A(_12624_),
    .B(_12625_),
    .Y(_12626_));
 sky130_fd_sc_hd__nor2_1 _20778_ (.A(_12624_),
    .B(_12625_),
    .Y(_12627_));
 sky130_fd_sc_hd__o21a_1 _20779_ (.A1(_12622_),
    .A2(_12627_),
    .B1(_12626_),
    .X(_12628_));
 sky130_fd_sc_hd__o21ai_1 _20780_ (.A1(net299),
    .A2(_12156_),
    .B1(_12611_),
    .Y(_12629_));
 sky130_fd_sc_hd__o21a_1 _20781_ (.A1(_12344_),
    .A2(_12623_),
    .B1(_11438_),
    .X(_12630_));
 sky130_fd_sc_hd__a221o_1 _20782_ (.A1(_12142_),
    .A2(_12623_),
    .B1(_12468_),
    .B2(net299),
    .C1(_12630_),
    .X(_12631_));
 sky130_fd_sc_hd__nor2_1 _20783_ (.A(_11408_),
    .B(_12631_),
    .Y(_12632_));
 sky130_fd_sc_hd__o21a_1 _20784_ (.A1(\top0.cordic0.vec[0][2] ),
    .A2(net285),
    .B1(net278),
    .X(_12633_));
 sky130_fd_sc_hd__o21a_1 _20785_ (.A1(net300),
    .A2(net292),
    .B1(net278),
    .X(_12634_));
 sky130_fd_sc_hd__o22a_1 _20786_ (.A1(_12611_),
    .A2(_12633_),
    .B1(_12634_),
    .B2(net285),
    .X(_12635_));
 sky130_fd_sc_hd__o311a_1 _20787_ (.A1(net299),
    .A2(net288),
    .A3(_12623_),
    .B1(_12635_),
    .C1(_11408_),
    .X(_12636_));
 sky130_fd_sc_hd__o22a_1 _20788_ (.A1(_12308_),
    .A2(_12629_),
    .B1(_12632_),
    .B2(_12636_),
    .X(_12637_));
 sky130_fd_sc_hd__o22a_1 _20789_ (.A1(_12622_),
    .A2(_12626_),
    .B1(_12628_),
    .B2(_12637_),
    .X(_12638_));
 sky130_fd_sc_hd__xnor2_1 _20790_ (.A(_11653_),
    .B(_12273_),
    .Y(_12639_));
 sky130_fd_sc_hd__xnor2_1 _20791_ (.A(_12588_),
    .B(_12639_),
    .Y(_12640_));
 sky130_fd_sc_hd__xor2_1 _20792_ (.A(_12587_),
    .B(_12640_),
    .X(_12641_));
 sky130_fd_sc_hd__xnor2_2 _20793_ (.A(_12598_),
    .B(_12641_),
    .Y(_12642_));
 sky130_fd_sc_hd__inv_2 _20794_ (.A(_12642_),
    .Y(_12643_));
 sky130_fd_sc_hd__a31o_1 _20795_ (.A1(_12618_),
    .A2(_12620_),
    .A3(_12638_),
    .B1(_12643_),
    .X(_12644_));
 sky130_fd_sc_hd__a21o_1 _20796_ (.A1(_12620_),
    .A2(_12638_),
    .B1(_12618_),
    .X(_12645_));
 sky130_fd_sc_hd__nand2_1 _20797_ (.A(_12583_),
    .B(_12605_),
    .Y(_12646_));
 sky130_fd_sc_hd__a21boi_1 _20798_ (.A1(_12644_),
    .A2(_12645_),
    .B1_N(_12646_),
    .Y(_12647_));
 sky130_fd_sc_hd__a211o_1 _20799_ (.A1(_12546_),
    .A2(_12579_),
    .B1(_12606_),
    .C1(_12647_),
    .X(_12648_));
 sky130_fd_sc_hd__a21o_1 _20800_ (.A1(_12575_),
    .A2(_12578_),
    .B1(_12546_),
    .X(_12649_));
 sky130_fd_sc_hd__and2_1 _20801_ (.A(_12552_),
    .B(_12555_),
    .X(_12650_));
 sky130_fd_sc_hd__nor2_1 _20802_ (.A(net254),
    .B(_12559_),
    .Y(_12651_));
 sky130_fd_sc_hd__nand2_1 _20803_ (.A(_11608_),
    .B(_12278_),
    .Y(_12652_));
 sky130_fd_sc_hd__nor2_1 _20804_ (.A(_11673_),
    .B(_12559_),
    .Y(_12653_));
 sky130_fd_sc_hd__or2_1 _20805_ (.A(_11608_),
    .B(_12278_),
    .X(_12654_));
 sky130_fd_sc_hd__o22ai_1 _20806_ (.A1(_12651_),
    .A2(_12652_),
    .B1(_12653_),
    .B2(_12654_),
    .Y(_12655_));
 sky130_fd_sc_hd__a32o_1 _20807_ (.A1(net273),
    .A2(_11673_),
    .A3(_12559_),
    .B1(_12650_),
    .B2(_12655_),
    .X(_12656_));
 sky130_fd_sc_hd__o2111a_1 _20808_ (.A1(net254),
    .A2(_12559_),
    .B1(_12650_),
    .C1(_12652_),
    .D1(_12654_),
    .X(_12657_));
 sky130_fd_sc_hd__a211o_1 _20809_ (.A1(net254),
    .A2(_12559_),
    .B1(_12657_),
    .C1(net285),
    .X(_12658_));
 sky130_fd_sc_hd__o21a_1 _20810_ (.A1(_11571_),
    .A2(_12656_),
    .B1(_12658_),
    .X(_12659_));
 sky130_fd_sc_hd__a31oi_4 _20811_ (.A1(_11608_),
    .A2(net254),
    .A3(_12559_),
    .B1(_12659_),
    .Y(_12660_));
 sky130_fd_sc_hd__a21o_1 _20812_ (.A1(_12648_),
    .A2(_12649_),
    .B1(_12660_),
    .X(_12661_));
 sky130_fd_sc_hd__a211o_1 _20813_ (.A1(_12575_),
    .A2(_12578_),
    .B1(_12606_),
    .C1(_12647_),
    .X(_12662_));
 sky130_fd_sc_hd__a21o_1 _20814_ (.A1(_12579_),
    .A2(_12662_),
    .B1(_12546_),
    .X(_12663_));
 sky130_fd_sc_hd__xnor2_1 _20815_ (.A(_12475_),
    .B(_12486_),
    .Y(_12664_));
 sky130_fd_sc_hd__xnor2_1 _20816_ (.A(_12463_),
    .B(_12664_),
    .Y(_12665_));
 sky130_fd_sc_hd__a32o_1 _20817_ (.A1(_12460_),
    .A2(_12461_),
    .A3(_12540_),
    .B1(_12533_),
    .B2(_12665_),
    .X(_12666_));
 sky130_fd_sc_hd__a221o_1 _20818_ (.A1(_12535_),
    .A2(_12539_),
    .B1(_12661_),
    .B2(_12663_),
    .C1(_12666_),
    .X(_12667_));
 sky130_fd_sc_hd__or2b_1 _20819_ (.A(_12543_),
    .B_N(_12667_),
    .X(_12668_));
 sky130_fd_sc_hd__or3_1 _20820_ (.A(_12172_),
    .B(_12173_),
    .C(_12243_),
    .X(_12669_));
 sky130_fd_sc_hd__nor2_1 _20821_ (.A(_12411_),
    .B(_12414_),
    .Y(_12670_));
 sky130_fd_sc_hd__a21o_1 _20822_ (.A1(_12400_),
    .A2(_12417_),
    .B1(_12670_),
    .X(_12671_));
 sky130_fd_sc_hd__a221o_1 _20823_ (.A1(_12670_),
    .A2(_12400_),
    .B1(_12671_),
    .B2(_12399_),
    .C1(_12408_),
    .X(_12672_));
 sky130_fd_sc_hd__nand2_1 _20824_ (.A(_12669_),
    .B(_12672_),
    .Y(_12673_));
 sky130_fd_sc_hd__a21o_1 _20825_ (.A1(_12420_),
    .A2(_12668_),
    .B1(_12673_),
    .X(_12674_));
 sky130_fd_sc_hd__and2_2 _20826_ (.A(_12244_),
    .B(_12674_),
    .X(_12675_));
 sky130_fd_sc_hd__a31o_1 _20827_ (.A1(_12228_),
    .A2(_12229_),
    .A3(_12240_),
    .B1(_12233_),
    .X(_12676_));
 sky130_fd_sc_hd__o21a_1 _20828_ (.A1(_12230_),
    .A2(_12240_),
    .B1(_12676_),
    .X(_12677_));
 sky130_fd_sc_hd__a21o_1 _20829_ (.A1(_12223_),
    .A2(_12226_),
    .B1(_12217_),
    .X(_12678_));
 sky130_fd_sc_hd__a311o_1 _20830_ (.A1(_12223_),
    .A2(_12226_),
    .A3(_12217_),
    .B1(_12211_),
    .C1(_12210_),
    .X(_12679_));
 sky130_fd_sc_hd__and3_1 _20831_ (.A(_12198_),
    .B(_12200_),
    .C(_12203_),
    .X(_12680_));
 sky130_fd_sc_hd__o21ai_2 _20832_ (.A1(_12209_),
    .A2(_12680_),
    .B1(_12204_),
    .Y(_12681_));
 sky130_fd_sc_hd__nand2_1 _20833_ (.A(net214),
    .B(_12238_),
    .Y(_12682_));
 sky130_fd_sc_hd__nand2_4 _20834_ (.A(net229),
    .B(net221),
    .Y(_12683_));
 sky130_fd_sc_hd__xor2_1 _20835_ (.A(_12682_),
    .B(_12683_),
    .X(_12684_));
 sky130_fd_sc_hd__xor2_2 _20836_ (.A(_12681_),
    .B(_12684_),
    .X(_12685_));
 sky130_fd_sc_hd__a21o_1 _20837_ (.A1(_12678_),
    .A2(_12679_),
    .B1(_12685_),
    .X(_12686_));
 sky130_fd_sc_hd__nand3_2 _20838_ (.A(_12678_),
    .B(_12679_),
    .C(_12685_),
    .Y(_12687_));
 sky130_fd_sc_hd__o21a_1 _20839_ (.A1(net277),
    .A2(_12040_),
    .B1(_12212_),
    .X(_12688_));
 sky130_fd_sc_hd__o2bb2a_1 _20840_ (.A1_N(_12066_),
    .A2_N(_12215_),
    .B1(_12212_),
    .B2(_12040_),
    .X(_12689_));
 sky130_fd_sc_hd__o21ai_1 _20841_ (.A1(_12215_),
    .A2(_12688_),
    .B1(_12689_),
    .Y(_12690_));
 sky130_fd_sc_hd__or2_1 _20842_ (.A(_11593_),
    .B(_12040_),
    .X(_12691_));
 sky130_fd_sc_hd__nand2_1 _20843_ (.A(_11593_),
    .B(_12040_),
    .Y(_12692_));
 sky130_fd_sc_hd__nor3_1 _20844_ (.A(net271),
    .B(_12040_),
    .C(_12215_),
    .Y(_12693_));
 sky130_fd_sc_hd__a41o_1 _20845_ (.A1(net271),
    .A2(_12215_),
    .A3(_12691_),
    .A4(_12692_),
    .B1(_12693_),
    .X(_12694_));
 sky130_fd_sc_hd__a21o_1 _20846_ (.A1(net296),
    .A2(_12690_),
    .B1(_12694_),
    .X(_12695_));
 sky130_fd_sc_hd__nor2b_2 _20847_ (.A(net227),
    .B_N(net218),
    .Y(_12696_));
 sky130_fd_sc_hd__nor2b_2 _20848_ (.A(net213),
    .B_N(net225),
    .Y(_12697_));
 sky130_fd_sc_hd__nor2_1 _20849_ (.A(_12696_),
    .B(_12697_),
    .Y(_12698_));
 sky130_fd_sc_hd__nor2b_2 _20850_ (.A(net238),
    .B_N(net234),
    .Y(_12699_));
 sky130_fd_sc_hd__xnor2_1 _20851_ (.A(net229),
    .B(_12699_),
    .Y(_12700_));
 sky130_fd_sc_hd__xor2_1 _20852_ (.A(_12698_),
    .B(_12700_),
    .X(_12701_));
 sky130_fd_sc_hd__xnor2_1 _20853_ (.A(net229),
    .B(net221),
    .Y(_12702_));
 sky130_fd_sc_hd__nor2_1 _20854_ (.A(net239),
    .B(net235),
    .Y(_12703_));
 sky130_fd_sc_hd__a21oi_1 _20855_ (.A1(net235),
    .A2(_12702_),
    .B1(_12703_),
    .Y(_12704_));
 sky130_fd_sc_hd__nand2_1 _20856_ (.A(net238),
    .B(net234),
    .Y(_12705_));
 sky130_fd_sc_hd__a21o_1 _20857_ (.A1(_12206_),
    .A2(_12705_),
    .B1(net246),
    .X(_12706_));
 sky130_fd_sc_hd__or2b_1 _20858_ (.A(net250),
    .B_N(net259),
    .X(_12707_));
 sky130_fd_sc_hd__a221o_2 _20859_ (.A1(net251),
    .A2(_12039_),
    .B1(_12707_),
    .B2(_12255_),
    .C1(_12085_),
    .X(_12708_));
 sky130_fd_sc_hd__nand3_1 _20860_ (.A(_12704_),
    .B(_12706_),
    .C(_12708_),
    .Y(_12709_));
 sky130_fd_sc_hd__a21o_1 _20861_ (.A1(_12704_),
    .A2(_12706_),
    .B1(_12708_),
    .X(_12710_));
 sky130_fd_sc_hd__nand3_1 _20862_ (.A(_12701_),
    .B(_12709_),
    .C(_12710_),
    .Y(_12711_));
 sky130_fd_sc_hd__a21o_1 _20863_ (.A1(_12709_),
    .A2(_12710_),
    .B1(_12701_),
    .X(_12712_));
 sky130_fd_sc_hd__and2b_1 _20864_ (.A_N(net265),
    .B(net271),
    .X(_12713_));
 sky130_fd_sc_hd__mux2_1 _20865_ (.A0(_12101_),
    .A1(_12713_),
    .S(net291),
    .X(_12714_));
 sky130_fd_sc_hd__xnor2_2 _20866_ (.A(net285),
    .B(net259),
    .Y(_12715_));
 sky130_fd_sc_hd__xnor2_1 _20867_ (.A(_12714_),
    .B(_12715_),
    .Y(_12716_));
 sky130_fd_sc_hd__xnor2_2 _20868_ (.A(_12095_),
    .B(_12716_),
    .Y(_12717_));
 sky130_fd_sc_hd__a21o_1 _20869_ (.A1(_12711_),
    .A2(_12712_),
    .B1(_12717_),
    .X(_12718_));
 sky130_fd_sc_hd__nand3_1 _20870_ (.A(_12717_),
    .B(_12711_),
    .C(_12712_),
    .Y(_12719_));
 sky130_fd_sc_hd__and3_1 _20871_ (.A(_12695_),
    .B(_12718_),
    .C(_12719_),
    .X(_12720_));
 sky130_fd_sc_hd__a21oi_2 _20872_ (.A1(_12718_),
    .A2(_12719_),
    .B1(_12695_),
    .Y(_12721_));
 sky130_fd_sc_hd__a211o_1 _20873_ (.A1(_12686_),
    .A2(_12687_),
    .B1(_12720_),
    .C1(_12721_),
    .X(_12722_));
 sky130_fd_sc_hd__o211ai_1 _20874_ (.A1(_12720_),
    .A2(_12721_),
    .B1(_12686_),
    .C1(_12687_),
    .Y(_12723_));
 sky130_fd_sc_hd__or2_1 _20875_ (.A(_12238_),
    .B(_12236_),
    .X(_12724_));
 sky130_fd_sc_hd__a31o_1 _20876_ (.A1(net235),
    .A2(\top0.cordic0.vec[0][15] ),
    .A3(net214),
    .B1(_12236_),
    .X(_12725_));
 sky130_fd_sc_hd__a22oi_2 _20877_ (.A1(_12724_),
    .A2(_12682_),
    .B1(_12725_),
    .B2(_12165_),
    .Y(_12726_));
 sky130_fd_sc_hd__and3_1 _20878_ (.A(_12722_),
    .B(_12723_),
    .C(_12726_),
    .X(_12727_));
 sky130_fd_sc_hd__a21o_1 _20879_ (.A1(_12722_),
    .A2(_12723_),
    .B1(_12726_),
    .X(_12728_));
 sky130_fd_sc_hd__and2b_1 _20880_ (.A_N(_12727_),
    .B(_12728_),
    .X(_12729_));
 sky130_fd_sc_hd__xnor2_1 _20881_ (.A(_12677_),
    .B(_12729_),
    .Y(_12730_));
 sky130_fd_sc_hd__o21ai_1 _20882_ (.A1(_12161_),
    .A2(_12192_),
    .B1(_12194_),
    .Y(_12731_));
 sky130_fd_sc_hd__o21ai_2 _20883_ (.A1(_12179_),
    .A2(_12242_),
    .B1(_12731_),
    .Y(_12732_));
 sky130_fd_sc_hd__a21oi_1 _20884_ (.A1(_12161_),
    .A2(_12192_),
    .B1(_12187_),
    .Y(_12733_));
 sky130_fd_sc_hd__o21ai_1 _20885_ (.A1(_12179_),
    .A2(_12733_),
    .B1(_12242_),
    .Y(_12734_));
 sky130_fd_sc_hd__o311ai_4 _20886_ (.A1(_12161_),
    .A2(_12187_),
    .A3(_12194_),
    .B1(_12732_),
    .C1(_12734_),
    .Y(_12735_));
 sky130_fd_sc_hd__nor2_2 _20887_ (.A(_12730_),
    .B(_12735_),
    .Y(_12736_));
 sky130_fd_sc_hd__and2_1 _20888_ (.A(_12730_),
    .B(_12735_),
    .X(_12737_));
 sky130_fd_sc_hd__nor2_2 _20889_ (.A(_12736_),
    .B(_12737_),
    .Y(_12738_));
 sky130_fd_sc_hd__xnor2_4 _20890_ (.A(_12675_),
    .B(_12738_),
    .Y(_12739_));
 sky130_fd_sc_hd__clkbuf_4 _20891_ (.A(_12035_),
    .X(_12740_));
 sky130_fd_sc_hd__nor2_1 _20892_ (.A(_12739_),
    .B(_12740_),
    .Y(_12741_));
 sky130_fd_sc_hd__a31o_1 _20893_ (.A1(net732),
    .A2(_12034_),
    .A3(_12037_),
    .B1(_12741_),
    .X(_00383_));
 sky130_fd_sc_hd__nor2_2 _20894_ (.A(_11433_),
    .B(_11648_),
    .Y(_12742_));
 sky130_fd_sc_hd__xnor2_1 _20895_ (.A(\top0.cordic0.domain[0] ),
    .B(net211),
    .Y(_12743_));
 sky130_fd_sc_hd__buf_1 _20896_ (.A(_12743_),
    .X(_12744_));
 sky130_fd_sc_hd__a21oi_1 _20897_ (.A1(_12678_),
    .A2(_12679_),
    .B1(_12685_),
    .Y(_12745_));
 sky130_fd_sc_hd__o31ai_4 _20898_ (.A1(_12720_),
    .A2(_12721_),
    .A3(_12745_),
    .B1(_12687_),
    .Y(_12746_));
 sky130_fd_sc_hd__a31o_1 _20899_ (.A1(net229),
    .A2(net221),
    .A3(net214),
    .B1(_12681_),
    .X(_12747_));
 sky130_fd_sc_hd__mux2_1 _20900_ (.A0(_12681_),
    .A1(_11788_),
    .S(_12683_),
    .X(_12748_));
 sky130_fd_sc_hd__a21o_1 _20901_ (.A1(_12238_),
    .A2(_12747_),
    .B1(_12748_),
    .X(_12749_));
 sky130_fd_sc_hd__nand2_1 _20902_ (.A(_12711_),
    .B(_12712_),
    .Y(_12750_));
 sky130_fd_sc_hd__o21a_1 _20903_ (.A1(_12717_),
    .A2(_12750_),
    .B1(_12695_),
    .X(_12751_));
 sky130_fd_sc_hd__a21oi_2 _20904_ (.A1(_12717_),
    .A2(_12750_),
    .B1(_12751_),
    .Y(_12752_));
 sky130_fd_sc_hd__o21ba_1 _20905_ (.A1(net271),
    .A2(_12095_),
    .B1_N(_12713_),
    .X(_12753_));
 sky130_fd_sc_hd__nand2_1 _20906_ (.A(_12101_),
    .B(_12715_),
    .Y(_12754_));
 sky130_fd_sc_hd__o31a_1 _20907_ (.A1(_11608_),
    .A2(net265),
    .A3(_12095_),
    .B1(_12754_),
    .X(_12755_));
 sky130_fd_sc_hd__o21ai_1 _20908_ (.A1(_12715_),
    .A2(_12753_),
    .B1(_12755_),
    .Y(_12756_));
 sky130_fd_sc_hd__xnor2_1 _20909_ (.A(net271),
    .B(_12095_),
    .Y(_12757_));
 sky130_fd_sc_hd__nor3_1 _20910_ (.A(net265),
    .B(_12095_),
    .C(_12715_),
    .Y(_12758_));
 sky130_fd_sc_hd__a31o_1 _20911_ (.A1(net265),
    .A2(_12715_),
    .A3(_12757_),
    .B1(_12758_),
    .X(_12759_));
 sky130_fd_sc_hd__a21oi_2 _20912_ (.A1(net291),
    .A2(_12756_),
    .B1(_12759_),
    .Y(_12760_));
 sky130_fd_sc_hd__nor2b_4 _20913_ (.A(net229),
    .B_N(net226),
    .Y(_12761_));
 sky130_fd_sc_hd__or2b_1 _20914_ (.A(net218),
    .B_N(net232),
    .X(_12762_));
 sky130_fd_sc_hd__and3b_1 _20915_ (.A_N(_12761_),
    .B(_12762_),
    .C(net241),
    .X(_12763_));
 sky130_fd_sc_hd__nand2b_1 _20916_ (.A_N(net232),
    .B(net218),
    .Y(_12764_));
 sky130_fd_sc_hd__nand2_1 _20917_ (.A(net232),
    .B(net228),
    .Y(_12765_));
 sky130_fd_sc_hd__a21oi_1 _20918_ (.A1(_12764_),
    .A2(_12765_),
    .B1(net241),
    .Y(_12766_));
 sky130_fd_sc_hd__or3b_1 _20919_ (.A(net236),
    .B(_12761_),
    .C_N(_12762_),
    .X(_12767_));
 sky130_fd_sc_hd__o31a_1 _20920_ (.A1(_11726_),
    .A2(_12763_),
    .A3(_12766_),
    .B1(_12767_),
    .X(_12768_));
 sky130_fd_sc_hd__and2b_1 _20921_ (.A_N(net223),
    .B(net218),
    .X(_12769_));
 sky130_fd_sc_hd__and2b_1 _20922_ (.A_N(net218),
    .B(net224),
    .X(_12770_));
 sky130_fd_sc_hd__or2_1 _20923_ (.A(_12769_),
    .B(_12770_),
    .X(_12771_));
 sky130_fd_sc_hd__or2b_1 _20924_ (.A(net244),
    .B_N(net254),
    .X(_12772_));
 sky130_fd_sc_hd__a221o_2 _20925_ (.A1(net244),
    .A2(_12094_),
    .B1(_12772_),
    .B2(_12293_),
    .C1(_12138_),
    .X(_12773_));
 sky130_fd_sc_hd__xnor2_1 _20926_ (.A(_12771_),
    .B(_12773_),
    .Y(_12774_));
 sky130_fd_sc_hd__xnor2_2 _20927_ (.A(_12768_),
    .B(_12774_),
    .Y(_12775_));
 sky130_fd_sc_hd__or2b_1 _20928_ (.A(net261),
    .B_N(net267),
    .X(_12776_));
 sky130_fd_sc_hd__mux2_1 _20929_ (.A0(_12126_),
    .A1(_12776_),
    .S(net284),
    .X(_12777_));
 sky130_fd_sc_hd__xor2_2 _20930_ (.A(net276),
    .B(net256),
    .X(_12778_));
 sky130_fd_sc_hd__xor2_1 _20931_ (.A(_12777_),
    .B(_12778_),
    .X(_12779_));
 sky130_fd_sc_hd__xnor2_2 _20932_ (.A(_12135_),
    .B(_12779_),
    .Y(_12780_));
 sky130_fd_sc_hd__xor2_1 _20933_ (.A(_12775_),
    .B(_12780_),
    .X(_12781_));
 sky130_fd_sc_hd__xnor2_2 _20934_ (.A(_12760_),
    .B(_12781_),
    .Y(_12782_));
 sky130_fd_sc_hd__nand2_1 _20935_ (.A(_12704_),
    .B(_12706_),
    .Y(_12783_));
 sky130_fd_sc_hd__and2_1 _20936_ (.A(_12783_),
    .B(_12708_),
    .X(_12784_));
 sky130_fd_sc_hd__clkbuf_4 _20937_ (.A(_12700_),
    .X(_12785_));
 sky130_fd_sc_hd__or2_1 _20938_ (.A(_12785_),
    .B(_12683_),
    .X(_12786_));
 sky130_fd_sc_hd__nand2_1 _20939_ (.A(_12785_),
    .B(_12683_),
    .Y(_12787_));
 sky130_fd_sc_hd__mux2_1 _20940_ (.A0(_12786_),
    .A1(_12787_),
    .S(_11758_),
    .X(_12788_));
 sky130_fd_sc_hd__mux2_1 _20941_ (.A0(_12786_),
    .A1(_12787_),
    .S(net225),
    .X(_12789_));
 sky130_fd_sc_hd__a21o_1 _20942_ (.A1(net235),
    .A2(_12702_),
    .B1(_12703_),
    .X(_12790_));
 sky130_fd_sc_hd__nor3b_1 _20943_ (.A(_12790_),
    .B(_12708_),
    .C_N(_12706_),
    .Y(_12791_));
 sky130_fd_sc_hd__xnor2_1 _20944_ (.A(_11758_),
    .B(_12683_),
    .Y(_12792_));
 sky130_fd_sc_hd__nand2_1 _20945_ (.A(_12792_),
    .B(_12791_),
    .Y(_12793_));
 sky130_fd_sc_hd__o221a_1 _20946_ (.A1(_12784_),
    .A2(_12788_),
    .B1(_12789_),
    .B2(_12791_),
    .C1(_12793_),
    .X(_12794_));
 sky130_fd_sc_hd__nand2_1 _20947_ (.A(_12783_),
    .B(_12708_),
    .Y(_12795_));
 sky130_fd_sc_hd__or2_1 _20948_ (.A(_11758_),
    .B(_12785_),
    .X(_12796_));
 sky130_fd_sc_hd__nand2_1 _20949_ (.A(_11758_),
    .B(_12785_),
    .Y(_12797_));
 sky130_fd_sc_hd__a311o_1 _20950_ (.A1(_12795_),
    .A2(_12796_),
    .A3(_12797_),
    .B1(_12791_),
    .C1(net213),
    .X(_12798_));
 sky130_fd_sc_hd__or2_1 _20951_ (.A(_12795_),
    .B(_12792_),
    .X(_12799_));
 sky130_fd_sc_hd__o211a_1 _20952_ (.A1(_11788_),
    .A2(_12794_),
    .B1(_12798_),
    .C1(_12799_),
    .X(_12800_));
 sky130_fd_sc_hd__xor2_1 _20953_ (.A(_12782_),
    .B(_12800_),
    .X(_12801_));
 sky130_fd_sc_hd__xnor2_2 _20954_ (.A(_12752_),
    .B(_12801_),
    .Y(_12802_));
 sky130_fd_sc_hd__xnor2_1 _20955_ (.A(_12749_),
    .B(_12802_),
    .Y(_12803_));
 sky130_fd_sc_hd__xnor2_2 _20956_ (.A(_12746_),
    .B(_12803_),
    .Y(_12804_));
 sky130_fd_sc_hd__a21o_1 _20957_ (.A1(_12677_),
    .A2(_12728_),
    .B1(_12727_),
    .X(_12805_));
 sky130_fd_sc_hd__xnor2_2 _20958_ (.A(_12804_),
    .B(_12805_),
    .Y(_12806_));
 sky130_fd_sc_hd__inv_2 _20959_ (.A(_12737_),
    .Y(_12807_));
 sky130_fd_sc_hd__o21a_2 _20960_ (.A1(_12675_),
    .A2(_12736_),
    .B1(_12807_),
    .X(_12808_));
 sky130_fd_sc_hd__xor2_2 _20961_ (.A(_12806_),
    .B(_12808_),
    .X(_12809_));
 sky130_fd_sc_hd__or3_1 _20962_ (.A(_12739_),
    .B(net1021),
    .C(_12809_),
    .X(_12810_));
 sky130_fd_sc_hd__o21ai_1 _20963_ (.A1(_12739_),
    .A2(net1021),
    .B1(_12809_),
    .Y(_12811_));
 sky130_fd_sc_hd__and2_1 _20964_ (.A(_12003_),
    .B(_12035_),
    .X(_12812_));
 sky130_fd_sc_hd__clkbuf_4 _20965_ (.A(_12812_),
    .X(_12813_));
 sky130_fd_sc_hd__a32o_1 _20966_ (.A1(_12742_),
    .A2(_12810_),
    .A3(_12811_),
    .B1(_12813_),
    .B2(net715),
    .X(_00384_));
 sky130_fd_sc_hd__nor2_1 _20967_ (.A(net236),
    .B(net231),
    .Y(_12814_));
 sky130_fd_sc_hd__nor2_1 _20968_ (.A(_11726_),
    .B(_11739_),
    .Y(_12815_));
 sky130_fd_sc_hd__o21ba_1 _20969_ (.A1(_12698_),
    .A2(_12815_),
    .B1_N(net241),
    .X(_12816_));
 sky130_fd_sc_hd__a211o_1 _20970_ (.A1(net231),
    .A2(_12698_),
    .B1(_12814_),
    .C1(_12816_),
    .X(_12817_));
 sky130_fd_sc_hd__nand2_1 _20971_ (.A(_12773_),
    .B(_12817_),
    .Y(_12818_));
 sky130_fd_sc_hd__nand2_1 _20972_ (.A(_11726_),
    .B(net230),
    .Y(_12819_));
 sky130_fd_sc_hd__nor2_2 _20973_ (.A(net236),
    .B(_11739_),
    .Y(_12820_));
 sky130_fd_sc_hd__or3_1 _20974_ (.A(net222),
    .B(net213),
    .C(_12820_),
    .X(_12821_));
 sky130_fd_sc_hd__o21ai_1 _20975_ (.A1(_12072_),
    .A2(_12819_),
    .B1(_12821_),
    .Y(_12822_));
 sky130_fd_sc_hd__xnor2_1 _20976_ (.A(_12072_),
    .B(_12820_),
    .Y(_12823_));
 sky130_fd_sc_hd__nor2_1 _20977_ (.A(net227),
    .B(net219),
    .Y(_12824_));
 sky130_fd_sc_hd__a22o_1 _20978_ (.A1(net227),
    .A2(_12822_),
    .B1(_12823_),
    .B2(_12824_),
    .X(_12825_));
 sky130_fd_sc_hd__nor2_1 _20979_ (.A(net225),
    .B(net222),
    .Y(_12826_));
 sky130_fd_sc_hd__or2_1 _20980_ (.A(_12817_),
    .B(_12820_),
    .X(_12827_));
 sky130_fd_sc_hd__and3_1 _20981_ (.A(net225),
    .B(net222),
    .C(_12817_),
    .X(_12828_));
 sky130_fd_sc_hd__a21o_1 _20982_ (.A1(_12826_),
    .A2(_12827_),
    .B1(_12828_),
    .X(_12829_));
 sky130_fd_sc_hd__nor2_1 _20983_ (.A(_12826_),
    .B(_12819_),
    .Y(_12830_));
 sky130_fd_sc_hd__a22o_1 _20984_ (.A1(_12773_),
    .A2(_12829_),
    .B1(_12830_),
    .B2(_12818_),
    .X(_12831_));
 sky130_fd_sc_hd__nand2_1 _20985_ (.A(_11757_),
    .B(net221),
    .Y(_12832_));
 sky130_fd_sc_hd__nand2_1 _20986_ (.A(net227),
    .B(_12180_),
    .Y(_12833_));
 sky130_fd_sc_hd__a311oi_1 _20987_ (.A1(net213),
    .A2(_12832_),
    .A3(_12833_),
    .B1(_12817_),
    .C1(_12773_),
    .Y(_12834_));
 sky130_fd_sc_hd__a221o_2 _20988_ (.A1(_12818_),
    .A2(_12825_),
    .B1(_12831_),
    .B2(net213),
    .C1(_12834_),
    .X(_12835_));
 sky130_fd_sc_hd__nor2_1 _20989_ (.A(net262),
    .B(_12135_),
    .Y(_12836_));
 sky130_fd_sc_hd__or2_1 _20990_ (.A(net267),
    .B(_12135_),
    .X(_12837_));
 sky130_fd_sc_hd__nand2_1 _20991_ (.A(_12776_),
    .B(_12837_),
    .Y(_12838_));
 sky130_fd_sc_hd__nor2_1 _20992_ (.A(_12126_),
    .B(_12778_),
    .Y(_12839_));
 sky130_fd_sc_hd__a221o_1 _20993_ (.A1(net267),
    .A2(_12836_),
    .B1(_12838_),
    .B2(_12778_),
    .C1(_12839_),
    .X(_12840_));
 sky130_fd_sc_hd__nand2_1 _20994_ (.A(net267),
    .B(_12135_),
    .Y(_12841_));
 sky130_fd_sc_hd__a211oi_1 _20995_ (.A1(_12837_),
    .A2(_12841_),
    .B1(_11653_),
    .C1(_12778_),
    .Y(_12842_));
 sky130_fd_sc_hd__a221o_2 _20996_ (.A1(_12778_),
    .A2(_12836_),
    .B1(_12840_),
    .B2(net284),
    .C1(_12842_),
    .X(_12843_));
 sky130_fd_sc_hd__or2b_1 _20997_ (.A(net255),
    .B_N(net259),
    .X(_12844_));
 sky130_fd_sc_hd__or3b_1 _20998_ (.A(net277),
    .B(net259),
    .C_N(net255),
    .X(_12845_));
 sky130_fd_sc_hd__o21a_1 _20999_ (.A1(_11592_),
    .A2(_12844_),
    .B1(_12845_),
    .X(_12846_));
 sky130_fd_sc_hd__xor2_2 _21000_ (.A(net271),
    .B(net251),
    .X(_12847_));
 sky130_fd_sc_hd__xor2_1 _21001_ (.A(_12846_),
    .B(_12847_),
    .X(_12848_));
 sky130_fd_sc_hd__xnor2_1 _21002_ (.A(_12208_),
    .B(_12848_),
    .Y(_12849_));
 sky130_fd_sc_hd__or2_1 _21003_ (.A(_11689_),
    .B(net238),
    .X(_12850_));
 sky130_fd_sc_hd__a221o_4 _21004_ (.A1(net238),
    .A2(_12134_),
    .B1(_12269_),
    .B2(_12850_),
    .C1(_12197_),
    .X(_12851_));
 sky130_fd_sc_hd__a211o_1 _21005_ (.A1(net225),
    .A2(net221),
    .B1(_12696_),
    .C1(net234),
    .X(_12852_));
 sky130_fd_sc_hd__nor2b_2 _21006_ (.A(net225),
    .B_N(net222),
    .Y(_12853_));
 sky130_fd_sc_hd__o21ai_1 _21007_ (.A1(_12697_),
    .A2(_12853_),
    .B1(net234),
    .Y(_12854_));
 sky130_fd_sc_hd__o21a_1 _21008_ (.A1(_12697_),
    .A2(_12853_),
    .B1(_11739_),
    .X(_12855_));
 sky130_fd_sc_hd__a31o_1 _21009_ (.A1(net229),
    .A2(_12852_),
    .A3(_12854_),
    .B1(_12855_),
    .X(_12856_));
 sky130_fd_sc_hd__xor2_2 _21010_ (.A(_12851_),
    .B(_12856_),
    .X(_12857_));
 sky130_fd_sc_hd__and2_1 _21011_ (.A(_12849_),
    .B(_12857_),
    .X(_12858_));
 sky130_fd_sc_hd__nor2_1 _21012_ (.A(_12849_),
    .B(_12857_),
    .Y(_12859_));
 sky130_fd_sc_hd__nor2_1 _21013_ (.A(_12858_),
    .B(_12859_),
    .Y(_12860_));
 sky130_fd_sc_hd__xnor2_2 _21014_ (.A(_12843_),
    .B(_12860_),
    .Y(_12861_));
 sky130_fd_sc_hd__o21a_1 _21015_ (.A1(_12775_),
    .A2(_12780_),
    .B1(_12760_),
    .X(_12862_));
 sky130_fd_sc_hd__a21o_1 _21016_ (.A1(_12775_),
    .A2(_12780_),
    .B1(_12862_),
    .X(_12863_));
 sky130_fd_sc_hd__xnor2_2 _21017_ (.A(_12861_),
    .B(_12863_),
    .Y(_12864_));
 sky130_fd_sc_hd__xnor2_4 _21018_ (.A(_12835_),
    .B(_12864_),
    .Y(_12865_));
 sky130_fd_sc_hd__nor2_1 _21019_ (.A(_12782_),
    .B(_12800_),
    .Y(_12866_));
 sky130_fd_sc_hd__nand2_1 _21020_ (.A(_12782_),
    .B(_12800_),
    .Y(_12867_));
 sky130_fd_sc_hd__o21ai_2 _21021_ (.A1(_12752_),
    .A2(_12866_),
    .B1(_12867_),
    .Y(_12868_));
 sky130_fd_sc_hd__inv_2 _21022_ (.A(_12785_),
    .Y(_12869_));
 sky130_fd_sc_hd__o21a_1 _21023_ (.A1(_12869_),
    .A2(_12783_),
    .B1(_12708_),
    .X(_12870_));
 sky130_fd_sc_hd__a211o_1 _21024_ (.A1(_12869_),
    .A2(_12783_),
    .B1(_12870_),
    .C1(net225),
    .X(_12871_));
 sky130_fd_sc_hd__a21oi_1 _21025_ (.A1(_12869_),
    .A2(_12795_),
    .B1(_11759_),
    .Y(_12872_));
 sky130_fd_sc_hd__a211oi_4 _21026_ (.A1(_12683_),
    .A2(_12871_),
    .B1(_12872_),
    .C1(_11789_),
    .Y(_12873_));
 sky130_fd_sc_hd__xnor2_2 _21027_ (.A(_12868_),
    .B(_12873_),
    .Y(_12874_));
 sky130_fd_sc_hd__xnor2_4 _21028_ (.A(_12865_),
    .B(_12874_),
    .Y(_12875_));
 sky130_fd_sc_hd__o21ba_1 _21029_ (.A1(_12749_),
    .A2(_12746_),
    .B1_N(_12802_),
    .X(_12876_));
 sky130_fd_sc_hd__a21oi_2 _21030_ (.A1(_12749_),
    .A2(_12746_),
    .B1(_12876_),
    .Y(_12877_));
 sky130_fd_sc_hd__xnor2_4 _21031_ (.A(_12875_),
    .B(_12877_),
    .Y(_12878_));
 sky130_fd_sc_hd__or2_1 _21032_ (.A(_12804_),
    .B(_12805_),
    .X(_12879_));
 sky130_fd_sc_hd__or2_1 _21033_ (.A(_12675_),
    .B(_12807_),
    .X(_12880_));
 sky130_fd_sc_hd__and2_1 _21034_ (.A(_12804_),
    .B(_12805_),
    .X(_12881_));
 sky130_fd_sc_hd__o21a_1 _21035_ (.A1(_12808_),
    .A2(_12881_),
    .B1(_12879_),
    .X(_12882_));
 sky130_fd_sc_hd__inv_2 _21036_ (.A(_12743_),
    .Y(_12883_));
 sky130_fd_sc_hd__a21o_1 _21037_ (.A1(_12736_),
    .A2(_12879_),
    .B1(_12881_),
    .X(_12884_));
 sky130_fd_sc_hd__a22o_1 _21038_ (.A1(_12807_),
    .A2(_12881_),
    .B1(_12884_),
    .B2(_12675_),
    .X(_12885_));
 sky130_fd_sc_hd__nand2_1 _21039_ (.A(_12883_),
    .B(_12885_),
    .Y(_12886_));
 sky130_fd_sc_hd__o221a_1 _21040_ (.A1(_12879_),
    .A2(_12880_),
    .B1(_12882_),
    .B2(_12883_),
    .C1(_12886_),
    .X(_12887_));
 sky130_fd_sc_hd__xor2_2 _21041_ (.A(_12878_),
    .B(_12887_),
    .X(_12888_));
 sky130_fd_sc_hd__nor2_1 _21042_ (.A(_12740_),
    .B(_12888_),
    .Y(_12889_));
 sky130_fd_sc_hd__a31o_1 _21043_ (.A1(net756),
    .A2(_12034_),
    .A3(_12037_),
    .B1(_12889_),
    .X(_00385_));
 sky130_fd_sc_hd__or2b_1 _21044_ (.A(_12863_),
    .B_N(_12835_),
    .X(_12890_));
 sky130_fd_sc_hd__and2b_1 _21045_ (.A_N(_12835_),
    .B(_12863_),
    .X(_12891_));
 sky130_fd_sc_hd__a21o_1 _21046_ (.A1(_12861_),
    .A2(_12890_),
    .B1(_12891_),
    .X(_12892_));
 sky130_fd_sc_hd__nor2_1 _21047_ (.A(_11758_),
    .B(_12820_),
    .Y(_12893_));
 sky130_fd_sc_hd__nor2_1 _21048_ (.A(_12180_),
    .B(_12893_),
    .Y(_12894_));
 sky130_fd_sc_hd__a21o_1 _21049_ (.A1(net221),
    .A2(_12827_),
    .B1(_11759_),
    .X(_12895_));
 sky130_fd_sc_hd__o221a_1 _21050_ (.A1(net222),
    .A2(_12827_),
    .B1(_12894_),
    .B2(_12773_),
    .C1(_12895_),
    .X(_12896_));
 sky130_fd_sc_hd__or2_1 _21051_ (.A(_11789_),
    .B(_12896_),
    .X(_12897_));
 sky130_fd_sc_hd__nand2_1 _21052_ (.A(_12849_),
    .B(_12857_),
    .Y(_12898_));
 sky130_fd_sc_hd__a21oi_2 _21053_ (.A1(_12843_),
    .A2(_12898_),
    .B1(_12859_),
    .Y(_12899_));
 sky130_fd_sc_hd__nor2_1 _21054_ (.A(net255),
    .B(_12208_),
    .Y(_12900_));
 sky130_fd_sc_hd__nor2_1 _21055_ (.A(_12039_),
    .B(_12847_),
    .Y(_12901_));
 sky130_fd_sc_hd__or2_1 _21056_ (.A(net262),
    .B(_12208_),
    .X(_12902_));
 sky130_fd_sc_hd__and3_1 _21057_ (.A(_12844_),
    .B(_12847_),
    .C(_12902_),
    .X(_12903_));
 sky130_fd_sc_hd__o2bb2a_1 _21058_ (.A1_N(net259),
    .A2_N(_12900_),
    .B1(_12901_),
    .B2(_12903_),
    .X(_12904_));
 sky130_fd_sc_hd__nand2_1 _21059_ (.A(net262),
    .B(_12208_),
    .Y(_12905_));
 sky130_fd_sc_hd__a21o_1 _21060_ (.A1(_12902_),
    .A2(_12905_),
    .B1(_11673_),
    .X(_12906_));
 sky130_fd_sc_hd__nand2_1 _21061_ (.A(_12847_),
    .B(_12900_),
    .Y(_12907_));
 sky130_fd_sc_hd__o221a_1 _21062_ (.A1(_11593_),
    .A2(_12904_),
    .B1(_12906_),
    .B2(_12847_),
    .C1(_12907_),
    .X(_12908_));
 sky130_fd_sc_hd__a21oi_1 _21063_ (.A1(net247),
    .A2(_11726_),
    .B1(_12045_),
    .Y(_12909_));
 sky130_fd_sc_hd__a211o_2 _21064_ (.A1(net235),
    .A2(_12207_),
    .B1(_12703_),
    .C1(_12909_),
    .X(_12910_));
 sky130_fd_sc_hd__nand2_1 _21065_ (.A(net230),
    .B(_12072_),
    .Y(_12911_));
 sky130_fd_sc_hd__o21a_1 _21066_ (.A1(_11757_),
    .A2(_12911_),
    .B1(_12832_),
    .X(_12912_));
 sky130_fd_sc_hd__xnor2_1 _21067_ (.A(_11787_),
    .B(_12912_),
    .Y(_12913_));
 sky130_fd_sc_hd__xnor2_2 _21068_ (.A(_12910_),
    .B(_12913_),
    .Y(_12914_));
 sky130_fd_sc_hd__nor2_1 _21069_ (.A(_11672_),
    .B(net251),
    .Y(_12915_));
 sky130_fd_sc_hd__mux2_1 _21070_ (.A0(_12094_),
    .A1(_12915_),
    .S(net272),
    .X(_12916_));
 sky130_fd_sc_hd__xnor2_2 _21071_ (.A(net265),
    .B(net244),
    .Y(_12917_));
 sky130_fd_sc_hd__xor2_1 _21072_ (.A(_12785_),
    .B(_12917_),
    .X(_12918_));
 sky130_fd_sc_hd__xnor2_2 _21073_ (.A(_12916_),
    .B(_12918_),
    .Y(_12919_));
 sky130_fd_sc_hd__xor2_1 _21074_ (.A(_12914_),
    .B(_12919_),
    .X(_12920_));
 sky130_fd_sc_hd__xnor2_2 _21075_ (.A(_12908_),
    .B(_12920_),
    .Y(_12921_));
 sky130_fd_sc_hd__nor2_1 _21076_ (.A(net234),
    .B(_12696_),
    .Y(_12922_));
 sky130_fd_sc_hd__or3_1 _21077_ (.A(_12697_),
    .B(_12851_),
    .C(_12922_),
    .X(_12923_));
 sky130_fd_sc_hd__nor2_1 _21078_ (.A(_11726_),
    .B(net226),
    .Y(_12924_));
 sky130_fd_sc_hd__or2b_1 _21079_ (.A(_12924_),
    .B_N(_12851_),
    .X(_12925_));
 sky130_fd_sc_hd__nor2_1 _21080_ (.A(_12072_),
    .B(_11788_),
    .Y(_12926_));
 sky130_fd_sc_hd__a221o_1 _21081_ (.A1(_12180_),
    .A2(_12923_),
    .B1(_12925_),
    .B2(_12926_),
    .C1(_11739_),
    .X(_12927_));
 sky130_fd_sc_hd__o21ai_1 _21082_ (.A1(_11788_),
    .A2(_12851_),
    .B1(net221),
    .Y(_12928_));
 sky130_fd_sc_hd__a221o_1 _21083_ (.A1(_11788_),
    .A2(_12851_),
    .B1(_12928_),
    .B2(_11758_),
    .C1(net229),
    .X(_12929_));
 sky130_fd_sc_hd__and4_1 _21084_ (.A(_11727_),
    .B(net225),
    .C(_11788_),
    .D(_12851_),
    .X(_12930_));
 sky130_fd_sc_hd__a21oi_2 _21085_ (.A1(_12927_),
    .A2(_12929_),
    .B1(_12930_),
    .Y(_12931_));
 sky130_fd_sc_hd__xnor2_1 _21086_ (.A(_12921_),
    .B(_12931_),
    .Y(_12932_));
 sky130_fd_sc_hd__xnor2_2 _21087_ (.A(_12899_),
    .B(_12932_),
    .Y(_12933_));
 sky130_fd_sc_hd__xnor2_1 _21088_ (.A(_12897_),
    .B(_12933_),
    .Y(_12934_));
 sky130_fd_sc_hd__xnor2_1 _21089_ (.A(_12892_),
    .B(_12934_),
    .Y(_12935_));
 sky130_fd_sc_hd__o21a_1 _21090_ (.A1(_12865_),
    .A2(_12873_),
    .B1(_12868_),
    .X(_12936_));
 sky130_fd_sc_hd__a21oi_1 _21091_ (.A1(_12865_),
    .A2(_12873_),
    .B1(_12936_),
    .Y(_12937_));
 sky130_fd_sc_hd__and2_1 _21092_ (.A(_12935_),
    .B(_12937_),
    .X(_12938_));
 sky130_fd_sc_hd__or2_1 _21093_ (.A(_12935_),
    .B(_12937_),
    .X(_12939_));
 sky130_fd_sc_hd__or2b_1 _21094_ (.A(_12938_),
    .B_N(_12939_),
    .X(_12940_));
 sky130_fd_sc_hd__or2_1 _21095_ (.A(_12806_),
    .B(_12878_),
    .X(_12941_));
 sky130_fd_sc_hd__inv_2 _21096_ (.A(_12941_),
    .Y(_12942_));
 sky130_fd_sc_hd__a21oi_2 _21097_ (.A1(_12677_),
    .A2(_12728_),
    .B1(_12727_),
    .Y(_12943_));
 sky130_fd_sc_hd__nand2_1 _21098_ (.A(_12746_),
    .B(_12943_),
    .Y(_12944_));
 sky130_fd_sc_hd__nor2_1 _21099_ (.A(_12746_),
    .B(_12943_),
    .Y(_12945_));
 sky130_fd_sc_hd__and2b_1 _21100_ (.A_N(_12749_),
    .B(_12802_),
    .X(_12946_));
 sky130_fd_sc_hd__o21a_1 _21101_ (.A1(_12875_),
    .A2(_12945_),
    .B1(_12946_),
    .X(_12947_));
 sky130_fd_sc_hd__a21oi_1 _21102_ (.A1(_12746_),
    .A2(_12943_),
    .B1(_12749_),
    .Y(_12948_));
 sky130_fd_sc_hd__o21a_1 _21103_ (.A1(_12945_),
    .A2(_12948_),
    .B1(_12875_),
    .X(_12949_));
 sky130_fd_sc_hd__a311oi_2 _21104_ (.A1(_12802_),
    .A2(_12875_),
    .A3(_12944_),
    .B1(_12947_),
    .C1(_12949_),
    .Y(_12950_));
 sky130_fd_sc_hd__a21boi_2 _21105_ (.A1(_12808_),
    .A2(_12942_),
    .B1_N(_12950_),
    .Y(_12951_));
 sky130_fd_sc_hd__xor2_2 _21106_ (.A(_12940_),
    .B(_12951_),
    .X(_12952_));
 sky130_fd_sc_hd__inv_2 _21107_ (.A(_12736_),
    .Y(_12953_));
 sky130_fd_sc_hd__inv_2 _21108_ (.A(_12738_),
    .Y(_12954_));
 sky130_fd_sc_hd__mux2_1 _21109_ (.A0(_12953_),
    .A1(_12954_),
    .S(_12675_),
    .X(_12955_));
 sky130_fd_sc_hd__or3b_1 _21110_ (.A(_12805_),
    .B(_12880_),
    .C_N(_12878_),
    .X(_12956_));
 sky130_fd_sc_hd__o31ai_1 _21111_ (.A1(_12943_),
    .A2(_12878_),
    .A3(_12955_),
    .B1(_12956_),
    .Y(_12957_));
 sky130_fd_sc_hd__mux2_1 _21112_ (.A0(_12880_),
    .A1(_12955_),
    .S(_12943_),
    .X(_12958_));
 sky130_fd_sc_hd__nor2_1 _21113_ (.A(_12878_),
    .B(_12958_),
    .Y(_12959_));
 sky130_fd_sc_hd__mux2_1 _21114_ (.A0(_12957_),
    .A1(_12959_),
    .S(_12804_),
    .X(_12960_));
 sky130_fd_sc_hd__or2_1 _21115_ (.A(net1021),
    .B(_12960_),
    .X(_12961_));
 sky130_fd_sc_hd__xnor2_2 _21116_ (.A(_12952_),
    .B(_12961_),
    .Y(_12962_));
 sky130_fd_sc_hd__clkbuf_4 _21117_ (.A(_12742_),
    .X(_12963_));
 sky130_fd_sc_hd__a22o_1 _21118_ (.A1(net718),
    .A2(_12813_),
    .B1(_12962_),
    .B2(_12963_),
    .X(_00386_));
 sky130_fd_sc_hd__o21a_1 _21119_ (.A1(_12897_),
    .A2(_12933_),
    .B1(_12892_),
    .X(_12964_));
 sky130_fd_sc_hd__a21oi_2 _21120_ (.A1(_12897_),
    .A2(_12933_),
    .B1(_12964_),
    .Y(_12965_));
 sky130_fd_sc_hd__a21o_1 _21121_ (.A1(_12914_),
    .A2(_12919_),
    .B1(_12908_),
    .X(_12966_));
 sky130_fd_sc_hd__o21ai_2 _21122_ (.A1(_12914_),
    .A2(_12919_),
    .B1(_12966_),
    .Y(_12967_));
 sky130_fd_sc_hd__or2_2 _21123_ (.A(_11788_),
    .B(_12765_),
    .X(_12968_));
 sky130_fd_sc_hd__o21ai_1 _21124_ (.A1(net227),
    .A2(_12910_),
    .B1(_12968_),
    .Y(_12969_));
 sky130_fd_sc_hd__nor3b_1 _21125_ (.A(_11759_),
    .B(_12910_),
    .C_N(_12911_),
    .Y(_12970_));
 sky130_fd_sc_hd__a221o_1 _21126_ (.A1(_11788_),
    .A2(_12910_),
    .B1(_12969_),
    .B2(_12180_),
    .C1(_12970_),
    .X(_12971_));
 sky130_fd_sc_hd__nor2_1 _21127_ (.A(net251),
    .B(_12785_),
    .Y(_12972_));
 sky130_fd_sc_hd__nor2_1 _21128_ (.A(net255),
    .B(_12785_),
    .Y(_12973_));
 sky130_fd_sc_hd__o21ba_1 _21129_ (.A1(_12915_),
    .A2(_12973_),
    .B1_N(_12917_),
    .X(_12974_));
 sky130_fd_sc_hd__a221o_1 _21130_ (.A1(_12094_),
    .A2(_12917_),
    .B1(_12972_),
    .B2(net255),
    .C1(_12974_),
    .X(_12975_));
 sky130_fd_sc_hd__nand2_1 _21131_ (.A(_11673_),
    .B(_12785_),
    .Y(_12976_));
 sky130_fd_sc_hd__or2_1 _21132_ (.A(_11673_),
    .B(_12785_),
    .X(_12977_));
 sky130_fd_sc_hd__and2b_1 _21133_ (.A_N(_12917_),
    .B(_12972_),
    .X(_12978_));
 sky130_fd_sc_hd__a41o_1 _21134_ (.A1(net251),
    .A2(_12917_),
    .A3(_12976_),
    .A4(_12977_),
    .B1(_12978_),
    .X(_12979_));
 sky130_fd_sc_hd__a21oi_2 _21135_ (.A1(net272),
    .A2(_12975_),
    .B1(_12979_),
    .Y(_12980_));
 sky130_fd_sc_hd__nor2_1 _21136_ (.A(_11739_),
    .B(net228),
    .Y(_12981_));
 sky130_fd_sc_hd__a21oi_4 _21137_ (.A1(_11727_),
    .A2(_12981_),
    .B1(_12893_),
    .Y(_12982_));
 sky130_fd_sc_hd__nor2_1 _21138_ (.A(_11689_),
    .B(net246),
    .Y(_12983_));
 sky130_fd_sc_hd__mux2_1 _21139_ (.A0(_12134_),
    .A1(_12983_),
    .S(net267),
    .X(_12984_));
 sky130_fd_sc_hd__xnor2_2 _21140_ (.A(net262),
    .B(net238),
    .Y(_12985_));
 sky130_fd_sc_hd__xor2_1 _21141_ (.A(_12984_),
    .B(_12985_),
    .X(_12986_));
 sky130_fd_sc_hd__xnor2_2 _21142_ (.A(_12982_),
    .B(_12986_),
    .Y(_12987_));
 sky130_fd_sc_hd__nand2_1 _21143_ (.A(net257),
    .B(net251),
    .Y(_12988_));
 sky130_fd_sc_hd__nand2_1 _21144_ (.A(net242),
    .B(_11739_),
    .Y(_12989_));
 sky130_fd_sc_hd__a221o_1 _21145_ (.A1(_12988_),
    .A2(_12989_),
    .B1(_12699_),
    .B2(net231),
    .C1(_12814_),
    .X(_12990_));
 sky130_fd_sc_hd__or2_1 _21146_ (.A(_12180_),
    .B(_12824_),
    .X(_12991_));
 sky130_fd_sc_hd__xnor2_1 _21147_ (.A(_12990_),
    .B(_12991_),
    .Y(_12992_));
 sky130_fd_sc_hd__xnor2_1 _21148_ (.A(_12987_),
    .B(_12992_),
    .Y(_12993_));
 sky130_fd_sc_hd__xnor2_1 _21149_ (.A(_12980_),
    .B(_12993_),
    .Y(_12994_));
 sky130_fd_sc_hd__nor2_1 _21150_ (.A(_12971_),
    .B(_12994_),
    .Y(_12995_));
 sky130_fd_sc_hd__nand2_1 _21151_ (.A(_12971_),
    .B(_12994_),
    .Y(_12996_));
 sky130_fd_sc_hd__or2b_1 _21152_ (.A(_12995_),
    .B_N(_12996_),
    .X(_12997_));
 sky130_fd_sc_hd__xnor2_2 _21153_ (.A(_12967_),
    .B(_12997_),
    .Y(_12998_));
 sky130_fd_sc_hd__o21ba_1 _21154_ (.A1(_12921_),
    .A2(_12931_),
    .B1_N(_12899_),
    .X(_12999_));
 sky130_fd_sc_hd__a21o_1 _21155_ (.A1(_12921_),
    .A2(_12931_),
    .B1(_12999_),
    .X(_13000_));
 sky130_fd_sc_hd__nand2_2 _21156_ (.A(net223),
    .B(net219),
    .Y(_13001_));
 sky130_fd_sc_hd__o2bb2a_1 _21157_ (.A1_N(net230),
    .A2_N(_12925_),
    .B1(_12851_),
    .B2(net225),
    .X(_13002_));
 sky130_fd_sc_hd__nor2_1 _21158_ (.A(_13001_),
    .B(_13002_),
    .Y(_13003_));
 sky130_fd_sc_hd__and2_1 _21159_ (.A(_13000_),
    .B(_13003_),
    .X(_13004_));
 sky130_fd_sc_hd__or2_1 _21160_ (.A(_13000_),
    .B(_13003_),
    .X(_13005_));
 sky130_fd_sc_hd__or2b_1 _21161_ (.A(_13004_),
    .B_N(_13005_),
    .X(_13006_));
 sky130_fd_sc_hd__xnor2_2 _21162_ (.A(_12998_),
    .B(_13006_),
    .Y(_13007_));
 sky130_fd_sc_hd__xnor2_2 _21163_ (.A(_12965_),
    .B(_13007_),
    .Y(_13008_));
 sky130_fd_sc_hd__a21oi_1 _21164_ (.A1(_12939_),
    .A2(_12951_),
    .B1(_12938_),
    .Y(_13009_));
 sky130_fd_sc_hd__xor2_2 _21165_ (.A(_13008_),
    .B(_13009_),
    .X(_13010_));
 sky130_fd_sc_hd__inv_2 _21166_ (.A(_12960_),
    .Y(_13011_));
 sky130_fd_sc_hd__o21a_1 _21167_ (.A1(_12952_),
    .A2(_13011_),
    .B1(_12883_),
    .X(_13012_));
 sky130_fd_sc_hd__xnor2_2 _21168_ (.A(_13010_),
    .B(_13012_),
    .Y(_13013_));
 sky130_fd_sc_hd__a22o_1 _21169_ (.A1(net731),
    .A2(_12813_),
    .B1(_13013_),
    .B2(_12963_),
    .X(_00387_));
 sky130_fd_sc_hd__and3b_1 _21170_ (.A_N(_12952_),
    .B(_12960_),
    .C(_13010_),
    .X(_13014_));
 sky130_fd_sc_hd__nor2_1 _21171_ (.A(net1021),
    .B(_13014_),
    .Y(_13015_));
 sky130_fd_sc_hd__a21oi_2 _21172_ (.A1(_12998_),
    .A2(_13005_),
    .B1(_13004_),
    .Y(_13016_));
 sky130_fd_sc_hd__o21a_1 _21173_ (.A1(_12987_),
    .A2(_12992_),
    .B1(_12980_),
    .X(_13017_));
 sky130_fd_sc_hd__a21o_1 _21174_ (.A1(_12987_),
    .A2(_12992_),
    .B1(_13017_),
    .X(_13018_));
 sky130_fd_sc_hd__nor2_1 _21175_ (.A(net246),
    .B(_12982_),
    .Y(_13019_));
 sky130_fd_sc_hd__nor2_1 _21176_ (.A(net252),
    .B(_12982_),
    .Y(_13020_));
 sky130_fd_sc_hd__o21ba_1 _21177_ (.A1(_12983_),
    .A2(_13020_),
    .B1_N(_12985_),
    .X(_13021_));
 sky130_fd_sc_hd__a221o_1 _21178_ (.A1(_12134_),
    .A2(_12985_),
    .B1(_13019_),
    .B2(net252),
    .C1(_13021_),
    .X(_13022_));
 sky130_fd_sc_hd__nand2_1 _21179_ (.A(_11689_),
    .B(_12982_),
    .Y(_13023_));
 sky130_fd_sc_hd__or2_1 _21180_ (.A(_11689_),
    .B(_12982_),
    .X(_13024_));
 sky130_fd_sc_hd__and2b_1 _21181_ (.A_N(_12985_),
    .B(_13019_),
    .X(_13025_));
 sky130_fd_sc_hd__a41o_1 _21182_ (.A1(net246),
    .A2(_12985_),
    .A3(_13023_),
    .A4(_13024_),
    .B1(_13025_),
    .X(_13026_));
 sky130_fd_sc_hd__a21oi_2 _21183_ (.A1(net267),
    .A2(_13022_),
    .B1(_13026_),
    .Y(_13027_));
 sky130_fd_sc_hd__xnor2_2 _21184_ (.A(net221),
    .B(_12761_),
    .Y(_13028_));
 sky130_fd_sc_hd__and2b_1 _21185_ (.A_N(net238),
    .B(net246),
    .X(_13029_));
 sky130_fd_sc_hd__mux2_1 _21186_ (.A0(_12207_),
    .A1(_13029_),
    .S(net262),
    .X(_13030_));
 sky130_fd_sc_hd__xnor2_2 _21187_ (.A(net257),
    .B(net234),
    .Y(_13031_));
 sky130_fd_sc_hd__xor2_1 _21188_ (.A(_13030_),
    .B(_13031_),
    .X(_13032_));
 sky130_fd_sc_hd__xnor2_2 _21189_ (.A(_13028_),
    .B(_13032_),
    .Y(_13033_));
 sky130_fd_sc_hd__mux2_1 _21190_ (.A0(net230),
    .A1(_12819_),
    .S(net226),
    .X(_13034_));
 sky130_fd_sc_hd__o21ai_2 _21191_ (.A1(_12924_),
    .A2(_12140_),
    .B1(_13034_),
    .Y(_13035_));
 sky130_fd_sc_hd__nand2_2 _21192_ (.A(net213),
    .B(_13035_),
    .Y(_13036_));
 sky130_fd_sc_hd__or2_1 _21193_ (.A(net213),
    .B(_13035_),
    .X(_13037_));
 sky130_fd_sc_hd__nand2_1 _21194_ (.A(_13036_),
    .B(_13037_),
    .Y(_13038_));
 sky130_fd_sc_hd__xnor2_1 _21195_ (.A(_13033_),
    .B(_13038_),
    .Y(_13039_));
 sky130_fd_sc_hd__xnor2_2 _21196_ (.A(_13027_),
    .B(_13039_),
    .Y(_13040_));
 sky130_fd_sc_hd__nor2_1 _21197_ (.A(_12180_),
    .B(_12990_),
    .Y(_13041_));
 sky130_fd_sc_hd__mux2_1 _21198_ (.A0(net213),
    .A1(_12697_),
    .S(_13041_),
    .X(_13042_));
 sky130_fd_sc_hd__xnor2_1 _21199_ (.A(_13040_),
    .B(_13042_),
    .Y(_13043_));
 sky130_fd_sc_hd__xnor2_2 _21200_ (.A(_13018_),
    .B(_13043_),
    .Y(_13044_));
 sky130_fd_sc_hd__a21oi_1 _21201_ (.A1(_12967_),
    .A2(_12996_),
    .B1(_12995_),
    .Y(_13045_));
 sky130_fd_sc_hd__a21o_1 _21202_ (.A1(_12911_),
    .A2(_12910_),
    .B1(_11759_),
    .X(_13046_));
 sky130_fd_sc_hd__or2_1 _21203_ (.A(net222),
    .B(_12910_),
    .X(_13047_));
 sky130_fd_sc_hd__a21o_1 _21204_ (.A1(_13046_),
    .A2(_13047_),
    .B1(_11789_),
    .X(_13048_));
 sky130_fd_sc_hd__nand2_1 _21205_ (.A(_13045_),
    .B(_13048_),
    .Y(_13049_));
 sky130_fd_sc_hd__nor2_1 _21206_ (.A(_13045_),
    .B(_13048_),
    .Y(_13050_));
 sky130_fd_sc_hd__inv_2 _21207_ (.A(_13050_),
    .Y(_13051_));
 sky130_fd_sc_hd__nand2_1 _21208_ (.A(_13049_),
    .B(_13051_),
    .Y(_13052_));
 sky130_fd_sc_hd__xnor2_1 _21209_ (.A(_13044_),
    .B(_13052_),
    .Y(_13053_));
 sky130_fd_sc_hd__a21o_1 _21210_ (.A1(_12531_),
    .A2(_12532_),
    .B1(_12515_),
    .X(_13054_));
 sky130_fd_sc_hd__nand3_1 _21211_ (.A(_12515_),
    .B(_12531_),
    .C(_12532_),
    .Y(_13055_));
 sky130_fd_sc_hd__nand2_1 _21212_ (.A(_12660_),
    .B(_12575_),
    .Y(_13056_));
 sky130_fd_sc_hd__a21o_1 _21213_ (.A1(_13054_),
    .A2(_13055_),
    .B1(_13056_),
    .X(_13057_));
 sky130_fd_sc_hd__or2_1 _21214_ (.A(_12660_),
    .B(_12575_),
    .X(_13058_));
 sky130_fd_sc_hd__or3_1 _21215_ (.A(_12544_),
    .B(_12545_),
    .C(_13058_),
    .X(_13059_));
 sky130_fd_sc_hd__or2_1 _21216_ (.A(_12646_),
    .B(_12577_),
    .X(_13060_));
 sky130_fd_sc_hd__nand2_1 _21217_ (.A(_12646_),
    .B(_12577_),
    .Y(_13061_));
 sky130_fd_sc_hd__a22o_1 _21218_ (.A1(_13057_),
    .A2(_13059_),
    .B1(_13060_),
    .B2(_13061_),
    .X(_13062_));
 sky130_fd_sc_hd__o211a_1 _21219_ (.A1(_12544_),
    .A2(_12545_),
    .B1(_12578_),
    .C1(_12646_),
    .X(_13063_));
 sky130_fd_sc_hd__and4b_1 _21220_ (.A_N(_12646_),
    .B(_13054_),
    .C(_13055_),
    .D(_12577_),
    .X(_13064_));
 sky130_fd_sc_hd__o211ai_1 _21221_ (.A1(_13063_),
    .A2(_13064_),
    .B1(_13056_),
    .C1(_13058_),
    .Y(_13065_));
 sky130_fd_sc_hd__inv_2 _21222_ (.A(_12620_),
    .Y(_13066_));
 sky130_fd_sc_hd__xnor2_1 _21223_ (.A(_12643_),
    .B(_12618_),
    .Y(_13067_));
 sky130_fd_sc_hd__inv_2 _21224_ (.A(_12626_),
    .Y(_13068_));
 sky130_fd_sc_hd__or3_1 _21225_ (.A(_12622_),
    .B(_13068_),
    .C(_12627_),
    .X(_13069_));
 sky130_fd_sc_hd__mux2_1 _21226_ (.A0(_12627_),
    .A1(_13068_),
    .S(_12620_),
    .X(_13070_));
 sky130_fd_sc_hd__and2_1 _21227_ (.A(_12620_),
    .B(_12627_),
    .X(_13071_));
 sky130_fd_sc_hd__mux2_1 _21228_ (.A0(_13070_),
    .A1(_13071_),
    .S(_13067_),
    .X(_13072_));
 sky130_fd_sc_hd__nand2_1 _21229_ (.A(_12622_),
    .B(_13072_),
    .Y(_13073_));
 sky130_fd_sc_hd__o31a_1 _21230_ (.A1(_13066_),
    .A2(_13067_),
    .A3(_13069_),
    .B1(_13073_),
    .X(_13074_));
 sky130_fd_sc_hd__and2_1 _21231_ (.A(_12643_),
    .B(_12618_),
    .X(_13075_));
 sky130_fd_sc_hd__xnor2_1 _21232_ (.A(_12583_),
    .B(_13075_),
    .Y(_13076_));
 sky130_fd_sc_hd__xnor2_1 _21233_ (.A(_12605_),
    .B(_13076_),
    .Y(_13077_));
 sky130_fd_sc_hd__nand2_1 _21234_ (.A(_12637_),
    .B(_13077_),
    .Y(_13078_));
 sky130_fd_sc_hd__a211o_1 _21235_ (.A1(_13062_),
    .A2(_13065_),
    .B1(_13074_),
    .C1(_13078_),
    .X(_13079_));
 sky130_fd_sc_hd__inv_2 _21236_ (.A(_12616_),
    .Y(_13080_));
 sky130_fd_sc_hd__or2b_1 _21237_ (.A(_12610_),
    .B_N(_12628_),
    .X(_13081_));
 sky130_fd_sc_hd__inv_2 _21238_ (.A(_12628_),
    .Y(_13082_));
 sky130_fd_sc_hd__a21o_1 _21239_ (.A1(_12610_),
    .A2(_13082_),
    .B1(_12642_),
    .X(_13083_));
 sky130_fd_sc_hd__a211o_1 _21240_ (.A1(_12642_),
    .A2(_13081_),
    .B1(_13080_),
    .C1(_12609_),
    .X(_13084_));
 sky130_fd_sc_hd__a32o_1 _21241_ (.A1(_12609_),
    .A2(_13080_),
    .A3(_13081_),
    .B1(_13083_),
    .B2(_13084_),
    .X(_13085_));
 sky130_fd_sc_hd__a21boi_1 _21242_ (.A1(_12583_),
    .A2(_12605_),
    .B1_N(_13085_),
    .Y(_13086_));
 sky130_fd_sc_hd__o21a_1 _21243_ (.A1(_12606_),
    .A2(_13086_),
    .B1(_12578_),
    .X(_13087_));
 sky130_fd_sc_hd__a211oi_1 _21244_ (.A1(_12660_),
    .A2(_12575_),
    .B1(_13087_),
    .C1(_12546_),
    .Y(_13088_));
 sky130_fd_sc_hd__or3_1 _21245_ (.A(_12606_),
    .B(_12578_),
    .C(_13086_),
    .X(_13089_));
 sky130_fd_sc_hd__a21oi_1 _21246_ (.A1(_13058_),
    .A2(_13089_),
    .B1(_12546_),
    .Y(_13090_));
 sky130_fd_sc_hd__or2_1 _21247_ (.A(_12533_),
    .B(_12665_),
    .X(_13091_));
 sky130_fd_sc_hd__o211ai_1 _21248_ (.A1(_13088_),
    .A2(_13090_),
    .B1(_13091_),
    .C1(_12541_),
    .Y(_13092_));
 sky130_fd_sc_hd__xnor2_1 _21249_ (.A(_12535_),
    .B(_12539_),
    .Y(_13093_));
 sky130_fd_sc_hd__a211oi_2 _21250_ (.A1(_13079_),
    .A2(_13092_),
    .B1(_13093_),
    .C1(_12666_),
    .Y(_13094_));
 sky130_fd_sc_hd__and2_1 _21251_ (.A(_12244_),
    .B(_12669_),
    .X(_13095_));
 sky130_fd_sc_hd__o2111ai_2 _21252_ (.A1(_12543_),
    .A2(_13094_),
    .B1(_13095_),
    .C1(_12738_),
    .D1(_12420_),
    .Y(_13096_));
 sky130_fd_sc_hd__a31oi_1 _21253_ (.A1(_12244_),
    .A2(_12673_),
    .A3(_12807_),
    .B1(_12736_),
    .Y(_13097_));
 sky130_fd_sc_hd__a2111o_1 _21254_ (.A1(_13096_),
    .A2(_13097_),
    .B1(_12940_),
    .C1(_12941_),
    .D1(_13008_),
    .X(_13098_));
 sky130_fd_sc_hd__nand2_1 _21255_ (.A(_12965_),
    .B(_13007_),
    .Y(_13099_));
 sky130_fd_sc_hd__a21o_1 _21256_ (.A1(_12939_),
    .A2(_12950_),
    .B1(_12938_),
    .X(_13100_));
 sky130_fd_sc_hd__nor2_1 _21257_ (.A(_12965_),
    .B(_13007_),
    .Y(_13101_));
 sky130_fd_sc_hd__a21o_1 _21258_ (.A1(_13099_),
    .A2(_13100_),
    .B1(_13101_),
    .X(_13102_));
 sky130_fd_sc_hd__and3_1 _21259_ (.A(_13053_),
    .B(_13098_),
    .C(_13102_),
    .X(_13103_));
 sky130_fd_sc_hd__a21oi_2 _21260_ (.A1(_13098_),
    .A2(_13102_),
    .B1(_13053_),
    .Y(_13104_));
 sky130_fd_sc_hd__nor2_1 _21261_ (.A(_13103_),
    .B(_13104_),
    .Y(_13105_));
 sky130_fd_sc_hd__xnor2_1 _21262_ (.A(_13016_),
    .B(_13105_),
    .Y(_13106_));
 sky130_fd_sc_hd__xnor2_2 _21263_ (.A(_13015_),
    .B(_13106_),
    .Y(_13107_));
 sky130_fd_sc_hd__nor2_1 _21264_ (.A(_12740_),
    .B(_13107_),
    .Y(_13108_));
 sky130_fd_sc_hd__a31o_1 _21265_ (.A1(net762),
    .A2(_12034_),
    .A3(_12037_),
    .B1(_13108_),
    .X(_00388_));
 sky130_fd_sc_hd__nand2_1 _21266_ (.A(_13044_),
    .B(_13051_),
    .Y(_13109_));
 sky130_fd_sc_hd__nand2_2 _21267_ (.A(_13049_),
    .B(_13109_),
    .Y(_13110_));
 sky130_fd_sc_hd__o21ba_1 _21268_ (.A1(_13027_),
    .A2(_13033_),
    .B1_N(_13038_),
    .X(_13111_));
 sky130_fd_sc_hd__a21o_2 _21269_ (.A1(_13027_),
    .A2(_13033_),
    .B1(_13111_),
    .X(_13112_));
 sky130_fd_sc_hd__nor2_1 _21270_ (.A(net239),
    .B(_13028_),
    .Y(_13113_));
 sky130_fd_sc_hd__nor2_1 _21271_ (.A(net246),
    .B(_13028_),
    .Y(_13114_));
 sky130_fd_sc_hd__o21ba_1 _21272_ (.A1(_13029_),
    .A2(_13114_),
    .B1_N(_13031_),
    .X(_13115_));
 sky130_fd_sc_hd__a221o_1 _21273_ (.A1(_12207_),
    .A2(_13031_),
    .B1(_13113_),
    .B2(net247),
    .C1(_13115_),
    .X(_13116_));
 sky130_fd_sc_hd__and2_1 _21274_ (.A(net247),
    .B(_13028_),
    .X(_13117_));
 sky130_fd_sc_hd__or2_1 _21275_ (.A(_13114_),
    .B(_13117_),
    .X(_13118_));
 sky130_fd_sc_hd__and2b_1 _21276_ (.A_N(_13031_),
    .B(_13113_),
    .X(_13119_));
 sky130_fd_sc_hd__a31o_1 _21277_ (.A1(net239),
    .A2(_13031_),
    .A3(_13118_),
    .B1(_13119_),
    .X(_13120_));
 sky130_fd_sc_hd__a21oi_2 _21278_ (.A1(net262),
    .A2(_13116_),
    .B1(_13120_),
    .Y(_13121_));
 sky130_fd_sc_hd__and2_1 _21279_ (.A(net242),
    .B(_11727_),
    .X(_13122_));
 sky130_fd_sc_hd__mux2_1 _21280_ (.A0(_12699_),
    .A1(_13122_),
    .S(net257),
    .X(_13123_));
 sky130_fd_sc_hd__xnor2_2 _21281_ (.A(net214),
    .B(_12853_),
    .Y(_13124_));
 sky130_fd_sc_hd__xnor2_2 _21282_ (.A(net251),
    .B(net229),
    .Y(_13125_));
 sky130_fd_sc_hd__xor2_1 _21283_ (.A(_13124_),
    .B(_13125_),
    .X(_13126_));
 sky130_fd_sc_hd__xnor2_2 _21284_ (.A(_13123_),
    .B(_13126_),
    .Y(_13127_));
 sky130_fd_sc_hd__nand2_1 _21285_ (.A(net248),
    .B(net242),
    .Y(_13128_));
 sky130_fd_sc_hd__a221o_1 _21286_ (.A1(_12911_),
    .A2(_13128_),
    .B1(_12761_),
    .B2(net222),
    .C1(_12826_),
    .X(_13129_));
 sky130_fd_sc_hd__nand2_2 _21287_ (.A(net213),
    .B(_13129_),
    .Y(_13130_));
 sky130_fd_sc_hd__or2_1 _21288_ (.A(net214),
    .B(_13129_),
    .X(_13131_));
 sky130_fd_sc_hd__nand2_1 _21289_ (.A(_13130_),
    .B(_13131_),
    .Y(_13132_));
 sky130_fd_sc_hd__xor2_1 _21290_ (.A(_13127_),
    .B(_13132_),
    .X(_13133_));
 sky130_fd_sc_hd__xnor2_2 _21291_ (.A(_13121_),
    .B(_13133_),
    .Y(_13134_));
 sky130_fd_sc_hd__xor2_2 _21292_ (.A(_13036_),
    .B(_13134_),
    .X(_13135_));
 sky130_fd_sc_hd__xnor2_4 _21293_ (.A(_13112_),
    .B(_13135_),
    .Y(_13136_));
 sky130_fd_sc_hd__o21ba_1 _21294_ (.A1(_13040_),
    .A2(_13042_),
    .B1_N(_13018_),
    .X(_13137_));
 sky130_fd_sc_hd__a21o_1 _21295_ (.A1(_13040_),
    .A2(_13042_),
    .B1(_13137_),
    .X(_13138_));
 sky130_fd_sc_hd__or2_1 _21296_ (.A(_13001_),
    .B(_12990_),
    .X(_13139_));
 sky130_fd_sc_hd__xnor2_2 _21297_ (.A(_13138_),
    .B(_13139_),
    .Y(_13140_));
 sky130_fd_sc_hd__xnor2_4 _21298_ (.A(_13136_),
    .B(_13140_),
    .Y(_13141_));
 sky130_fd_sc_hd__xor2_2 _21299_ (.A(_13110_),
    .B(_13141_),
    .X(_13142_));
 sky130_fd_sc_hd__nand2_1 _21300_ (.A(_13016_),
    .B(_13103_),
    .Y(_13143_));
 sky130_fd_sc_hd__inv_2 _21301_ (.A(_13143_),
    .Y(_13144_));
 sky130_fd_sc_hd__inv_2 _21302_ (.A(_13016_),
    .Y(_13145_));
 sky130_fd_sc_hd__o21bai_2 _21303_ (.A1(_13145_),
    .A2(_13104_),
    .B1_N(_13103_),
    .Y(_13146_));
 sky130_fd_sc_hd__a2bb2o_1 _21304_ (.A1_N(_13014_),
    .A2_N(_13146_),
    .B1(_13145_),
    .B2(_13104_),
    .X(_13147_));
 sky130_fd_sc_hd__mux2_1 _21305_ (.A0(_13146_),
    .A1(_13147_),
    .S(_12883_),
    .X(_13148_));
 sky130_fd_sc_hd__a21oi_1 _21306_ (.A1(_13014_),
    .A2(_13144_),
    .B1(_13148_),
    .Y(_13149_));
 sky130_fd_sc_hd__xnor2_2 _21307_ (.A(_13142_),
    .B(_13149_),
    .Y(_13150_));
 sky130_fd_sc_hd__nor2_1 _21308_ (.A(_12036_),
    .B(_13150_),
    .Y(_13151_));
 sky130_fd_sc_hd__a31o_1 _21309_ (.A1(net738),
    .A2(_12034_),
    .A3(_12037_),
    .B1(_13151_),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _21310_ (.A0(_13104_),
    .A1(_13105_),
    .S(_13145_),
    .X(_13152_));
 sky130_fd_sc_hd__mux2_1 _21311_ (.A0(_13144_),
    .A1(_13152_),
    .S(_13142_),
    .X(_13153_));
 sky130_fd_sc_hd__and2_1 _21312_ (.A(_13014_),
    .B(_13153_),
    .X(_13154_));
 sky130_fd_sc_hd__nor2_1 _21313_ (.A(net1021),
    .B(_13154_),
    .Y(_13155_));
 sky130_fd_sc_hd__a21bo_1 _21314_ (.A1(_13138_),
    .A2(_13136_),
    .B1_N(_13139_),
    .X(_13156_));
 sky130_fd_sc_hd__o21a_1 _21315_ (.A1(_13138_),
    .A2(_13136_),
    .B1(_13156_),
    .X(_13157_));
 sky130_fd_sc_hd__o21a_1 _21316_ (.A1(_13112_),
    .A2(_13134_),
    .B1(_13036_),
    .X(_13158_));
 sky130_fd_sc_hd__a21o_1 _21317_ (.A1(_13112_),
    .A2(_13134_),
    .B1(_13158_),
    .X(_13159_));
 sky130_fd_sc_hd__o21ba_1 _21318_ (.A1(_13121_),
    .A2(_13127_),
    .B1_N(_13132_),
    .X(_13160_));
 sky130_fd_sc_hd__a21o_1 _21319_ (.A1(_13121_),
    .A2(_13127_),
    .B1(_13160_),
    .X(_13161_));
 sky130_fd_sc_hd__nor2_1 _21320_ (.A(net235),
    .B(_13124_),
    .Y(_13162_));
 sky130_fd_sc_hd__nor2_1 _21321_ (.A(net242),
    .B(_13124_),
    .Y(_13163_));
 sky130_fd_sc_hd__o21ba_1 _21322_ (.A1(_13122_),
    .A2(_13163_),
    .B1_N(_13125_),
    .X(_13164_));
 sky130_fd_sc_hd__a221o_1 _21323_ (.A1(_12699_),
    .A2(_13125_),
    .B1(_13162_),
    .B2(net242),
    .C1(_13164_),
    .X(_13165_));
 sky130_fd_sc_hd__and2_1 _21324_ (.A(net242),
    .B(_13124_),
    .X(_13166_));
 sky130_fd_sc_hd__o21a_1 _21325_ (.A1(_13163_),
    .A2(_13166_),
    .B1(net235),
    .X(_13167_));
 sky130_fd_sc_hd__mux2_1 _21326_ (.A0(_13162_),
    .A1(_13167_),
    .S(_13125_),
    .X(_13168_));
 sky130_fd_sc_hd__a21oi_2 _21327_ (.A1(net257),
    .A2(_13165_),
    .B1(_13168_),
    .Y(_13169_));
 sky130_fd_sc_hd__xnor2_2 _21328_ (.A(net248),
    .B(net227),
    .Y(_13170_));
 sky130_fd_sc_hd__or2_1 _21329_ (.A(_13001_),
    .B(_13170_),
    .X(_13171_));
 sky130_fd_sc_hd__nand2_1 _21330_ (.A(_13001_),
    .B(_13170_),
    .Y(_13172_));
 sky130_fd_sc_hd__and2_1 _21331_ (.A(_13171_),
    .B(_13172_),
    .X(_13173_));
 sky130_fd_sc_hd__or2_1 _21332_ (.A(_11727_),
    .B(net231),
    .X(_13174_));
 sky130_fd_sc_hd__mux2_1 _21333_ (.A0(_12819_),
    .A1(_13174_),
    .S(\top0.cordic0.vec[0][10] ),
    .X(_13175_));
 sky130_fd_sc_hd__xnor2_1 _21334_ (.A(_13173_),
    .B(_13175_),
    .Y(_13176_));
 sky130_fd_sc_hd__a31o_1 _21335_ (.A1(net242),
    .A2(net236),
    .A3(_11759_),
    .B1(_12697_),
    .X(_13177_));
 sky130_fd_sc_hd__a22o_1 _21336_ (.A1(net213),
    .A2(_12705_),
    .B1(_13177_),
    .B2(net222),
    .X(_13178_));
 sky130_fd_sc_hd__nor2_1 _21337_ (.A(_13176_),
    .B(_13178_),
    .Y(_13179_));
 sky130_fd_sc_hd__nand2_1 _21338_ (.A(_13176_),
    .B(_13178_),
    .Y(_13180_));
 sky130_fd_sc_hd__and2b_1 _21339_ (.A_N(_13179_),
    .B(_13180_),
    .X(_13181_));
 sky130_fd_sc_hd__xnor2_2 _21340_ (.A(_13169_),
    .B(_13181_),
    .Y(_13182_));
 sky130_fd_sc_hd__xor2_1 _21341_ (.A(_13130_),
    .B(_13182_),
    .X(_13183_));
 sky130_fd_sc_hd__xnor2_2 _21342_ (.A(_13161_),
    .B(_13183_),
    .Y(_13184_));
 sky130_fd_sc_hd__nor2_1 _21343_ (.A(_11789_),
    .B(_13035_),
    .Y(_13185_));
 sky130_fd_sc_hd__xnor2_1 _21344_ (.A(_13184_),
    .B(_13185_),
    .Y(_13186_));
 sky130_fd_sc_hd__xnor2_1 _21345_ (.A(_13159_),
    .B(_13186_),
    .Y(_13187_));
 sky130_fd_sc_hd__nor2_1 _21346_ (.A(_13157_),
    .B(_13187_),
    .Y(_13188_));
 sky130_fd_sc_hd__nand2_2 _21347_ (.A(_13157_),
    .B(_13187_),
    .Y(_00916_));
 sky130_fd_sc_hd__or2b_1 _21348_ (.A(_13188_),
    .B_N(_00916_),
    .X(_00917_));
 sky130_fd_sc_hd__or2_1 _21349_ (.A(_13141_),
    .B(_13146_),
    .X(_00918_));
 sky130_fd_sc_hd__and2_1 _21350_ (.A(_13141_),
    .B(_13146_),
    .X(_00919_));
 sky130_fd_sc_hd__a21o_1 _21351_ (.A1(_13110_),
    .A2(_00918_),
    .B1(_00919_),
    .X(_00920_));
 sky130_fd_sc_hd__xnor2_1 _21352_ (.A(_00917_),
    .B(_00920_),
    .Y(_00921_));
 sky130_fd_sc_hd__xnor2_2 _21353_ (.A(_13155_),
    .B(_00921_),
    .Y(_00922_));
 sky130_fd_sc_hd__a22o_1 _21354_ (.A1(net763),
    .A2(_12813_),
    .B1(_00922_),
    .B2(_12963_),
    .X(_00390_));
 sky130_fd_sc_hd__a21o_1 _21355_ (.A1(_13141_),
    .A2(_13146_),
    .B1(_13110_),
    .X(_00923_));
 sky130_fd_sc_hd__nand2_1 _21356_ (.A(_00918_),
    .B(_00923_),
    .Y(_00924_));
 sky130_fd_sc_hd__xor2_1 _21357_ (.A(_00917_),
    .B(_00924_),
    .X(_00925_));
 sky130_fd_sc_hd__nand2_1 _21358_ (.A(_13154_),
    .B(_00925_),
    .Y(_00926_));
 sky130_fd_sc_hd__a21o_1 _21359_ (.A1(_00918_),
    .A2(_00923_),
    .B1(_13188_),
    .X(_00927_));
 sky130_fd_sc_hd__nand2_1 _21360_ (.A(_00916_),
    .B(_00927_),
    .Y(_00928_));
 sky130_fd_sc_hd__inv_2 _21361_ (.A(_13161_),
    .Y(_00929_));
 sky130_fd_sc_hd__nor2_1 _21362_ (.A(_00929_),
    .B(_13182_),
    .Y(_00930_));
 sky130_fd_sc_hd__nand2_1 _21363_ (.A(_00929_),
    .B(_13182_),
    .Y(_00931_));
 sky130_fd_sc_hd__o21ai_4 _21364_ (.A1(_13130_),
    .A2(_00930_),
    .B1(_00931_),
    .Y(_00932_));
 sky130_fd_sc_hd__o21a_1 _21365_ (.A1(_13169_),
    .A2(_13179_),
    .B1(_13180_),
    .X(_00933_));
 sky130_fd_sc_hd__xnor2_1 _21366_ (.A(_11727_),
    .B(_13001_),
    .Y(_00934_));
 sky130_fd_sc_hd__nand2_1 _21367_ (.A(net231),
    .B(_13170_),
    .Y(_00935_));
 sky130_fd_sc_hd__nor2_1 _21368_ (.A(_13001_),
    .B(_13174_),
    .Y(_00936_));
 sky130_fd_sc_hd__o21ai_1 _21369_ (.A1(net236),
    .A2(_13001_),
    .B1(_13174_),
    .Y(_00937_));
 sky130_fd_sc_hd__mux2_1 _21370_ (.A0(_00937_),
    .A1(_12820_),
    .S(_13170_),
    .X(_00938_));
 sky130_fd_sc_hd__o21ai_1 _21371_ (.A1(_00936_),
    .A2(_00938_),
    .B1(net252),
    .Y(_00939_));
 sky130_fd_sc_hd__o221a_1 _21372_ (.A1(net231),
    .A2(_13171_),
    .B1(_00934_),
    .B2(_00935_),
    .C1(_00939_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _21373_ (.A0(_12761_),
    .A1(_12981_),
    .S(net248),
    .X(_00941_));
 sky130_fd_sc_hd__xnor2_2 _21374_ (.A(net241),
    .B(net223),
    .Y(_00942_));
 sky130_fd_sc_hd__xnor2_1 _21375_ (.A(net218),
    .B(_00942_),
    .Y(_00943_));
 sky130_fd_sc_hd__xnor2_2 _21376_ (.A(_00941_),
    .B(_00943_),
    .Y(_00944_));
 sky130_fd_sc_hd__a21o_1 _21377_ (.A1(net223),
    .A2(_12815_),
    .B1(_11789_),
    .X(_00945_));
 sky130_fd_sc_hd__xor2_1 _21378_ (.A(_00944_),
    .B(_00945_),
    .X(_00946_));
 sky130_fd_sc_hd__xnor2_1 _21379_ (.A(_00940_),
    .B(_00946_),
    .Y(_00947_));
 sky130_fd_sc_hd__nor2_1 _21380_ (.A(_12705_),
    .B(_12853_),
    .Y(_00948_));
 sky130_fd_sc_hd__or2_1 _21381_ (.A(_11789_),
    .B(_00948_),
    .X(_00949_));
 sky130_fd_sc_hd__xnor2_1 _21382_ (.A(_00947_),
    .B(_00949_),
    .Y(_00950_));
 sky130_fd_sc_hd__xnor2_2 _21383_ (.A(_00933_),
    .B(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__nor2_1 _21384_ (.A(_11789_),
    .B(_13129_),
    .Y(_00952_));
 sky130_fd_sc_hd__xor2_1 _21385_ (.A(_00951_),
    .B(_00952_),
    .X(_00953_));
 sky130_fd_sc_hd__xnor2_2 _21386_ (.A(_00932_),
    .B(_00953_),
    .Y(_00954_));
 sky130_fd_sc_hd__o21ba_1 _21387_ (.A1(_13159_),
    .A2(_13184_),
    .B1_N(_13185_),
    .X(_00955_));
 sky130_fd_sc_hd__a21o_2 _21388_ (.A1(_13159_),
    .A2(_13184_),
    .B1(_00955_),
    .X(_00956_));
 sky130_fd_sc_hd__xnor2_2 _21389_ (.A(_00954_),
    .B(_00956_),
    .Y(_00957_));
 sky130_fd_sc_hd__xnor2_2 _21390_ (.A(_00928_),
    .B(_00957_),
    .Y(_00958_));
 sky130_fd_sc_hd__a21bo_1 _21391_ (.A1(_12883_),
    .A2(_00926_),
    .B1_N(_00958_),
    .X(_00959_));
 sky130_fd_sc_hd__or3b_1 _21392_ (.A(net1021),
    .B(_00958_),
    .C_N(_00926_),
    .X(_00960_));
 sky130_fd_sc_hd__a21oi_1 _21393_ (.A1(_00959_),
    .A2(_00960_),
    .B1(_12740_),
    .Y(_00961_));
 sky130_fd_sc_hd__a31o_1 _21394_ (.A1(net771),
    .A2(_12034_),
    .A3(_12037_),
    .B1(_00961_),
    .X(_00391_));
 sky130_fd_sc_hd__or2_1 _21395_ (.A(_00954_),
    .B(_00956_),
    .X(_00962_));
 sky130_fd_sc_hd__and2_1 _21396_ (.A(_00954_),
    .B(_00956_),
    .X(_00963_));
 sky130_fd_sc_hd__a31o_2 _21397_ (.A1(_00916_),
    .A2(_00927_),
    .A3(_00962_),
    .B1(_00963_),
    .X(_00964_));
 sky130_fd_sc_hd__a21o_1 _21398_ (.A1(_00932_),
    .A2(_00951_),
    .B1(_00952_),
    .X(_00965_));
 sky130_fd_sc_hd__o21ai_4 _21399_ (.A1(_00932_),
    .A2(_00951_),
    .B1(_00965_),
    .Y(_00966_));
 sky130_fd_sc_hd__o21a_1 _21400_ (.A1(_00944_),
    .A2(_00945_),
    .B1(_00940_),
    .X(_00967_));
 sky130_fd_sc_hd__a21o_1 _21401_ (.A1(_00944_),
    .A2(_00945_),
    .B1(_00967_),
    .X(_00968_));
 sky130_fd_sc_hd__nand2_1 _21402_ (.A(net232),
    .B(_11759_),
    .Y(_00969_));
 sky130_fd_sc_hd__a21oi_1 _21403_ (.A1(_00969_),
    .A2(_12764_),
    .B1(_00942_),
    .Y(_00970_));
 sky130_fd_sc_hd__a221o_1 _21404_ (.A1(net232),
    .A2(_12696_),
    .B1(_12761_),
    .B2(_00942_),
    .C1(_00970_),
    .X(_00971_));
 sky130_fd_sc_hd__and2b_1 _21405_ (.A_N(_00942_),
    .B(_12696_),
    .X(_00972_));
 sky130_fd_sc_hd__nand2_1 _21406_ (.A(_12762_),
    .B(_12764_),
    .Y(_00973_));
 sky130_fd_sc_hd__and3_1 _21407_ (.A(net228),
    .B(_00942_),
    .C(_00973_),
    .X(_00974_));
 sky130_fd_sc_hd__a211o_1 _21408_ (.A1(net248),
    .A2(_00971_),
    .B1(_00972_),
    .C1(_00974_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _21409_ (.A0(_12832_),
    .A1(_12833_),
    .S(net241),
    .X(_00976_));
 sky130_fd_sc_hd__xnor2_2 _21410_ (.A(net236),
    .B(_00976_),
    .Y(_00977_));
 sky130_fd_sc_hd__nand2_1 _21411_ (.A(net218),
    .B(_12765_),
    .Y(_00978_));
 sky130_fd_sc_hd__or2_1 _21412_ (.A(_00977_),
    .B(_00978_),
    .X(_00979_));
 sky130_fd_sc_hd__nand2_1 _21413_ (.A(_00977_),
    .B(_00978_),
    .Y(_00980_));
 sky130_fd_sc_hd__nand2_1 _21414_ (.A(_00979_),
    .B(_00980_),
    .Y(_00981_));
 sky130_fd_sc_hd__xnor2_2 _21415_ (.A(_00975_),
    .B(_00981_),
    .Y(_00982_));
 sky130_fd_sc_hd__xor2_1 _21416_ (.A(_00945_),
    .B(_00982_),
    .X(_00983_));
 sky130_fd_sc_hd__xnor2_1 _21417_ (.A(_00968_),
    .B(_00983_),
    .Y(_00984_));
 sky130_fd_sc_hd__o21ai_1 _21418_ (.A1(_00947_),
    .A2(_00948_),
    .B1(net219),
    .Y(_00985_));
 sky130_fd_sc_hd__o2bb2a_1 _21419_ (.A1_N(_00933_),
    .A2_N(_00985_),
    .B1(_00947_),
    .B2(net218),
    .X(_00986_));
 sky130_fd_sc_hd__nand2_1 _21420_ (.A(_00984_),
    .B(_00986_),
    .Y(_00987_));
 sky130_fd_sc_hd__or2_1 _21421_ (.A(_00984_),
    .B(_00986_),
    .X(_00988_));
 sky130_fd_sc_hd__nand2_1 _21422_ (.A(_00987_),
    .B(_00988_),
    .Y(_00989_));
 sky130_fd_sc_hd__xnor2_1 _21423_ (.A(_00966_),
    .B(_00989_),
    .Y(_00990_));
 sky130_fd_sc_hd__xnor2_2 _21424_ (.A(_00964_),
    .B(_00990_),
    .Y(_00991_));
 sky130_fd_sc_hd__o21a_1 _21425_ (.A1(_00958_),
    .A2(_00926_),
    .B1(_12883_),
    .X(_00992_));
 sky130_fd_sc_hd__xnor2_2 _21426_ (.A(_00991_),
    .B(_00992_),
    .Y(_00993_));
 sky130_fd_sc_hd__a22o_1 _21427_ (.A1(net785),
    .A2(_12813_),
    .B1(_00993_),
    .B2(_12963_),
    .X(_00392_));
 sky130_fd_sc_hd__and4b_2 _21428_ (.A_N(_00958_),
    .B(_00925_),
    .C(_00991_),
    .D(_13154_),
    .X(_00994_));
 sky130_fd_sc_hd__nor2_1 _21429_ (.A(_00984_),
    .B(_00986_),
    .Y(_00995_));
 sky130_fd_sc_hd__o21ai_1 _21430_ (.A1(_00966_),
    .A2(_00995_),
    .B1(_00987_),
    .Y(_00996_));
 sky130_fd_sc_hd__inv_2 _21431_ (.A(_00996_),
    .Y(_00997_));
 sky130_fd_sc_hd__a31o_1 _21432_ (.A1(_00916_),
    .A2(_00927_),
    .A3(_00956_),
    .B1(_00954_),
    .X(_00998_));
 sky130_fd_sc_hd__a21o_1 _21433_ (.A1(_00916_),
    .A2(_00927_),
    .B1(_00956_),
    .X(_00999_));
 sky130_fd_sc_hd__a21oi_1 _21434_ (.A1(_00998_),
    .A2(_00999_),
    .B1(_00987_),
    .Y(_01000_));
 sky130_fd_sc_hd__mux2_1 _21435_ (.A0(_01000_),
    .A1(_00995_),
    .S(_00966_),
    .X(_01001_));
 sky130_fd_sc_hd__a21oi_2 _21436_ (.A1(_00964_),
    .A2(_00997_),
    .B1(_01001_),
    .Y(_01002_));
 sky130_fd_sc_hd__a21o_1 _21437_ (.A1(_00967_),
    .A2(_00982_),
    .B1(_00945_),
    .X(_01003_));
 sky130_fd_sc_hd__o21a_1 _21438_ (.A1(_00968_),
    .A2(_00982_),
    .B1(_01003_),
    .X(_01004_));
 sky130_fd_sc_hd__nand2_1 _21439_ (.A(_12180_),
    .B(_12238_),
    .Y(_01005_));
 sky130_fd_sc_hd__or2_1 _21440_ (.A(net236),
    .B(net227),
    .X(_01006_));
 sky130_fd_sc_hd__a22o_1 _21441_ (.A1(net241),
    .A2(_01005_),
    .B1(_01006_),
    .B2(net223),
    .X(_01007_));
 sky130_fd_sc_hd__xor2_2 _21442_ (.A(_00973_),
    .B(_01007_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _21443_ (.A0(_00979_),
    .A1(_00980_),
    .S(_00975_),
    .X(_01009_));
 sky130_fd_sc_hd__xor2_1 _21444_ (.A(_01008_),
    .B(_01009_),
    .X(_01010_));
 sky130_fd_sc_hd__a2bb2o_1 _21445_ (.A1_N(_01004_),
    .A2_N(_01010_),
    .B1(_12815_),
    .B2(_12926_),
    .X(_01011_));
 sky130_fd_sc_hd__nand2_1 _21446_ (.A(_01004_),
    .B(_01010_),
    .Y(_01012_));
 sky130_fd_sc_hd__and2b_1 _21447_ (.A_N(_01011_),
    .B(_01012_),
    .X(_01013_));
 sky130_fd_sc_hd__xnor2_4 _21448_ (.A(_01002_),
    .B(_01013_),
    .Y(_01014_));
 sky130_fd_sc_hd__or3b_1 _21449_ (.A(net1021),
    .B(_00994_),
    .C_N(_01014_),
    .X(_01015_));
 sky130_fd_sc_hd__o21bai_1 _21450_ (.A1(net1021),
    .A2(_00994_),
    .B1_N(_01014_),
    .Y(_01016_));
 sky130_fd_sc_hd__a21oi_1 _21451_ (.A1(_01015_),
    .A2(_01016_),
    .B1(_12740_),
    .Y(_01017_));
 sky130_fd_sc_hd__a31o_1 _21452_ (.A1(net794),
    .A2(_12034_),
    .A3(_12037_),
    .B1(_01017_),
    .X(_00393_));
 sky130_fd_sc_hd__and2_1 _21453_ (.A(_00984_),
    .B(_00986_),
    .X(_01018_));
 sky130_fd_sc_hd__nor2_1 _21454_ (.A(_01018_),
    .B(_01012_),
    .Y(_01019_));
 sky130_fd_sc_hd__o2bb2a_1 _21455_ (.A1_N(_00988_),
    .A2_N(_01012_),
    .B1(_01019_),
    .B2(_00966_),
    .X(_01020_));
 sky130_fd_sc_hd__a21oi_1 _21456_ (.A1(_00996_),
    .A2(_01012_),
    .B1(_01011_),
    .Y(_01021_));
 sky130_fd_sc_hd__o21ai_2 _21457_ (.A1(_00964_),
    .A2(_01020_),
    .B1(_01021_),
    .Y(_01022_));
 sky130_fd_sc_hd__and4bb_1 _21458_ (.A_N(_00964_),
    .B_N(_00966_),
    .C(_01018_),
    .D(_01011_),
    .X(_01023_));
 sky130_fd_sc_hd__inv_2 _21459_ (.A(_01023_),
    .Y(_01024_));
 sky130_fd_sc_hd__nand2_1 _21460_ (.A(_01022_),
    .B(_01024_),
    .Y(_01025_));
 sky130_fd_sc_hd__nor2_1 _21461_ (.A(_11727_),
    .B(_12180_),
    .Y(_01026_));
 sky130_fd_sc_hd__a2bb2o_1 _21462_ (.A1_N(_01026_),
    .A2_N(_12764_),
    .B1(_12770_),
    .B2(net231),
    .X(_01027_));
 sky130_fd_sc_hd__nand2_1 _21463_ (.A(_11759_),
    .B(_01027_),
    .Y(_01028_));
 sky130_fd_sc_hd__a221o_1 _21464_ (.A1(net231),
    .A2(_12770_),
    .B1(_12814_),
    .B2(_12769_),
    .C1(_11759_),
    .X(_01029_));
 sky130_fd_sc_hd__a22o_1 _21465_ (.A1(_12769_),
    .A2(_12761_),
    .B1(_12820_),
    .B2(_11759_),
    .X(_01030_));
 sky130_fd_sc_hd__a2bb2o_1 _21466_ (.A1_N(net232),
    .A2_N(_12832_),
    .B1(_12815_),
    .B2(_12697_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _21467_ (.A0(_01030_),
    .A1(_01031_),
    .S(net241),
    .X(_01032_));
 sky130_fd_sc_hd__a21oi_1 _21468_ (.A1(_01028_),
    .A2(_01029_),
    .B1(_01032_),
    .Y(_01033_));
 sky130_fd_sc_hd__nor2_1 _21469_ (.A(_00977_),
    .B(_01008_),
    .Y(_01034_));
 sky130_fd_sc_hd__a21o_1 _21470_ (.A1(_00977_),
    .A2(_01008_),
    .B1(net218),
    .X(_01035_));
 sky130_fd_sc_hd__a2bb2o_1 _21471_ (.A1_N(_00978_),
    .A2_N(_01034_),
    .B1(_01035_),
    .B2(_00975_),
    .X(_01036_));
 sky130_fd_sc_hd__or2_1 _21472_ (.A(_01033_),
    .B(_01036_),
    .X(_01037_));
 sky130_fd_sc_hd__nand2_1 _21473_ (.A(_01033_),
    .B(_01036_),
    .Y(_01038_));
 sky130_fd_sc_hd__and3_1 _21474_ (.A(_12968_),
    .B(_01037_),
    .C(_01038_),
    .X(_01039_));
 sky130_fd_sc_hd__xor2_2 _21475_ (.A(_01025_),
    .B(_01039_),
    .X(_01040_));
 sky130_fd_sc_hd__a21oi_1 _21476_ (.A1(_01014_),
    .A2(_00994_),
    .B1(net1021),
    .Y(_01041_));
 sky130_fd_sc_hd__xnor2_1 _21477_ (.A(_01040_),
    .B(_01041_),
    .Y(_01042_));
 sky130_fd_sc_hd__and3_1 _21478_ (.A(\top0.cordic0.cos[11] ),
    .B(_12004_),
    .C(_12036_),
    .X(_01043_));
 sky130_fd_sc_hd__a21o_1 _21479_ (.A1(_12963_),
    .A2(_01042_),
    .B1(_01043_),
    .X(_00394_));
 sky130_fd_sc_hd__clkinvlp_2 _21480_ (.A(_12968_),
    .Y(_01044_));
 sky130_fd_sc_hd__o21a_1 _21481_ (.A1(net242),
    .A2(_01006_),
    .B1(net218),
    .X(_01045_));
 sky130_fd_sc_hd__nor2_1 _21482_ (.A(net231),
    .B(_01045_),
    .Y(_01046_));
 sky130_fd_sc_hd__a31o_1 _21483_ (.A1(net242),
    .A2(net236),
    .A3(net227),
    .B1(net219),
    .X(_01047_));
 sky130_fd_sc_hd__a221o_1 _21484_ (.A1(net227),
    .A2(net219),
    .B1(_01047_),
    .B2(net231),
    .C1(net223),
    .X(_01048_));
 sky130_fd_sc_hd__o31a_1 _21485_ (.A1(_12180_),
    .A2(_12824_),
    .A3(_01046_),
    .B1(_01048_),
    .X(_01049_));
 sky130_fd_sc_hd__a21o_1 _21486_ (.A1(_01022_),
    .A2(_01036_),
    .B1(_01033_),
    .X(_01050_));
 sky130_fd_sc_hd__o21a_1 _21487_ (.A1(_01022_),
    .A2(_01036_),
    .B1(_01050_),
    .X(_01051_));
 sky130_fd_sc_hd__o2111ai_1 _21488_ (.A1(_01023_),
    .A2(_01037_),
    .B1(_01038_),
    .C1(_01049_),
    .D1(_01022_),
    .Y(_01052_));
 sky130_fd_sc_hd__o31a_1 _21489_ (.A1(_01023_),
    .A2(_01049_),
    .A3(_01051_),
    .B1(_01052_),
    .X(_01053_));
 sky130_fd_sc_hd__or3b_1 _21490_ (.A(_01024_),
    .B(_01049_),
    .C_N(_01022_),
    .X(_01054_));
 sky130_fd_sc_hd__nand2_1 _21491_ (.A(_01024_),
    .B(_01049_),
    .Y(_01055_));
 sky130_fd_sc_hd__a22o_1 _21492_ (.A1(_12968_),
    .A2(_01038_),
    .B1(_01054_),
    .B2(_01055_),
    .X(_01056_));
 sky130_fd_sc_hd__o21a_1 _21493_ (.A1(_01044_),
    .A2(_01053_),
    .B1(_01056_),
    .X(_01057_));
 sky130_fd_sc_hd__a31o_1 _21494_ (.A1(_01014_),
    .A2(_00994_),
    .A3(_01040_),
    .B1(_12744_),
    .X(_01058_));
 sky130_fd_sc_hd__xnor2_1 _21495_ (.A(_01057_),
    .B(_01058_),
    .Y(_01059_));
 sky130_fd_sc_hd__a22o_1 _21496_ (.A1(net761),
    .A2(_12813_),
    .B1(_01059_),
    .B2(_12963_),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _21497_ (.A0(_01058_),
    .A1(_12883_),
    .S(_01057_),
    .X(_01060_));
 sky130_fd_sc_hd__nand3_1 _21498_ (.A(net863),
    .B(_12034_),
    .C(_12037_),
    .Y(_01061_));
 sky130_fd_sc_hd__o21ai_1 _21499_ (.A1(_12037_),
    .A2(_01060_),
    .B1(_01061_),
    .Y(_00396_));
 sky130_fd_sc_hd__inv_2 _21500_ (.A(net97),
    .Y(_01062_));
 sky130_fd_sc_hd__clkbuf_4 _21501_ (.A(_01062_),
    .X(_01063_));
 sky130_fd_sc_hd__nand2_2 _21502_ (.A(net110),
    .B(net93),
    .Y(_01064_));
 sky130_fd_sc_hd__inv_2 _21503_ (.A(net116),
    .Y(_01065_));
 sky130_fd_sc_hd__clkinv_4 _21504_ (.A(net99),
    .Y(_01066_));
 sky130_fd_sc_hd__nor2_1 _21505_ (.A(_01065_),
    .B(_01066_),
    .Y(_01067_));
 sky130_fd_sc_hd__nand2_1 _21506_ (.A(_01064_),
    .B(_01067_),
    .Y(_01068_));
 sky130_fd_sc_hd__xnor2_4 _21507_ (.A(net115),
    .B(net97),
    .Y(_01069_));
 sky130_fd_sc_hd__a21o_1 _21508_ (.A1(net124),
    .A2(net118),
    .B1(_01069_),
    .X(_01070_));
 sky130_fd_sc_hd__inv_2 _21509_ (.A(net126),
    .Y(_01071_));
 sky130_fd_sc_hd__nor2_1 _21510_ (.A(net124),
    .B(net118),
    .Y(_01072_));
 sky130_fd_sc_hd__a221o_2 _21511_ (.A1(net118),
    .A2(_01069_),
    .B1(_01070_),
    .B2(_01071_),
    .C1(_01072_),
    .X(_01073_));
 sky130_fd_sc_hd__xnor2_4 _21512_ (.A(net111),
    .B(net94),
    .Y(_01074_));
 sky130_fd_sc_hd__and2b_2 _21513_ (.A_N(net123),
    .B(net118),
    .X(_01075_));
 sky130_fd_sc_hd__xnor2_4 _21514_ (.A(net114),
    .B(_01075_),
    .Y(_01076_));
 sky130_fd_sc_hd__xnor2_2 _21515_ (.A(_01074_),
    .B(_01076_),
    .Y(_01077_));
 sky130_fd_sc_hd__nor2b_4 _21516_ (.A(net143),
    .B_N(net139),
    .Y(_01078_));
 sky130_fd_sc_hd__nor2_2 _21517_ (.A(net139),
    .B(net131),
    .Y(_01079_));
 sky130_fd_sc_hd__inv_2 _21518_ (.A(net142),
    .Y(_01080_));
 sky130_fd_sc_hd__nand2_2 _21519_ (.A(net160),
    .B(net155),
    .Y(_01081_));
 sky130_fd_sc_hd__o21a_1 _21520_ (.A1(_01080_),
    .A2(net131),
    .B1(_01081_),
    .X(_01082_));
 sky130_fd_sc_hd__a211oi_4 _21521_ (.A1(net131),
    .A2(_01078_),
    .B1(_01079_),
    .C1(_01082_),
    .Y(_01083_));
 sky130_fd_sc_hd__o21bai_1 _21522_ (.A1(_01073_),
    .A2(_01077_),
    .B1_N(_01083_),
    .Y(_01084_));
 sky130_fd_sc_hd__a21bo_1 _21523_ (.A1(_01073_),
    .A2(_01077_),
    .B1_N(_01084_),
    .X(_01085_));
 sky130_fd_sc_hd__nor3_1 _21524_ (.A(_01063_),
    .B(_01064_),
    .C(_01067_),
    .Y(_01086_));
 sky130_fd_sc_hd__a221oi_4 _21525_ (.A1(_01063_),
    .A2(_01064_),
    .B1(_01068_),
    .B2(_01085_),
    .C1(_01086_),
    .Y(_01087_));
 sky130_fd_sc_hd__xor2_4 _21526_ (.A(net159),
    .B(net139),
    .X(_01088_));
 sky130_fd_sc_hd__nor2b_2 _21527_ (.A(net132),
    .B_N(net127),
    .Y(_01089_));
 sky130_fd_sc_hd__xnor2_4 _21528_ (.A(net122),
    .B(_01089_),
    .Y(_01090_));
 sky130_fd_sc_hd__or2b_1 _21529_ (.A(net143),
    .B_N(net146),
    .X(_01091_));
 sky130_fd_sc_hd__o21ai_1 _21530_ (.A1(net146),
    .A2(_01090_),
    .B1(_01091_),
    .Y(_01092_));
 sky130_fd_sc_hd__or2b_1 _21531_ (.A(net148),
    .B_N(net141),
    .X(_01093_));
 sky130_fd_sc_hd__o22a_1 _21532_ (.A1(_01093_),
    .A2(_01088_),
    .B1(_01090_),
    .B2(_01091_),
    .X(_01094_));
 sky130_fd_sc_hd__a21bo_1 _21533_ (.A1(_01088_),
    .A2(_01092_),
    .B1_N(_01094_),
    .X(_01095_));
 sky130_fd_sc_hd__xnor2_1 _21534_ (.A(net146),
    .B(_01090_),
    .Y(_01096_));
 sky130_fd_sc_hd__a21oi_1 _21535_ (.A1(\top0.cordic0.vec[1][4] ),
    .A2(_01096_),
    .B1(_01088_),
    .Y(_01097_));
 sky130_fd_sc_hd__o21a_1 _21536_ (.A1(net143),
    .A2(_01090_),
    .B1(_01088_),
    .X(_01098_));
 sky130_fd_sc_hd__o2bb2a_2 _21537_ (.A1_N(net164),
    .A2_N(_01095_),
    .B1(_01097_),
    .B2(_01098_),
    .X(_01099_));
 sky130_fd_sc_hd__nor2b_2 _21538_ (.A(net126),
    .B_N(net123),
    .Y(_01100_));
 sky130_fd_sc_hd__xnor2_4 _21539_ (.A(net118),
    .B(_01100_),
    .Y(_01101_));
 sky130_fd_sc_hd__buf_4 _21540_ (.A(_01080_),
    .X(_01102_));
 sky130_fd_sc_hd__nor2_1 _21541_ (.A(_01102_),
    .B(net139),
    .Y(_01103_));
 sky130_fd_sc_hd__mux2_1 _21542_ (.A0(_01078_),
    .A1(_01103_),
    .S(net158),
    .X(_01104_));
 sky130_fd_sc_hd__inv_2 _21543_ (.A(net133),
    .Y(_01105_));
 sky130_fd_sc_hd__and2_1 _21544_ (.A(net155),
    .B(_01105_),
    .X(_01106_));
 sky130_fd_sc_hd__nor2_1 _21545_ (.A(net155),
    .B(_01105_),
    .Y(_01107_));
 sky130_fd_sc_hd__or2_1 _21546_ (.A(_01106_),
    .B(_01107_),
    .X(_01108_));
 sky130_fd_sc_hd__xnor2_1 _21547_ (.A(_01104_),
    .B(_01108_),
    .Y(_01109_));
 sky130_fd_sc_hd__xnor2_2 _21548_ (.A(_01101_),
    .B(_01109_),
    .Y(_01110_));
 sky130_fd_sc_hd__xor2_1 _21549_ (.A(net77),
    .B(net102),
    .X(_01111_));
 sky130_fd_sc_hd__and2b_2 _21550_ (.A_N(net115),
    .B(net109),
    .X(_01112_));
 sky130_fd_sc_hd__xnor2_4 _21551_ (.A(net104),
    .B(_01112_),
    .Y(_01113_));
 sky130_fd_sc_hd__xnor2_1 _21552_ (.A(_01111_),
    .B(_01113_),
    .Y(_01114_));
 sky130_fd_sc_hd__xnor2_4 _21553_ (.A(net105),
    .B(net86),
    .Y(_01115_));
 sky130_fd_sc_hd__nor2_1 _21554_ (.A(net114),
    .B(net109),
    .Y(_01116_));
 sky130_fd_sc_hd__a21oi_1 _21555_ (.A1(net109),
    .A2(_01115_),
    .B1(_01116_),
    .Y(_01117_));
 sky130_fd_sc_hd__xor2_2 _21556_ (.A(net105),
    .B(net86),
    .X(_01118_));
 sky130_fd_sc_hd__nand2_1 _21557_ (.A(net115),
    .B(net110),
    .Y(_01119_));
 sky130_fd_sc_hd__a21o_1 _21558_ (.A1(_01118_),
    .A2(_01119_),
    .B1(net119),
    .X(_01120_));
 sky130_fd_sc_hd__nand2_1 _21559_ (.A(_01117_),
    .B(_01120_),
    .Y(_01121_));
 sky130_fd_sc_hd__inv_2 _21560_ (.A(net122),
    .Y(_01122_));
 sky130_fd_sc_hd__and2_2 _21561_ (.A(net151),
    .B(net145),
    .X(_01123_));
 sky130_fd_sc_hd__a21oi_1 _21562_ (.A1(net132),
    .A2(_01122_),
    .B1(_01123_),
    .Y(_01124_));
 sky130_fd_sc_hd__nor2_1 _21563_ (.A(net127),
    .B(net124),
    .Y(_01125_));
 sky130_fd_sc_hd__a211oi_2 _21564_ (.A1(net124),
    .A2(_01089_),
    .B1(_01124_),
    .C1(_01125_),
    .Y(_01126_));
 sky130_fd_sc_hd__xor2_1 _21565_ (.A(_01121_),
    .B(_01126_),
    .X(_01127_));
 sky130_fd_sc_hd__xnor2_1 _21566_ (.A(_01114_),
    .B(_01127_),
    .Y(_01128_));
 sky130_fd_sc_hd__xor2_1 _21567_ (.A(_01110_),
    .B(_01128_),
    .X(_01129_));
 sky130_fd_sc_hd__xnor2_2 _21568_ (.A(_01099_),
    .B(_01129_),
    .Y(_01130_));
 sky130_fd_sc_hd__nand2_1 _21569_ (.A(net118),
    .B(net114),
    .Y(_01131_));
 sky130_fd_sc_hd__or2b_1 _21570_ (.A(_01074_),
    .B_N(_01131_),
    .X(_01132_));
 sky130_fd_sc_hd__nor2_1 _21571_ (.A(net120),
    .B(net114),
    .Y(_01133_));
 sky130_fd_sc_hd__a221o_2 _21572_ (.A1(net114),
    .A2(_01074_),
    .B1(_01132_),
    .B2(_01122_),
    .C1(_01133_),
    .X(_01134_));
 sky130_fd_sc_hd__clkbuf_4 _21573_ (.A(_01071_),
    .X(_01135_));
 sky130_fd_sc_hd__and2_2 _21574_ (.A(net154),
    .B(net149),
    .X(_01136_));
 sky130_fd_sc_hd__a21oi_1 _21575_ (.A1(net139),
    .A2(_01135_),
    .B1(_01136_),
    .Y(_01137_));
 sky130_fd_sc_hd__nor2_1 _21576_ (.A(net131),
    .B(net126),
    .Y(_01138_));
 sky130_fd_sc_hd__nand2b_2 _21577_ (.A_N(net139),
    .B(net131),
    .Y(_01139_));
 sky130_fd_sc_hd__nor2_1 _21578_ (.A(_01135_),
    .B(_01139_),
    .Y(_01140_));
 sky130_fd_sc_hd__or3_2 _21579_ (.A(_01137_),
    .B(_01138_),
    .C(_01140_),
    .X(_01141_));
 sky130_fd_sc_hd__xor2_2 _21580_ (.A(_01134_),
    .B(_01141_),
    .X(_01142_));
 sky130_fd_sc_hd__nor2b_2 _21581_ (.A(net119),
    .B_N(net116),
    .Y(_01143_));
 sky130_fd_sc_hd__xnor2_4 _21582_ (.A(net109),
    .B(_01143_),
    .Y(_01144_));
 sky130_fd_sc_hd__xnor2_2 _21583_ (.A(_01144_),
    .B(_01115_),
    .Y(_01145_));
 sky130_fd_sc_hd__xnor2_2 _21584_ (.A(_01142_),
    .B(_01145_),
    .Y(_01146_));
 sky130_fd_sc_hd__and2b_1 _21585_ (.A_N(net164),
    .B(net143),
    .X(_01147_));
 sky130_fd_sc_hd__and2b_1 _21586_ (.A_N(net143),
    .B(net164),
    .X(_01148_));
 sky130_fd_sc_hd__nor2_1 _21587_ (.A(_01147_),
    .B(_01148_),
    .Y(_01149_));
 sky130_fd_sc_hd__xnor2_2 _21588_ (.A(net149),
    .B(_01149_),
    .Y(_01150_));
 sky130_fd_sc_hd__xnor2_4 _21589_ (.A(_01071_),
    .B(_01139_),
    .Y(_01151_));
 sky130_fd_sc_hd__xnor2_2 _21590_ (.A(_01136_),
    .B(_01151_),
    .Y(_01152_));
 sky130_fd_sc_hd__and2_1 _21591_ (.A(_01150_),
    .B(_01152_),
    .X(_01153_));
 sky130_fd_sc_hd__xor2_2 _21592_ (.A(_01088_),
    .B(_01090_),
    .X(_01154_));
 sky130_fd_sc_hd__and2b_1 _21593_ (.A_N(net141),
    .B(net148),
    .X(_01155_));
 sky130_fd_sc_hd__nor2_1 _21594_ (.A(net164),
    .B(_01093_),
    .Y(_01156_));
 sky130_fd_sc_hd__a21o_1 _21595_ (.A1(net164),
    .A2(_01155_),
    .B1(_01156_),
    .X(_01157_));
 sky130_fd_sc_hd__xnor2_1 _21596_ (.A(_01154_),
    .B(_01157_),
    .Y(_01158_));
 sky130_fd_sc_hd__o21a_1 _21597_ (.A1(_01146_),
    .A2(_01153_),
    .B1(_01158_),
    .X(_01159_));
 sky130_fd_sc_hd__a21o_2 _21598_ (.A1(_01146_),
    .A2(_01153_),
    .B1(_01159_),
    .X(_01160_));
 sky130_fd_sc_hd__a21o_1 _21599_ (.A1(_01141_),
    .A2(_01145_),
    .B1(_01134_),
    .X(_01161_));
 sky130_fd_sc_hd__o21a_1 _21600_ (.A1(_01141_),
    .A2(_01145_),
    .B1(_01161_),
    .X(_01162_));
 sky130_fd_sc_hd__nand2_1 _21601_ (.A(net105),
    .B(net86),
    .Y(_01163_));
 sky130_fd_sc_hd__a21oi_1 _21602_ (.A1(net110),
    .A2(net96),
    .B1(_01163_),
    .Y(_01164_));
 sky130_fd_sc_hd__mux2_2 _21603_ (.A0(_01163_),
    .A1(_01164_),
    .S(net90),
    .X(_01165_));
 sky130_fd_sc_hd__clkinv_4 _21604_ (.A(net94),
    .Y(_01166_));
 sky130_fd_sc_hd__nor2_1 _21605_ (.A(_01063_),
    .B(_01166_),
    .Y(_01167_));
 sky130_fd_sc_hd__and3_1 _21606_ (.A(net110),
    .B(_01163_),
    .C(_01167_),
    .X(_01168_));
 sky130_fd_sc_hd__or2_1 _21607_ (.A(_01165_),
    .B(_01168_),
    .X(_01169_));
 sky130_fd_sc_hd__xnor2_1 _21608_ (.A(_01162_),
    .B(_01169_),
    .Y(_01170_));
 sky130_fd_sc_hd__xnor2_1 _21609_ (.A(_01160_),
    .B(_01170_),
    .Y(_01171_));
 sky130_fd_sc_hd__xnor2_2 _21610_ (.A(_01130_),
    .B(_01171_),
    .Y(_01172_));
 sky130_fd_sc_hd__xnor2_2 _21611_ (.A(_01073_),
    .B(_01077_),
    .Y(_01173_));
 sky130_fd_sc_hd__xnor2_4 _21612_ (.A(_01083_),
    .B(_01173_),
    .Y(_01174_));
 sky130_fd_sc_hd__xnor2_4 _21613_ (.A(net131),
    .B(_01078_),
    .Y(_01175_));
 sky130_fd_sc_hd__xnor2_1 _21614_ (.A(net158),
    .B(_01175_),
    .Y(_01176_));
 sky130_fd_sc_hd__nor2b_2 _21615_ (.A(net146),
    .B_N(net154),
    .Y(_01177_));
 sky130_fd_sc_hd__inv_2 _21616_ (.A(net146),
    .Y(_01178_));
 sky130_fd_sc_hd__or2_1 _21617_ (.A(net152),
    .B(_01178_),
    .X(_01179_));
 sky130_fd_sc_hd__o2bb2a_2 _21618_ (.A1_N(_01176_),
    .A2_N(_01177_),
    .B1(_01175_),
    .B2(_01179_),
    .X(_01180_));
 sky130_fd_sc_hd__xnor2_2 _21619_ (.A(_01150_),
    .B(_01152_),
    .Y(_01181_));
 sky130_fd_sc_hd__nand2_1 _21620_ (.A(_01180_),
    .B(_01181_),
    .Y(_01182_));
 sky130_fd_sc_hd__nor2_1 _21621_ (.A(_01180_),
    .B(_01181_),
    .Y(_01183_));
 sky130_fd_sc_hd__a21oi_2 _21622_ (.A1(_01174_),
    .A2(_01182_),
    .B1(_01183_),
    .Y(_01184_));
 sky130_fd_sc_hd__xor2_1 _21623_ (.A(net154),
    .B(_01151_),
    .X(_01185_));
 sky130_fd_sc_hd__o21bai_1 _21624_ (.A1(_01147_),
    .A2(_01185_),
    .B1_N(_01148_),
    .Y(_01186_));
 sky130_fd_sc_hd__mux2_1 _21625_ (.A0(_01148_),
    .A1(_01156_),
    .S(_01151_),
    .X(_01187_));
 sky130_fd_sc_hd__a21oi_1 _21626_ (.A1(net149),
    .A2(_01186_),
    .B1(_01187_),
    .Y(_01188_));
 sky130_fd_sc_hd__xor2_1 _21627_ (.A(_01154_),
    .B(_01146_),
    .X(_01189_));
 sky130_fd_sc_hd__xnor2_2 _21628_ (.A(_01188_),
    .B(_01189_),
    .Y(_01190_));
 sky130_fd_sc_hd__or2_1 _21629_ (.A(_01062_),
    .B(_01067_),
    .X(_01191_));
 sky130_fd_sc_hd__xor2_1 _21630_ (.A(_01064_),
    .B(_01191_),
    .X(_01192_));
 sky130_fd_sc_hd__xnor2_1 _21631_ (.A(_01085_),
    .B(_01192_),
    .Y(_01193_));
 sky130_fd_sc_hd__o21ba_1 _21632_ (.A1(_01184_),
    .A2(_01190_),
    .B1_N(_01193_),
    .X(_01194_));
 sky130_fd_sc_hd__a21o_1 _21633_ (.A1(_01184_),
    .A2(_01190_),
    .B1(_01194_),
    .X(_01195_));
 sky130_fd_sc_hd__a21bo_1 _21634_ (.A1(_01087_),
    .A2(_01172_),
    .B1_N(_01195_),
    .X(_01196_));
 sky130_fd_sc_hd__o21ai_1 _21635_ (.A1(_01087_),
    .A2(_01172_),
    .B1(_01196_),
    .Y(_01197_));
 sky130_fd_sc_hd__nor2_1 _21636_ (.A(net138),
    .B(_01101_),
    .Y(_01198_));
 sky130_fd_sc_hd__nor2_1 _21637_ (.A(_01106_),
    .B(_01107_),
    .Y(_01199_));
 sky130_fd_sc_hd__nor2_1 _21638_ (.A(net144),
    .B(_01101_),
    .Y(_01200_));
 sky130_fd_sc_hd__o21a_1 _21639_ (.A1(_01103_),
    .A2(_01200_),
    .B1(_01108_),
    .X(_01201_));
 sky130_fd_sc_hd__a221o_1 _21640_ (.A1(_01078_),
    .A2(_01199_),
    .B1(_01198_),
    .B2(net144),
    .C1(_01201_),
    .X(_01202_));
 sky130_fd_sc_hd__and2_1 _21641_ (.A(net144),
    .B(_01101_),
    .X(_01203_));
 sky130_fd_sc_hd__o211a_1 _21642_ (.A1(_01200_),
    .A2(_01203_),
    .B1(net138),
    .C1(_01199_),
    .X(_01204_));
 sky130_fd_sc_hd__a221o_4 _21643_ (.A1(_01108_),
    .A2(_01198_),
    .B1(_01202_),
    .B2(net160),
    .C1(_01204_),
    .X(_01205_));
 sky130_fd_sc_hd__nand2_1 _21644_ (.A(net138),
    .B(_01105_),
    .Y(_01206_));
 sky130_fd_sc_hd__mux2_2 _21645_ (.A0(_01139_),
    .A1(_01206_),
    .S(net155),
    .X(_01207_));
 sky130_fd_sc_hd__xnor2_4 _21646_ (.A(net150),
    .B(net128),
    .Y(_01208_));
 sky130_fd_sc_hd__xnor2_2 _21647_ (.A(_01076_),
    .B(_01208_),
    .Y(_01209_));
 sky130_fd_sc_hd__xnor2_4 _21648_ (.A(_01207_),
    .B(_01209_),
    .Y(_01210_));
 sky130_fd_sc_hd__clkinv_4 _21649_ (.A(net105),
    .Y(_01211_));
 sky130_fd_sc_hd__a21oi_1 _21650_ (.A1(net114),
    .A2(_01211_),
    .B1(_01111_),
    .Y(_01212_));
 sky130_fd_sc_hd__clkinv_4 _21651_ (.A(net109),
    .Y(_01213_));
 sky130_fd_sc_hd__mux2_1 _21652_ (.A0(_01213_),
    .A1(_01112_),
    .S(net105),
    .X(_01214_));
 sky130_fd_sc_hd__or2_1 _21653_ (.A(_01212_),
    .B(_01214_),
    .X(_01215_));
 sky130_fd_sc_hd__nand2_1 _21654_ (.A(net143),
    .B(net139),
    .Y(_01216_));
 sky130_fd_sc_hd__clkinv_4 _21655_ (.A(net121),
    .Y(_01217_));
 sky130_fd_sc_hd__nand2_1 _21656_ (.A(net126),
    .B(_01217_),
    .Y(_01218_));
 sky130_fd_sc_hd__a221o_2 _21657_ (.A1(net118),
    .A2(_01100_),
    .B1(_01216_),
    .B2(_01218_),
    .C1(_01072_),
    .X(_01219_));
 sky130_fd_sc_hd__xnor2_1 _21658_ (.A(_01215_),
    .B(_01219_),
    .Y(_01220_));
 sky130_fd_sc_hd__nand2b_2 _21659_ (.A_N(net96),
    .B(net78),
    .Y(_01221_));
 sky130_fd_sc_hd__or2b_1 _21660_ (.A(net81),
    .B_N(net96),
    .X(_01222_));
 sky130_fd_sc_hd__nand2_4 _21661_ (.A(_01221_),
    .B(_01222_),
    .Y(_01223_));
 sky130_fd_sc_hd__nand2b_4 _21662_ (.A_N(net111),
    .B(net107),
    .Y(_01224_));
 sky130_fd_sc_hd__xnor2_4 _21663_ (.A(_01066_),
    .B(_01224_),
    .Y(_01225_));
 sky130_fd_sc_hd__xor2_1 _21664_ (.A(_01223_),
    .B(_01225_),
    .X(_01226_));
 sky130_fd_sc_hd__xnor2_2 _21665_ (.A(_01220_),
    .B(_01226_),
    .Y(_01227_));
 sky130_fd_sc_hd__xnor2_2 _21666_ (.A(_01210_),
    .B(_01227_),
    .Y(_01228_));
 sky130_fd_sc_hd__xnor2_4 _21667_ (.A(_01205_),
    .B(_01228_),
    .Y(_01229_));
 sky130_fd_sc_hd__clkinv_4 _21668_ (.A(net88),
    .Y(_01230_));
 sky130_fd_sc_hd__a21o_1 _21669_ (.A1(net105),
    .A2(net90),
    .B1(_01230_),
    .X(_01231_));
 sky130_fd_sc_hd__nor2_1 _21670_ (.A(_11444_),
    .B(_01066_),
    .Y(_01232_));
 sky130_fd_sc_hd__a21o_1 _21671_ (.A1(_01117_),
    .A2(_01120_),
    .B1(_01126_),
    .X(_01233_));
 sky130_fd_sc_hd__and3_1 _21672_ (.A(_01117_),
    .B(_01120_),
    .C(_01126_),
    .X(_01234_));
 sky130_fd_sc_hd__a21o_1 _21673_ (.A1(_01114_),
    .A2(_01233_),
    .B1(_01234_),
    .X(_01235_));
 sky130_fd_sc_hd__o21a_1 _21674_ (.A1(net99),
    .A2(_01113_),
    .B1(net77),
    .X(_01236_));
 sky130_fd_sc_hd__or2_1 _21675_ (.A(_01066_),
    .B(_01113_),
    .X(_01237_));
 sky130_fd_sc_hd__nand2_1 _21676_ (.A(_01066_),
    .B(_01113_),
    .Y(_01238_));
 sky130_fd_sc_hd__and3_1 _21677_ (.A(_11444_),
    .B(_01237_),
    .C(_01238_),
    .X(_01239_));
 sky130_fd_sc_hd__o32a_1 _21678_ (.A1(_01234_),
    .A2(_01236_),
    .A3(_01239_),
    .B1(_01232_),
    .B2(_01233_),
    .X(_01240_));
 sky130_fd_sc_hd__a21bo_1 _21679_ (.A1(_01232_),
    .A2(_01235_),
    .B1_N(_01240_),
    .X(_01241_));
 sky130_fd_sc_hd__xor2_2 _21680_ (.A(_01231_),
    .B(_01241_),
    .X(_01242_));
 sky130_fd_sc_hd__and2b_1 _21681_ (.A_N(_01128_),
    .B(_01110_),
    .X(_01243_));
 sky130_fd_sc_hd__or2b_1 _21682_ (.A(_01110_),
    .B_N(_01128_),
    .X(_01244_));
 sky130_fd_sc_hd__o21ai_2 _21683_ (.A1(_01099_),
    .A2(_01243_),
    .B1(_01244_),
    .Y(_01245_));
 sky130_fd_sc_hd__xor2_2 _21684_ (.A(_01242_),
    .B(_01245_),
    .X(_01246_));
 sky130_fd_sc_hd__xnor2_4 _21685_ (.A(_01229_),
    .B(_01246_),
    .Y(_01247_));
 sky130_fd_sc_hd__nand2_2 _21686_ (.A(net96),
    .B(net90),
    .Y(_01248_));
 sky130_fd_sc_hd__or3b_2 _21687_ (.A(_01213_),
    .B(_01248_),
    .C_N(_01163_),
    .X(_01249_));
 sky130_fd_sc_hd__and2_1 _21688_ (.A(_01130_),
    .B(_01162_),
    .X(_01250_));
 sky130_fd_sc_hd__a21o_1 _21689_ (.A1(_01130_),
    .A2(_01249_),
    .B1(_01162_),
    .X(_01251_));
 sky130_fd_sc_hd__a221o_1 _21690_ (.A1(_01249_),
    .A2(_01250_),
    .B1(_01251_),
    .B2(_01165_),
    .C1(_01160_),
    .X(_01252_));
 sky130_fd_sc_hd__or2_1 _21691_ (.A(_01130_),
    .B(_01162_),
    .X(_01253_));
 sky130_fd_sc_hd__o221ai_1 _21692_ (.A1(_01165_),
    .A2(_01253_),
    .B1(_01250_),
    .B2(_01249_),
    .C1(_01160_),
    .Y(_01254_));
 sky130_fd_sc_hd__a2bb2o_1 _21693_ (.A1_N(_01249_),
    .A2_N(_01253_),
    .B1(_01250_),
    .B2(_01165_),
    .X(_01255_));
 sky130_fd_sc_hd__a21o_1 _21694_ (.A1(_01252_),
    .A2(_01254_),
    .B1(_01255_),
    .X(_01256_));
 sky130_fd_sc_hd__xnor2_1 _21695_ (.A(_01247_),
    .B(_01256_),
    .Y(_01257_));
 sky130_fd_sc_hd__or2_1 _21696_ (.A(_01197_),
    .B(_01257_),
    .X(_01258_));
 sky130_fd_sc_hd__xnor2_4 _21697_ (.A(net129),
    .B(net113),
    .Y(_01259_));
 sky130_fd_sc_hd__nand2_1 _21698_ (.A(net139),
    .B(net131),
    .Y(_01260_));
 sky130_fd_sc_hd__or2b_1 _21699_ (.A(_01259_),
    .B_N(_01260_),
    .X(_01261_));
 sky130_fd_sc_hd__a221o_4 _21700_ (.A1(net131),
    .A2(_01259_),
    .B1(_01261_),
    .B2(_01080_),
    .C1(_01079_),
    .X(_01262_));
 sky130_fd_sc_hd__xnor2_2 _21701_ (.A(net122),
    .B(net106),
    .Y(_01263_));
 sky130_fd_sc_hd__xnor2_2 _21702_ (.A(_01151_),
    .B(_01263_),
    .Y(_01264_));
 sky130_fd_sc_hd__nor2_2 _21703_ (.A(net146),
    .B(_01081_),
    .Y(_01265_));
 sky130_fd_sc_hd__inv_2 _21704_ (.A(net158),
    .Y(_01266_));
 sky130_fd_sc_hd__clkbuf_4 _21705_ (.A(_01266_),
    .X(_01267_));
 sky130_fd_sc_hd__and2b_1 _21706_ (.A_N(net152),
    .B(net146),
    .X(_01268_));
 sky130_fd_sc_hd__xnor2_2 _21707_ (.A(net152),
    .B(net146),
    .Y(_01269_));
 sky130_fd_sc_hd__mux2_1 _21708_ (.A0(_01268_),
    .A1(_01269_),
    .S(net162),
    .X(_01270_));
 sky130_fd_sc_hd__nand2_1 _21709_ (.A(net141),
    .B(_01270_),
    .Y(_01271_));
 sky130_fd_sc_hd__or3_1 _21710_ (.A(net162),
    .B(net141),
    .C(_01268_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _21711_ (.A0(_01091_),
    .A1(_01102_),
    .S(net154),
    .X(_01273_));
 sky130_fd_sc_hd__o221a_1 _21712_ (.A1(net149),
    .A2(_01149_),
    .B1(_01273_),
    .B2(net164),
    .C1(net158),
    .X(_01274_));
 sky130_fd_sc_hd__a31o_1 _21713_ (.A1(_01267_),
    .A2(_01271_),
    .A3(_01272_),
    .B1(_01274_),
    .X(_01275_));
 sky130_fd_sc_hd__nor2_1 _21714_ (.A(_01265_),
    .B(_01275_),
    .Y(_01276_));
 sky130_fd_sc_hd__o21a_1 _21715_ (.A1(_01262_),
    .A2(_01264_),
    .B1(_01276_),
    .X(_01277_));
 sky130_fd_sc_hd__and2_1 _21716_ (.A(_01262_),
    .B(_01264_),
    .X(_01278_));
 sky130_fd_sc_hd__nor2_1 _21717_ (.A(_01262_),
    .B(_01264_),
    .Y(_01279_));
 sky130_fd_sc_hd__nor2_1 _21718_ (.A(net147),
    .B(net142),
    .Y(_01280_));
 sky130_fd_sc_hd__nor2_2 _21719_ (.A(net163),
    .B(_01266_),
    .Y(_01281_));
 sky130_fd_sc_hd__mux4_1 _21720_ (.A0(_01155_),
    .A1(_01123_),
    .A2(net142),
    .A3(_01280_),
    .S0(_01266_),
    .S1(net153),
    .X(_01282_));
 sky130_fd_sc_hd__a32o_1 _21721_ (.A1(net153),
    .A2(_01280_),
    .A3(_01281_),
    .B1(_01282_),
    .B2(net167),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _21722_ (.A0(_01278_),
    .A1(_01279_),
    .S(_01283_),
    .X(_01284_));
 sky130_fd_sc_hd__nor2_1 _21723_ (.A(_01277_),
    .B(_01284_),
    .Y(_01285_));
 sky130_fd_sc_hd__nand2_2 _21724_ (.A(net122),
    .B(net106),
    .Y(_01286_));
 sky130_fd_sc_hd__nand2_2 _21725_ (.A(net129),
    .B(net1031),
    .Y(_01287_));
 sky130_fd_sc_hd__nand2_1 _21726_ (.A(net113),
    .B(_01287_),
    .Y(_01288_));
 sky130_fd_sc_hd__xor2_2 _21727_ (.A(_01286_),
    .B(_01288_),
    .X(_01289_));
 sky130_fd_sc_hd__a21o_1 _21728_ (.A1(net126),
    .A2(_01263_),
    .B1(_01138_),
    .X(_01290_));
 sky130_fd_sc_hd__nand2_1 _21729_ (.A(net131),
    .B(net126),
    .Y(_01291_));
 sky130_fd_sc_hd__xor2_2 _21730_ (.A(net123),
    .B(net108),
    .X(_01292_));
 sky130_fd_sc_hd__a21oi_2 _21731_ (.A1(_01291_),
    .A2(_01292_),
    .B1(net139),
    .Y(_01293_));
 sky130_fd_sc_hd__nand2_1 _21732_ (.A(net152),
    .B(net147),
    .Y(_01294_));
 sky130_fd_sc_hd__nor2_1 _21733_ (.A(net141),
    .B(_01294_),
    .Y(_01295_));
 sky130_fd_sc_hd__o21ai_1 _21734_ (.A1(_01290_),
    .A2(_01293_),
    .B1(_01295_),
    .Y(_01296_));
 sky130_fd_sc_hd__or3_1 _21735_ (.A(_01290_),
    .B(_01293_),
    .C(_01295_),
    .X(_01297_));
 sky130_fd_sc_hd__nand2_1 _21736_ (.A(_01296_),
    .B(_01297_),
    .Y(_01298_));
 sky130_fd_sc_hd__nand2_2 _21737_ (.A(net147),
    .B(net142),
    .Y(_01299_));
 sky130_fd_sc_hd__or2_1 _21738_ (.A(net154),
    .B(net148),
    .X(_01300_));
 sky130_fd_sc_hd__clkbuf_2 _21739_ (.A(_01300_),
    .X(_01301_));
 sky130_fd_sc_hd__a32o_1 _21740_ (.A1(_01266_),
    .A2(_01299_),
    .A3(_01301_),
    .B1(net152),
    .B2(_01102_),
    .X(_01302_));
 sky130_fd_sc_hd__or3_1 _21741_ (.A(_01266_),
    .B(_01177_),
    .C(_01155_),
    .X(_01303_));
 sky130_fd_sc_hd__o22a_1 _21742_ (.A1(net159),
    .A2(_01294_),
    .B1(_01093_),
    .B2(net157),
    .X(_01304_));
 sky130_fd_sc_hd__a21oi_1 _21743_ (.A1(_01303_),
    .A2(_01304_),
    .B1(net164),
    .Y(_01305_));
 sky130_fd_sc_hd__nor2_1 _21744_ (.A(net159),
    .B(net141),
    .Y(_01306_));
 sky130_fd_sc_hd__a2bb2o_1 _21745_ (.A1_N(net154),
    .A2_N(_01093_),
    .B1(_01136_),
    .B2(net164),
    .X(_01307_));
 sky130_fd_sc_hd__a22o_1 _21746_ (.A1(net154),
    .A2(_01306_),
    .B1(_01307_),
    .B2(net159),
    .X(_01308_));
 sky130_fd_sc_hd__a211o_1 _21747_ (.A1(net164),
    .A2(_01302_),
    .B1(_01305_),
    .C1(_01308_),
    .X(_01309_));
 sky130_fd_sc_hd__inv_2 _21748_ (.A(net136),
    .Y(_01310_));
 sky130_fd_sc_hd__clkbuf_4 _21749_ (.A(_01310_),
    .X(_01311_));
 sky130_fd_sc_hd__xnor2_4 _21750_ (.A(net119),
    .B(net102),
    .Y(_01312_));
 sky130_fd_sc_hd__xnor2_1 _21751_ (.A(_01090_),
    .B(_01312_),
    .Y(_01313_));
 sky130_fd_sc_hd__xnor2_1 _21752_ (.A(_01311_),
    .B(_01313_),
    .Y(_01314_));
 sky130_fd_sc_hd__xnor2_1 _21753_ (.A(_01309_),
    .B(_01314_),
    .Y(_01315_));
 sky130_fd_sc_hd__xnor2_2 _21754_ (.A(_01298_),
    .B(_01315_),
    .Y(_01316_));
 sky130_fd_sc_hd__xnor2_1 _21755_ (.A(_01289_),
    .B(_01316_),
    .Y(_01317_));
 sky130_fd_sc_hd__xnor2_2 _21756_ (.A(_01285_),
    .B(_01317_),
    .Y(_01318_));
 sky130_fd_sc_hd__inv_2 _21757_ (.A(net163),
    .Y(_01319_));
 sky130_fd_sc_hd__clkbuf_4 _21758_ (.A(_01319_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _21759_ (.A0(net147),
    .A1(_01177_),
    .S(net162),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _21760_ (.A0(_01177_),
    .A1(_01269_),
    .S(net162),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _21761_ (.A0(_01321_),
    .A1(_01322_),
    .S(_01266_),
    .X(_01323_));
 sky130_fd_sc_hd__a21o_1 _21762_ (.A1(_01320_),
    .A2(_01268_),
    .B1(_01323_),
    .X(_01324_));
 sky130_fd_sc_hd__nand2_1 _21763_ (.A(net166),
    .B(net158),
    .Y(_01325_));
 sky130_fd_sc_hd__nor2_1 _21764_ (.A(_01325_),
    .B(_01301_),
    .Y(_01326_));
 sky130_fd_sc_hd__xnor2_4 _21765_ (.A(net133),
    .B(net1031),
    .Y(_01327_));
 sky130_fd_sc_hd__xor2_4 _21766_ (.A(net133),
    .B(net1031),
    .X(_01328_));
 sky130_fd_sc_hd__a21oi_1 _21767_ (.A1(_01216_),
    .A2(_01328_),
    .B1(net147),
    .Y(_01329_));
 sky130_fd_sc_hd__nor2_1 _21768_ (.A(net142),
    .B(net135),
    .Y(_01330_));
 sky130_fd_sc_hd__a211o_2 _21769_ (.A1(net135),
    .A2(_01327_),
    .B1(_01329_),
    .C1(_01330_),
    .X(_01331_));
 sky130_fd_sc_hd__xnor2_4 _21770_ (.A(_01175_),
    .B(_01259_),
    .Y(_01332_));
 sky130_fd_sc_hd__xnor2_4 _21771_ (.A(_01331_),
    .B(_01332_),
    .Y(_01333_));
 sky130_fd_sc_hd__mux2_1 _21772_ (.A0(_01324_),
    .A1(_01326_),
    .S(_01333_),
    .X(_01334_));
 sky130_fd_sc_hd__inv_2 _21773_ (.A(_01334_),
    .Y(_01335_));
 sky130_fd_sc_hd__or2_1 _21774_ (.A(net152),
    .B(_01325_),
    .X(_01336_));
 sky130_fd_sc_hd__o21ai_1 _21775_ (.A1(_01331_),
    .A2(_01336_),
    .B1(_01332_),
    .Y(_01337_));
 sky130_fd_sc_hd__nor2b_4 _21776_ (.A(net147),
    .B_N(net141),
    .Y(_01338_));
 sky130_fd_sc_hd__a211o_1 _21777_ (.A1(net135),
    .A2(_01338_),
    .B1(_01330_),
    .C1(_01327_),
    .X(_01339_));
 sky130_fd_sc_hd__o211ai_2 _21778_ (.A1(net135),
    .A2(_01299_),
    .B1(_01336_),
    .C1(_01339_),
    .Y(_01340_));
 sky130_fd_sc_hd__and4_1 _21779_ (.A(net130),
    .B(net129),
    .C(net121),
    .D(net113),
    .X(_01341_));
 sky130_fd_sc_hd__nand2_1 _21780_ (.A(net129),
    .B(net113),
    .Y(_01342_));
 sky130_fd_sc_hd__and4_1 _21781_ (.A(net130),
    .B(net121),
    .C(net1031),
    .D(_01342_),
    .X(_01343_));
 sky130_fd_sc_hd__nor2_1 _21782_ (.A(net1031),
    .B(_01342_),
    .Y(_01344_));
 sky130_fd_sc_hd__and2_1 _21783_ (.A(net1031),
    .B(_01342_),
    .X(_01345_));
 sky130_fd_sc_hd__o211a_1 _21784_ (.A1(_01344_),
    .A2(_01345_),
    .B1(_01337_),
    .C1(_01340_),
    .X(_01346_));
 sky130_fd_sc_hd__a311o_1 _21785_ (.A1(_01337_),
    .A2(_01340_),
    .A3(_01341_),
    .B1(_01343_),
    .C1(_01346_),
    .X(_01347_));
 sky130_fd_sc_hd__inv_2 _21786_ (.A(_01347_),
    .Y(_01348_));
 sky130_fd_sc_hd__a21o_1 _21787_ (.A1(net132),
    .A2(net118),
    .B1(_01065_),
    .X(_01349_));
 sky130_fd_sc_hd__xor2_1 _21788_ (.A(_01342_),
    .B(_01349_),
    .X(_01350_));
 sky130_fd_sc_hd__and2_1 _21789_ (.A(_01337_),
    .B(_01340_),
    .X(_01351_));
 sky130_fd_sc_hd__xor2_1 _21790_ (.A(_01350_),
    .B(_01351_),
    .X(_01352_));
 sky130_fd_sc_hd__inv_2 _21791_ (.A(_01352_),
    .Y(_01353_));
 sky130_fd_sc_hd__xnor2_2 _21792_ (.A(_01265_),
    .B(_01264_),
    .Y(_01354_));
 sky130_fd_sc_hd__xnor2_4 _21793_ (.A(_01262_),
    .B(_01354_),
    .Y(_01355_));
 sky130_fd_sc_hd__nor2_1 _21794_ (.A(net166),
    .B(net161),
    .Y(_01356_));
 sky130_fd_sc_hd__mux2_1 _21795_ (.A0(net158),
    .A1(_01356_),
    .S(_01179_),
    .X(_01357_));
 sky130_fd_sc_hd__nor2_1 _21796_ (.A(_01266_),
    .B(net152),
    .Y(_01358_));
 sky130_fd_sc_hd__o21a_1 _21797_ (.A1(_01177_),
    .A2(_01358_),
    .B1(net162),
    .X(_01359_));
 sky130_fd_sc_hd__nor2_1 _21798_ (.A(_01357_),
    .B(_01359_),
    .Y(_01360_));
 sky130_fd_sc_hd__xnor2_2 _21799_ (.A(_01102_),
    .B(_01360_),
    .Y(_01361_));
 sky130_fd_sc_hd__xnor2_4 _21800_ (.A(_01355_),
    .B(_01361_),
    .Y(_01362_));
 sky130_fd_sc_hd__a211oi_2 _21801_ (.A1(_01335_),
    .A2(_01353_),
    .B1(_01348_),
    .C1(_01362_),
    .Y(_01363_));
 sky130_fd_sc_hd__o211a_1 _21802_ (.A1(_01335_),
    .A2(_01353_),
    .B1(_01348_),
    .C1(_01362_),
    .X(_01364_));
 sky130_fd_sc_hd__a311o_1 _21803_ (.A1(_01335_),
    .A2(_01348_),
    .A3(_01353_),
    .B1(_01363_),
    .C1(_01364_),
    .X(_01365_));
 sky130_fd_sc_hd__nand2_1 _21804_ (.A(_01318_),
    .B(_01365_),
    .Y(_01366_));
 sky130_fd_sc_hd__or3_1 _21805_ (.A(_01331_),
    .B(_01332_),
    .C(_01326_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _21806_ (.A0(net147),
    .A1(_01294_),
    .S(net162),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _21807_ (.A0(_01294_),
    .A1(_01269_),
    .S(net162),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _21808_ (.A0(_01368_),
    .A1(_01369_),
    .S(_01267_),
    .X(_01370_));
 sky130_fd_sc_hd__o221ai_1 _21809_ (.A1(_01331_),
    .A2(_01332_),
    .B1(_01301_),
    .B2(net162),
    .C1(_01370_),
    .Y(_01371_));
 sky130_fd_sc_hd__nand2b_2 _21810_ (.A_N(net155),
    .B(net160),
    .Y(_01372_));
 sky130_fd_sc_hd__o211a_1 _21811_ (.A1(net147),
    .A2(_01372_),
    .B1(_01332_),
    .C1(_01331_),
    .X(_01373_));
 sky130_fd_sc_hd__a21oi_1 _21812_ (.A1(_01367_),
    .A2(_01371_),
    .B1(_01373_),
    .Y(_01374_));
 sky130_fd_sc_hd__xnor2_1 _21813_ (.A(_01374_),
    .B(_01350_),
    .Y(_01375_));
 sky130_fd_sc_hd__xnor2_1 _21814_ (.A(_01362_),
    .B(_01375_),
    .Y(_01376_));
 sky130_fd_sc_hd__nand2_1 _21815_ (.A(net135),
    .B(net122),
    .Y(_01377_));
 sky130_fd_sc_hd__xnor2_4 _21816_ (.A(net135),
    .B(_01338_),
    .Y(_01378_));
 sky130_fd_sc_hd__xnor2_2 _21817_ (.A(_01328_),
    .B(_01378_),
    .Y(_01379_));
 sky130_fd_sc_hd__xnor2_2 _21818_ (.A(net135),
    .B(net121),
    .Y(_01380_));
 sky130_fd_sc_hd__a21oi_1 _21819_ (.A1(net142),
    .A2(_01380_),
    .B1(_01280_),
    .Y(_01381_));
 sky130_fd_sc_hd__o21bai_1 _21820_ (.A1(_01123_),
    .A2(_01380_),
    .B1_N(net152),
    .Y(_01382_));
 sky130_fd_sc_hd__and2_1 _21821_ (.A(_01381_),
    .B(_01382_),
    .X(_01383_));
 sky130_fd_sc_hd__nand2_1 _21822_ (.A(_01379_),
    .B(_01383_),
    .Y(_01384_));
 sky130_fd_sc_hd__nand2_2 _21823_ (.A(net130),
    .B(net1031),
    .Y(_01385_));
 sky130_fd_sc_hd__a22o_1 _21824_ (.A1(_01377_),
    .A2(_01384_),
    .B1(_01385_),
    .B2(_01217_),
    .X(_01386_));
 sky130_fd_sc_hd__nand2_2 _21825_ (.A(net121),
    .B(_01377_),
    .Y(_01387_));
 sky130_fd_sc_hd__a31o_1 _21826_ (.A1(_01379_),
    .A2(_01383_),
    .A3(_01387_),
    .B1(_01385_),
    .X(_01388_));
 sky130_fd_sc_hd__nor2b_1 _21827_ (.A(_01386_),
    .B_N(_01388_),
    .Y(_01389_));
 sky130_fd_sc_hd__xnor2_2 _21828_ (.A(net153),
    .B(_01281_),
    .Y(_01390_));
 sky130_fd_sc_hd__xnor2_4 _21829_ (.A(_01385_),
    .B(_01387_),
    .Y(_01391_));
 sky130_fd_sc_hd__nand2b_4 _21830_ (.A_N(net158),
    .B(net153),
    .Y(_01392_));
 sky130_fd_sc_hd__nand2_2 _21831_ (.A(_01372_),
    .B(_01392_),
    .Y(_01393_));
 sky130_fd_sc_hd__mux2_1 _21832_ (.A0(_01392_),
    .A1(_01393_),
    .S(net163),
    .X(_01394_));
 sky130_fd_sc_hd__xnor2_2 _21833_ (.A(_01178_),
    .B(_01394_),
    .Y(_01395_));
 sky130_fd_sc_hd__xnor2_4 _21834_ (.A(_01333_),
    .B(_01395_),
    .Y(_01396_));
 sky130_fd_sc_hd__o21ai_2 _21835_ (.A1(_01390_),
    .A2(_01391_),
    .B1(_01396_),
    .Y(_01397_));
 sky130_fd_sc_hd__xnor2_2 _21836_ (.A(_01327_),
    .B(_01378_),
    .Y(_01398_));
 sky130_fd_sc_hd__nand2_2 _21837_ (.A(_01381_),
    .B(_01382_),
    .Y(_01399_));
 sky130_fd_sc_hd__o211a_1 _21838_ (.A1(_01398_),
    .A2(_01399_),
    .B1(_01390_),
    .C1(_01391_),
    .X(_01400_));
 sky130_fd_sc_hd__o21bai_2 _21839_ (.A1(_01384_),
    .A2(_01391_),
    .B1_N(_01400_),
    .Y(_01401_));
 sky130_fd_sc_hd__and3_1 _21840_ (.A(_01398_),
    .B(_01399_),
    .C(_01391_),
    .X(_01402_));
 sky130_fd_sc_hd__a311oi_4 _21841_ (.A1(_01398_),
    .A2(_01399_),
    .A3(_01396_),
    .B1(_01401_),
    .C1(_01402_),
    .Y(_01403_));
 sky130_fd_sc_hd__nand3_1 _21842_ (.A(_01389_),
    .B(_01397_),
    .C(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hd__a21oi_1 _21843_ (.A1(_01397_),
    .A2(_01403_),
    .B1(_01389_),
    .Y(_01405_));
 sky130_fd_sc_hd__a21o_1 _21844_ (.A1(_01376_),
    .A2(_01404_),
    .B1(_01405_),
    .X(_01406_));
 sky130_fd_sc_hd__o21ba_1 _21845_ (.A1(_01318_),
    .A2(_01365_),
    .B1_N(_01406_),
    .X(_01407_));
 sky130_fd_sc_hd__clkbuf_4 _21846_ (.A(_01122_),
    .X(_01408_));
 sky130_fd_sc_hd__nand2_1 _21847_ (.A(net135),
    .B(net121),
    .Y(_01409_));
 sky130_fd_sc_hd__and2b_1 _21848_ (.A_N(net122),
    .B(net141),
    .X(_01410_));
 sky130_fd_sc_hd__and2b_1 _21849_ (.A_N(net141),
    .B(net122),
    .X(_01411_));
 sky130_fd_sc_hd__buf_4 _21850_ (.A(_01380_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _21851_ (.A0(_01410_),
    .A1(_01411_),
    .S(_01412_),
    .X(_01413_));
 sky130_fd_sc_hd__xnor2_1 _21852_ (.A(net141),
    .B(_01412_),
    .Y(_01414_));
 sky130_fd_sc_hd__mux2_1 _21853_ (.A0(_01411_),
    .A1(_01410_),
    .S(_01380_),
    .X(_01415_));
 sky130_fd_sc_hd__o21a_1 _21854_ (.A1(net158),
    .A2(_01178_),
    .B1(_01415_),
    .X(_01416_));
 sky130_fd_sc_hd__a31o_1 _21855_ (.A1(net158),
    .A2(_01178_),
    .A3(_01414_),
    .B1(_01416_),
    .X(_01417_));
 sky130_fd_sc_hd__a22o_2 _21856_ (.A1(_01268_),
    .A2(_01413_),
    .B1(_01417_),
    .B2(net152),
    .X(_01418_));
 sky130_fd_sc_hd__o21ai_1 _21857_ (.A1(_01408_),
    .A2(_01409_),
    .B1(_01418_),
    .Y(_01419_));
 sky130_fd_sc_hd__nand2_1 _21858_ (.A(net145),
    .B(net129),
    .Y(_01420_));
 sky130_fd_sc_hd__nor2_1 _21859_ (.A(_01418_),
    .B(_01409_),
    .Y(_01421_));
 sky130_fd_sc_hd__a221o_1 _21860_ (.A1(_01408_),
    .A2(_01409_),
    .B1(_01419_),
    .B2(_01420_),
    .C1(_01421_),
    .X(_01422_));
 sky130_fd_sc_hd__nor2_1 _21861_ (.A(_01399_),
    .B(_01390_),
    .Y(_01423_));
 sky130_fd_sc_hd__nand2_1 _21862_ (.A(_01399_),
    .B(_01390_),
    .Y(_01424_));
 sky130_fd_sc_hd__o21ai_1 _21863_ (.A1(_01379_),
    .A2(_01423_),
    .B1(_01424_),
    .Y(_01425_));
 sky130_fd_sc_hd__xnor2_1 _21864_ (.A(_01391_),
    .B(_01425_),
    .Y(_01426_));
 sky130_fd_sc_hd__xnor2_1 _21865_ (.A(_01396_),
    .B(_01426_),
    .Y(_01427_));
 sky130_fd_sc_hd__nor2_1 _21866_ (.A(_01422_),
    .B(_01427_),
    .Y(_01428_));
 sky130_fd_sc_hd__and2_1 _21867_ (.A(_01422_),
    .B(_01427_),
    .X(_01429_));
 sky130_fd_sc_hd__a21o_1 _21868_ (.A1(net145),
    .A2(net129),
    .B1(_01122_),
    .X(_01430_));
 sky130_fd_sc_hd__xor2_1 _21869_ (.A(_01409_),
    .B(_01430_),
    .X(_01431_));
 sky130_fd_sc_hd__xnor2_2 _21870_ (.A(_01418_),
    .B(_01431_),
    .Y(_01432_));
 sky130_fd_sc_hd__or2_1 _21871_ (.A(_01399_),
    .B(_01390_),
    .X(_01433_));
 sky130_fd_sc_hd__and2_1 _21872_ (.A(_01424_),
    .B(_01433_),
    .X(_01434_));
 sky130_fd_sc_hd__xnor2_2 _21873_ (.A(_01379_),
    .B(_01434_),
    .Y(_01435_));
 sky130_fd_sc_hd__a21o_1 _21874_ (.A1(net151),
    .A2(_01122_),
    .B1(_01338_),
    .X(_01436_));
 sky130_fd_sc_hd__xnor2_1 _21875_ (.A(_01412_),
    .B(_01436_),
    .Y(_01437_));
 sky130_fd_sc_hd__o21ai_1 _21876_ (.A1(net151),
    .A2(_01122_),
    .B1(_01299_),
    .Y(_01438_));
 sky130_fd_sc_hd__xor2_1 _21877_ (.A(_01412_),
    .B(_01438_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _21878_ (.A0(_01437_),
    .A1(_01439_),
    .S(net166),
    .X(_01440_));
 sky130_fd_sc_hd__or2b_1 _21879_ (.A(net161),
    .B_N(net166),
    .X(_01441_));
 sky130_fd_sc_hd__inv_2 _21880_ (.A(_01441_),
    .Y(_01442_));
 sky130_fd_sc_hd__o22ai_1 _21881_ (.A1(_01281_),
    .A2(_01442_),
    .B1(_01437_),
    .B2(net156),
    .Y(_01443_));
 sky130_fd_sc_hd__a21o_1 _21882_ (.A1(net156),
    .A2(_01440_),
    .B1(_01443_),
    .X(_01444_));
 sky130_fd_sc_hd__o21a_1 _21883_ (.A1(_01432_),
    .A2(_01435_),
    .B1(_01444_),
    .X(_01445_));
 sky130_fd_sc_hd__a21oi_1 _21884_ (.A1(_01432_),
    .A2(_01435_),
    .B1(_01445_),
    .Y(_01446_));
 sky130_fd_sc_hd__and2b_1 _21885_ (.A_N(_01429_),
    .B(_01446_),
    .X(_01447_));
 sky130_fd_sc_hd__nand2_1 _21886_ (.A(_01397_),
    .B(_01403_),
    .Y(_01448_));
 sky130_fd_sc_hd__xnor2_1 _21887_ (.A(_01376_),
    .B(_01389_),
    .Y(_01449_));
 sky130_fd_sc_hd__xnor2_1 _21888_ (.A(_01448_),
    .B(_01449_),
    .Y(_01450_));
 sky130_fd_sc_hd__o21a_1 _21889_ (.A1(_01428_),
    .A2(_01447_),
    .B1(_01450_),
    .X(_01451_));
 sky130_fd_sc_hd__a21oi_1 _21890_ (.A1(_01366_),
    .A2(_01407_),
    .B1(_01451_),
    .Y(_01452_));
 sky130_fd_sc_hd__xnor2_1 _21891_ (.A(_01444_),
    .B(_01435_),
    .Y(_01453_));
 sky130_fd_sc_hd__xnor2_1 _21892_ (.A(_01432_),
    .B(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__xor2_4 _21893_ (.A(net148),
    .B(_01392_),
    .X(_01455_));
 sky130_fd_sc_hd__nor2_4 _21894_ (.A(_01411_),
    .B(_01410_),
    .Y(_01456_));
 sky130_fd_sc_hd__xnor2_2 _21895_ (.A(_01455_),
    .B(_01456_),
    .Y(_01457_));
 sky130_fd_sc_hd__xor2_2 _21896_ (.A(net150),
    .B(net128),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _21897_ (.A0(net160),
    .A1(_01458_),
    .S(net155),
    .X(_01459_));
 sky130_fd_sc_hd__a21o_1 _21898_ (.A1(_01081_),
    .A2(_01458_),
    .B1(net167),
    .X(_01460_));
 sky130_fd_sc_hd__nand2_1 _21899_ (.A(_01459_),
    .B(_01460_),
    .Y(_01461_));
 sky130_fd_sc_hd__nor2_1 _21900_ (.A(_01457_),
    .B(_01461_),
    .Y(_01462_));
 sky130_fd_sc_hd__a21o_1 _21901_ (.A1(net151),
    .A2(net130),
    .B1(_01135_),
    .X(_01463_));
 sky130_fd_sc_hd__nand2_2 _21902_ (.A(net145),
    .B(net122),
    .Y(_01464_));
 sky130_fd_sc_hd__a21o_1 _21903_ (.A1(_01462_),
    .A2(_01463_),
    .B1(_01464_),
    .X(_01465_));
 sky130_fd_sc_hd__a21o_1 _21904_ (.A1(net151),
    .A2(net130),
    .B1(_01462_),
    .X(_01466_));
 sky130_fd_sc_hd__nand2_1 _21905_ (.A(_01135_),
    .B(_01464_),
    .Y(_01467_));
 sky130_fd_sc_hd__and3_1 _21906_ (.A(_01465_),
    .B(_01466_),
    .C(_01467_),
    .X(_01468_));
 sky130_fd_sc_hd__nand2_1 _21907_ (.A(_01358_),
    .B(_01436_),
    .Y(_01469_));
 sky130_fd_sc_hd__o221a_1 _21908_ (.A1(_01393_),
    .A2(_01436_),
    .B1(_01438_),
    .B2(_01392_),
    .C1(_01469_),
    .X(_01470_));
 sky130_fd_sc_hd__xnor2_2 _21909_ (.A(_01412_),
    .B(_01470_),
    .Y(_01471_));
 sky130_fd_sc_hd__xor2_2 _21910_ (.A(_01464_),
    .B(_01463_),
    .X(_01472_));
 sky130_fd_sc_hd__inv_2 _21911_ (.A(_01472_),
    .Y(_01473_));
 sky130_fd_sc_hd__inv_2 _21912_ (.A(_01462_),
    .Y(_01474_));
 sky130_fd_sc_hd__nand2_1 _21913_ (.A(_01457_),
    .B(_01461_),
    .Y(_01475_));
 sky130_fd_sc_hd__o21a_1 _21914_ (.A1(net166),
    .A2(_01462_),
    .B1(_01475_),
    .X(_01476_));
 sky130_fd_sc_hd__a21bo_1 _21915_ (.A1(_01472_),
    .A2(_01475_),
    .B1_N(_01471_),
    .X(_01477_));
 sky130_fd_sc_hd__o22a_1 _21916_ (.A1(_01472_),
    .A2(_01476_),
    .B1(_01477_),
    .B2(_01320_),
    .X(_01478_));
 sky130_fd_sc_hd__o221a_1 _21917_ (.A1(net166),
    .A2(_01471_),
    .B1(_01473_),
    .B2(_01474_),
    .C1(_01478_),
    .X(_01479_));
 sky130_fd_sc_hd__nor2_1 _21918_ (.A(_01468_),
    .B(_01479_),
    .Y(_01480_));
 sky130_fd_sc_hd__a21oi_1 _21919_ (.A1(_01458_),
    .A2(_01393_),
    .B1(net165),
    .Y(_01481_));
 sky130_fd_sc_hd__a21oi_1 _21920_ (.A1(net165),
    .A2(_01459_),
    .B1(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__xnor2_2 _21921_ (.A(_01457_),
    .B(_01482_),
    .Y(_01483_));
 sky130_fd_sc_hd__mux2_1 _21922_ (.A0(_01106_),
    .A1(_01107_),
    .S(_01208_),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _21923_ (.A0(_01106_),
    .A1(_01107_),
    .S(_01458_),
    .X(_01485_));
 sky130_fd_sc_hd__a22o_1 _21924_ (.A1(_01281_),
    .A2(_01484_),
    .B1(_01485_),
    .B2(_01442_),
    .X(_01486_));
 sky130_fd_sc_hd__nand2_1 _21925_ (.A(net156),
    .B(net137),
    .Y(_01487_));
 sky130_fd_sc_hd__nand2_1 _21926_ (.A(net151),
    .B(net129),
    .Y(_01488_));
 sky130_fd_sc_hd__a21oi_1 _21927_ (.A1(\top0.cordic0.vec[1][6] ),
    .A2(_01487_),
    .B1(_01488_),
    .Y(_01489_));
 sky130_fd_sc_hd__and3_1 _21928_ (.A(net130),
    .B(_01487_),
    .C(_01488_),
    .X(_01490_));
 sky130_fd_sc_hd__or2_1 _21929_ (.A(_01489_),
    .B(_01490_),
    .X(_01491_));
 sky130_fd_sc_hd__xor2_1 _21930_ (.A(_01486_),
    .B(_01491_),
    .X(_01492_));
 sky130_fd_sc_hd__xnor2_1 _21931_ (.A(_01483_),
    .B(_01492_),
    .Y(_01493_));
 sky130_fd_sc_hd__nand2_1 _21932_ (.A(net151),
    .B(net137),
    .Y(_01494_));
 sky130_fd_sc_hd__a21oi_1 _21933_ (.A1(net163),
    .A2(_01123_),
    .B1(_01280_),
    .Y(_01495_));
 sky130_fd_sc_hd__and2b_1 _21934_ (.A_N(net136),
    .B(net153),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _21935_ (.A0(net136),
    .A1(_01496_),
    .S(_01267_),
    .X(_01497_));
 sky130_fd_sc_hd__nand2_1 _21936_ (.A(_01267_),
    .B(_01330_),
    .Y(_01498_));
 sky130_fd_sc_hd__o31a_1 _21937_ (.A1(_01267_),
    .A2(net147),
    .A3(_01216_),
    .B1(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__o22a_1 _21938_ (.A1(_01495_),
    .A2(_01497_),
    .B1(_01499_),
    .B2(net162),
    .X(_01500_));
 sky130_fd_sc_hd__a21o_1 _21939_ (.A1(_01102_),
    .A2(_01301_),
    .B1(_01136_),
    .X(_01501_));
 sky130_fd_sc_hd__a21o_1 _21940_ (.A1(net164),
    .A2(_01501_),
    .B1(_01295_),
    .X(_01502_));
 sky130_fd_sc_hd__o31a_1 _21941_ (.A1(net159),
    .A2(net136),
    .A3(_01136_),
    .B1(_01301_),
    .X(_01503_));
 sky130_fd_sc_hd__o21ai_1 _21942_ (.A1(net151),
    .A2(net136),
    .B1(net165),
    .Y(_01504_));
 sky130_fd_sc_hd__or2_1 _21943_ (.A(_01320_),
    .B(net154),
    .X(_01505_));
 sky130_fd_sc_hd__a21o_1 _21944_ (.A1(_01311_),
    .A2(_01505_),
    .B1(_01267_),
    .X(_01506_));
 sky130_fd_sc_hd__o2111a_1 _21945_ (.A1(net165),
    .A2(_01503_),
    .B1(_01504_),
    .C1(net145),
    .D1(_01506_),
    .X(_01507_));
 sky130_fd_sc_hd__a21oi_1 _21946_ (.A1(net165),
    .A2(net137),
    .B1(_01356_),
    .Y(_01508_));
 sky130_fd_sc_hd__xnor2_1 _21947_ (.A(_01199_),
    .B(_01508_),
    .Y(_01509_));
 sky130_fd_sc_hd__a311o_1 _21948_ (.A1(net160),
    .A2(net137),
    .A3(_01502_),
    .B1(_01507_),
    .C1(_01509_),
    .X(_01510_));
 sky130_fd_sc_hd__o311a_1 _21949_ (.A1(net156),
    .A2(_01441_),
    .A3(_01494_),
    .B1(_01500_),
    .C1(_01510_),
    .X(_01511_));
 sky130_fd_sc_hd__nand2_1 _21950_ (.A(net161),
    .B(net137),
    .Y(_01512_));
 sky130_fd_sc_hd__and3_1 _21951_ (.A(net166),
    .B(_01123_),
    .C(_01512_),
    .X(_01513_));
 sky130_fd_sc_hd__nor2_1 _21952_ (.A(_01511_),
    .B(_01513_),
    .Y(_01514_));
 sky130_fd_sc_hd__nand2_1 _21953_ (.A(net156),
    .B(net130),
    .Y(_01515_));
 sky130_fd_sc_hd__or3b_1 _21954_ (.A(_01267_),
    .B(_01102_),
    .C_N(_01515_),
    .X(_01516_));
 sky130_fd_sc_hd__nor2_1 _21955_ (.A(net156),
    .B(net130),
    .Y(_01517_));
 sky130_fd_sc_hd__nand2_1 _21956_ (.A(_01442_),
    .B(_01517_),
    .Y(_01518_));
 sky130_fd_sc_hd__a21o_1 _21957_ (.A1(_01516_),
    .A2(_01518_),
    .B1(_01311_),
    .X(_01519_));
 sky130_fd_sc_hd__a21oi_1 _21958_ (.A1(net161),
    .A2(_01102_),
    .B1(_01356_),
    .Y(_01520_));
 sky130_fd_sc_hd__o211a_1 _21959_ (.A1(_01515_),
    .A2(_01520_),
    .B1(_01516_),
    .C1(net137),
    .X(_01521_));
 sky130_fd_sc_hd__a211oi_1 _21960_ (.A1(_01325_),
    .A2(_01515_),
    .B1(_01517_),
    .C1(net137),
    .Y(_01522_));
 sky130_fd_sc_hd__o21a_1 _21961_ (.A1(_01521_),
    .A2(_01522_),
    .B1(_01518_),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _21962_ (.A0(net155),
    .A1(_01105_),
    .S(net160),
    .X(_01524_));
 sky130_fd_sc_hd__o211a_1 _21963_ (.A1(net160),
    .A2(net130),
    .B1(_01372_),
    .C1(net165),
    .X(_01525_));
 sky130_fd_sc_hd__a21o_1 _21964_ (.A1(_01320_),
    .A2(_01524_),
    .B1(_01525_),
    .X(_01526_));
 sky130_fd_sc_hd__xnor2_1 _21965_ (.A(_01208_),
    .B(_01526_),
    .Y(_01527_));
 sky130_fd_sc_hd__nand2_1 _21966_ (.A(_01523_),
    .B(_01527_),
    .Y(_01528_));
 sky130_fd_sc_hd__o211a_1 _21967_ (.A1(_01493_),
    .A2(_01514_),
    .B1(_01519_),
    .C1(_01528_),
    .X(_01529_));
 sky130_fd_sc_hd__nor2_1 _21968_ (.A(_01523_),
    .B(_01527_),
    .Y(_01530_));
 sky130_fd_sc_hd__nand2_1 _21969_ (.A(_01511_),
    .B(_01513_),
    .Y(_01531_));
 sky130_fd_sc_hd__or2_1 _21970_ (.A(_01523_),
    .B(_01527_),
    .X(_01532_));
 sky130_fd_sc_hd__nand2_1 _21971_ (.A(_01528_),
    .B(_01532_),
    .Y(_01533_));
 sky130_fd_sc_hd__mux2_1 _21972_ (.A0(_01474_),
    .A1(_01475_),
    .S(net166),
    .X(_01534_));
 sky130_fd_sc_hd__xnor2_1 _21973_ (.A(_01471_),
    .B(_01472_),
    .Y(_01535_));
 sky130_fd_sc_hd__xnor2_1 _21974_ (.A(_01534_),
    .B(_01535_),
    .Y(_01536_));
 sky130_fd_sc_hd__a221o_1 _21975_ (.A1(net130),
    .A2(_01488_),
    .B1(_01486_),
    .B2(_01483_),
    .C1(_01489_),
    .X(_01537_));
 sky130_fd_sc_hd__a311o_1 _21976_ (.A1(net156),
    .A2(net137),
    .A3(_01488_),
    .B1(_01486_),
    .C1(_01483_),
    .X(_01538_));
 sky130_fd_sc_hd__nand2_1 _21977_ (.A(_01537_),
    .B(_01538_),
    .Y(_01539_));
 sky130_fd_sc_hd__a32o_1 _21978_ (.A1(_01493_),
    .A2(_01531_),
    .A3(_01533_),
    .B1(_01536_),
    .B2(_01539_),
    .X(_01540_));
 sky130_fd_sc_hd__a221o_1 _21979_ (.A1(_01493_),
    .A2(_01514_),
    .B1(_01519_),
    .B2(_01530_),
    .C1(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__o2bb2a_1 _21980_ (.A1_N(_01468_),
    .A2_N(_01479_),
    .B1(_01539_),
    .B2(_01536_),
    .X(_01542_));
 sky130_fd_sc_hd__o221a_1 _21981_ (.A1(_01454_),
    .A2(_01480_),
    .B1(_01529_),
    .B2(_01541_),
    .C1(_01542_),
    .X(_01543_));
 sky130_fd_sc_hd__nor2_1 _21982_ (.A(_01428_),
    .B(_01429_),
    .Y(_01544_));
 sky130_fd_sc_hd__mux2_1 _21983_ (.A0(_01544_),
    .A1(_01429_),
    .S(_01446_),
    .X(_01545_));
 sky130_fd_sc_hd__a22oi_1 _21984_ (.A1(_01446_),
    .A2(_01428_),
    .B1(_01545_),
    .B2(_01450_),
    .Y(_01546_));
 sky130_fd_sc_hd__a211o_1 _21985_ (.A1(_01454_),
    .A2(_01480_),
    .B1(_01543_),
    .C1(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__nand2_1 _21986_ (.A(net147),
    .B(_01311_),
    .Y(_01548_));
 sky130_fd_sc_hd__a221o_2 _21987_ (.A1(net135),
    .A2(_01338_),
    .B1(_01325_),
    .B2(_01548_),
    .C1(_01330_),
    .X(_01549_));
 sky130_fd_sc_hd__nand2_1 _21988_ (.A(net127),
    .B(net124),
    .Y(_01550_));
 sky130_fd_sc_hd__or2b_1 _21989_ (.A(_01312_),
    .B_N(_01550_),
    .X(_01551_));
 sky130_fd_sc_hd__a221o_1 _21990_ (.A1(net124),
    .A2(_01312_),
    .B1(_01551_),
    .B2(_01105_),
    .C1(_01125_),
    .X(_01552_));
 sky130_fd_sc_hd__xnor2_2 _21991_ (.A(_01069_),
    .B(_01101_),
    .Y(_01553_));
 sky130_fd_sc_hd__xor2_1 _21992_ (.A(_01552_),
    .B(_01553_),
    .X(_01554_));
 sky130_fd_sc_hd__xnor2_2 _21993_ (.A(_01549_),
    .B(_01554_),
    .Y(_01555_));
 sky130_fd_sc_hd__xnor2_1 _21994_ (.A(_01319_),
    .B(_01378_),
    .Y(_01556_));
 sky130_fd_sc_hd__o22a_2 _21995_ (.A1(_01378_),
    .A2(_01392_),
    .B1(_01556_),
    .B2(_01372_),
    .X(_01557_));
 sky130_fd_sc_hd__xnor2_4 _21996_ (.A(_01175_),
    .B(_01455_),
    .Y(_01558_));
 sky130_fd_sc_hd__xnor2_1 _21997_ (.A(_01557_),
    .B(_01558_),
    .Y(_01559_));
 sky130_fd_sc_hd__xnor2_2 _21998_ (.A(_01555_),
    .B(_01559_),
    .Y(_01560_));
 sky130_fd_sc_hd__or3b_1 _21999_ (.A(_01290_),
    .B(_01293_),
    .C_N(_01295_),
    .X(_01561_));
 sky130_fd_sc_hd__o21ba_1 _22000_ (.A1(_01290_),
    .A2(_01293_),
    .B1_N(_01295_),
    .X(_01562_));
 sky130_fd_sc_hd__a21o_1 _22001_ (.A1(_01313_),
    .A2(_01561_),
    .B1(_01562_),
    .X(_01563_));
 sky130_fd_sc_hd__nand2_1 _22002_ (.A(net118),
    .B(net102),
    .Y(_01564_));
 sky130_fd_sc_hd__nand2_1 _22003_ (.A(net124),
    .B(net109),
    .Y(_01565_));
 sky130_fd_sc_hd__nand2_1 _22004_ (.A(net106),
    .B(_01565_),
    .Y(_01566_));
 sky130_fd_sc_hd__xnor2_1 _22005_ (.A(_01564_),
    .B(_01566_),
    .Y(_01567_));
 sky130_fd_sc_hd__xnor2_1 _22006_ (.A(_01563_),
    .B(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__a2bb2o_1 _22007_ (.A1_N(net166),
    .A2_N(_01512_),
    .B1(_01311_),
    .B2(_01442_),
    .X(_01569_));
 sky130_fd_sc_hd__or3_1 _22008_ (.A(_01319_),
    .B(net158),
    .C(_01310_),
    .X(_01570_));
 sky130_fd_sc_hd__or3_1 _22009_ (.A(net163),
    .B(_01266_),
    .C(net136),
    .X(_01571_));
 sky130_fd_sc_hd__nand2_1 _22010_ (.A(_01570_),
    .B(_01571_),
    .Y(_01572_));
 sky130_fd_sc_hd__mux2_1 _22011_ (.A0(_01155_),
    .A1(_01338_),
    .S(net153),
    .X(_01573_));
 sky130_fd_sc_hd__a32o_1 _22012_ (.A1(net142),
    .A2(_01269_),
    .A3(_01569_),
    .B1(_01572_),
    .B2(_01573_),
    .X(_01574_));
 sky130_fd_sc_hd__xor2_1 _22013_ (.A(_01090_),
    .B(_01312_),
    .X(_01575_));
 sky130_fd_sc_hd__and3_1 _22014_ (.A(_01296_),
    .B(_01297_),
    .C(_01575_),
    .X(_01576_));
 sky130_fd_sc_hd__a21oi_1 _22015_ (.A1(_01296_),
    .A2(_01297_),
    .B1(_01575_),
    .Y(_01577_));
 sky130_fd_sc_hd__mux2_1 _22016_ (.A0(net136),
    .A1(_01512_),
    .S(_01319_),
    .X(_01578_));
 sky130_fd_sc_hd__xor2_1 _22017_ (.A(net153),
    .B(net135),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _22018_ (.A0(net151),
    .A1(_01338_),
    .S(_01579_),
    .X(_01580_));
 sky130_fd_sc_hd__or3b_1 _22019_ (.A(_01281_),
    .B(_01442_),
    .C_N(_01580_),
    .X(_01581_));
 sky130_fd_sc_hd__o21ba_1 _22020_ (.A1(_01310_),
    .A2(_01301_),
    .B1_N(_01496_),
    .X(_01582_));
 sky130_fd_sc_hd__o211a_1 _22021_ (.A1(net136),
    .A2(_01301_),
    .B1(_01487_),
    .C1(net166),
    .X(_01583_));
 sky130_fd_sc_hd__or2_1 _22022_ (.A(net152),
    .B(net136),
    .X(_01584_));
 sky130_fd_sc_hd__and3_1 _22023_ (.A(_01356_),
    .B(_01487_),
    .C(_01584_),
    .X(_01585_));
 sky130_fd_sc_hd__a2111o_1 _22024_ (.A1(_01281_),
    .A2(_01582_),
    .B1(_01583_),
    .C1(net145),
    .D1(_01585_),
    .X(_01586_));
 sky130_fd_sc_hd__o311a_1 _22025_ (.A1(net153),
    .A2(_01299_),
    .A3(_01578_),
    .B1(_01581_),
    .C1(_01586_),
    .X(_01587_));
 sky130_fd_sc_hd__o31a_1 _22026_ (.A1(_01574_),
    .A2(_01576_),
    .A3(_01577_),
    .B1(_01587_),
    .X(_01588_));
 sky130_fd_sc_hd__xnor2_1 _22027_ (.A(_01568_),
    .B(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__xnor2_2 _22028_ (.A(_01560_),
    .B(_01589_),
    .Y(_01590_));
 sky130_fd_sc_hd__inv_2 _22029_ (.A(_01590_),
    .Y(_01591_));
 sky130_fd_sc_hd__mux2_1 _22030_ (.A0(_01372_),
    .A1(_01393_),
    .S(net142),
    .X(_01592_));
 sky130_fd_sc_hd__inv_2 _22031_ (.A(_01592_),
    .Y(_01593_));
 sky130_fd_sc_hd__a22o_1 _22032_ (.A1(_01177_),
    .A2(_01306_),
    .B1(_01593_),
    .B2(net146),
    .X(_01594_));
 sky130_fd_sc_hd__a22o_1 _22033_ (.A1(_01355_),
    .A2(_01275_),
    .B1(_01594_),
    .B2(net162),
    .X(_01595_));
 sky130_fd_sc_hd__o21bai_2 _22034_ (.A1(_01265_),
    .A2(_01279_),
    .B1_N(_01278_),
    .Y(_01596_));
 sky130_fd_sc_hd__xnor2_1 _22035_ (.A(_01289_),
    .B(_01596_),
    .Y(_01597_));
 sky130_fd_sc_hd__a21bo_1 _22036_ (.A1(_01595_),
    .A2(_01597_),
    .B1_N(_01316_),
    .X(_01598_));
 sky130_fd_sc_hd__o21a_1 _22037_ (.A1(_01595_),
    .A2(_01597_),
    .B1(_01598_),
    .X(_01599_));
 sky130_fd_sc_hd__a31o_1 _22038_ (.A1(net122),
    .A2(net113),
    .A3(net106),
    .B1(_01596_),
    .X(_01600_));
 sky130_fd_sc_hd__or2_1 _22039_ (.A(net146),
    .B(_01081_),
    .X(_01601_));
 sky130_fd_sc_hd__a21o_1 _22040_ (.A1(_01262_),
    .A2(_01601_),
    .B1(_01151_),
    .X(_01602_));
 sky130_fd_sc_hd__o2111a_1 _22041_ (.A1(_01262_),
    .A2(_01601_),
    .B1(_01602_),
    .C1(net106),
    .D1(net122),
    .X(_01603_));
 sky130_fd_sc_hd__a221oi_2 _22042_ (.A1(_01213_),
    .A2(_01286_),
    .B1(_01287_),
    .B2(_01600_),
    .C1(_01603_),
    .Y(_01604_));
 sky130_fd_sc_hd__or2_1 _22043_ (.A(_01599_),
    .B(_01604_),
    .X(_01605_));
 sky130_fd_sc_hd__or2_1 _22044_ (.A(_01362_),
    .B(_01335_),
    .X(_01606_));
 sky130_fd_sc_hd__nor2_1 _22045_ (.A(_01334_),
    .B(_01347_),
    .Y(_01607_));
 sky130_fd_sc_hd__a32o_1 _22046_ (.A1(_01606_),
    .A2(_01348_),
    .A3(_01353_),
    .B1(_01607_),
    .B2(_01362_),
    .X(_01608_));
 sky130_fd_sc_hd__nor2_1 _22047_ (.A(_01318_),
    .B(_01608_),
    .Y(_01609_));
 sky130_fd_sc_hd__o22a_1 _22048_ (.A1(_01591_),
    .A2(_01605_),
    .B1(_01609_),
    .B2(_01363_),
    .X(_01610_));
 sky130_fd_sc_hd__nand2_1 _22049_ (.A(_01599_),
    .B(_01604_),
    .Y(_01611_));
 sky130_fd_sc_hd__a21boi_1 _22050_ (.A1(_01590_),
    .A2(_01611_),
    .B1_N(_01605_),
    .Y(_01612_));
 sky130_fd_sc_hd__xnor2_2 _22051_ (.A(_01180_),
    .B(_01181_),
    .Y(_01613_));
 sky130_fd_sc_hd__xnor2_4 _22052_ (.A(_01174_),
    .B(_01613_),
    .Y(_01614_));
 sky130_fd_sc_hd__nand2_2 _22053_ (.A(net115),
    .B(net97),
    .Y(_01615_));
 sky130_fd_sc_hd__nand2_2 _22054_ (.A(net119),
    .B(net105),
    .Y(_01616_));
 sky130_fd_sc_hd__nand2_2 _22055_ (.A(net102),
    .B(_01616_),
    .Y(_01617_));
 sky130_fd_sc_hd__xor2_4 _22056_ (.A(_01615_),
    .B(_01617_),
    .X(_01618_));
 sky130_fd_sc_hd__xnor2_4 _22057_ (.A(_01614_),
    .B(_01618_),
    .Y(_01619_));
 sky130_fd_sc_hd__inv_2 _22058_ (.A(_01558_),
    .Y(_01620_));
 sky130_fd_sc_hd__or2_1 _22059_ (.A(_01549_),
    .B(_01553_),
    .X(_01621_));
 sky130_fd_sc_hd__a21o_1 _22060_ (.A1(_01549_),
    .A2(_01553_),
    .B1(_01552_),
    .X(_01622_));
 sky130_fd_sc_hd__and3_1 _22061_ (.A(_01552_),
    .B(_01549_),
    .C(_01553_),
    .X(_01623_));
 sky130_fd_sc_hd__a31oi_1 _22062_ (.A1(_01557_),
    .A2(_01621_),
    .A3(_01622_),
    .B1(_01623_),
    .Y(_01624_));
 sky130_fd_sc_hd__a211o_1 _22063_ (.A1(_01557_),
    .A2(_01558_),
    .B1(_01621_),
    .C1(_01552_),
    .X(_01625_));
 sky130_fd_sc_hd__nand2_1 _22064_ (.A(_01557_),
    .B(_01623_),
    .Y(_01626_));
 sky130_fd_sc_hd__a211o_1 _22065_ (.A1(_01621_),
    .A2(_01622_),
    .B1(_01558_),
    .C1(_01557_),
    .X(_01627_));
 sky130_fd_sc_hd__o2111a_2 _22066_ (.A1(_01620_),
    .A2(_01624_),
    .B1(_01625_),
    .C1(_01626_),
    .D1(_01627_),
    .X(_01628_));
 sky130_fd_sc_hd__xor2_2 _22067_ (.A(_01619_),
    .B(_01628_),
    .X(_01629_));
 sky130_fd_sc_hd__a31o_1 _22068_ (.A1(net118),
    .A2(net106),
    .A3(net102),
    .B1(_01563_),
    .X(_01630_));
 sky130_fd_sc_hd__mux2_1 _22069_ (.A0(_01563_),
    .A1(_01211_),
    .S(_01564_),
    .X(_01631_));
 sky130_fd_sc_hd__a21oi_2 _22070_ (.A1(_01565_),
    .A2(_01630_),
    .B1(_01631_),
    .Y(_01632_));
 sky130_fd_sc_hd__nand2b_1 _22071_ (.A_N(_01588_),
    .B(_01568_),
    .Y(_01633_));
 sky130_fd_sc_hd__and2b_1 _22072_ (.A_N(_01568_),
    .B(_01588_),
    .X(_01634_));
 sky130_fd_sc_hd__a21oi_2 _22073_ (.A1(_01560_),
    .A2(_01633_),
    .B1(_01634_),
    .Y(_01635_));
 sky130_fd_sc_hd__xnor2_2 _22074_ (.A(_01632_),
    .B(_01635_),
    .Y(_01636_));
 sky130_fd_sc_hd__xnor2_4 _22075_ (.A(_01629_),
    .B(_01636_),
    .Y(_01637_));
 sky130_fd_sc_hd__o21ai_1 _22076_ (.A1(_01610_),
    .A2(_01612_),
    .B1(_01637_),
    .Y(_01638_));
 sky130_fd_sc_hd__xnor2_1 _22077_ (.A(_01193_),
    .B(_01184_),
    .Y(_01639_));
 sky130_fd_sc_hd__xnor2_2 _22078_ (.A(_01190_),
    .B(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hd__and2_1 _22079_ (.A(_01621_),
    .B(_01622_),
    .X(_01641_));
 sky130_fd_sc_hd__a31o_1 _22080_ (.A1(net115),
    .A2(net102),
    .A3(net97),
    .B1(_01641_),
    .X(_01642_));
 sky130_fd_sc_hd__clkbuf_4 _22081_ (.A(_01066_),
    .X(_01643_));
 sky130_fd_sc_hd__mux2_1 _22082_ (.A0(_01641_),
    .A1(_01643_),
    .S(_01615_),
    .X(_01644_));
 sky130_fd_sc_hd__a21oi_2 _22083_ (.A1(_01616_),
    .A2(_01642_),
    .B1(_01644_),
    .Y(_01645_));
 sky130_fd_sc_hd__or2_1 _22084_ (.A(_01640_),
    .B(_01645_),
    .X(_01646_));
 sky130_fd_sc_hd__nand2_1 _22085_ (.A(_01640_),
    .B(_01645_),
    .Y(_01647_));
 sky130_fd_sc_hd__nand2_1 _22086_ (.A(_01647_),
    .B(_01646_),
    .Y(_01648_));
 sky130_fd_sc_hd__o21ba_1 _22087_ (.A1(_01557_),
    .A2(_01558_),
    .B1_N(_01555_),
    .X(_01649_));
 sky130_fd_sc_hd__a21oi_1 _22088_ (.A1(_01557_),
    .A2(_01558_),
    .B1(_01649_),
    .Y(_01650_));
 sky130_fd_sc_hd__xnor2_1 _22089_ (.A(_01618_),
    .B(_01641_),
    .Y(_01651_));
 sky130_fd_sc_hd__o21a_1 _22090_ (.A1(_01650_),
    .A2(_01651_),
    .B1(_01614_),
    .X(_01652_));
 sky130_fd_sc_hd__a21o_1 _22091_ (.A1(_01650_),
    .A2(_01651_),
    .B1(_01652_),
    .X(_01653_));
 sky130_fd_sc_hd__nor2_1 _22092_ (.A(_01619_),
    .B(_01628_),
    .Y(_01654_));
 sky130_fd_sc_hd__and2_1 _22093_ (.A(_01619_),
    .B(_01628_),
    .X(_01655_));
 sky130_fd_sc_hd__inv_2 _22094_ (.A(_01635_),
    .Y(_01656_));
 sky130_fd_sc_hd__and2b_1 _22095_ (.A_N(_01628_),
    .B(_01632_),
    .X(_01657_));
 sky130_fd_sc_hd__and2_1 _22096_ (.A(_01628_),
    .B(_01632_),
    .X(_01658_));
 sky130_fd_sc_hd__mux2_1 _22097_ (.A0(_01657_),
    .A1(_01658_),
    .S(_01619_),
    .X(_01659_));
 sky130_fd_sc_hd__o32a_2 _22098_ (.A1(_01654_),
    .A2(_01655_),
    .A3(_01632_),
    .B1(_01656_),
    .B2(_01659_),
    .X(_01660_));
 sky130_fd_sc_hd__nor2_1 _22099_ (.A(_01653_),
    .B(_01660_),
    .Y(_01661_));
 sky130_fd_sc_hd__mux2_1 _22100_ (.A0(_01646_),
    .A1(_01648_),
    .S(_01661_),
    .X(_01662_));
 sky130_fd_sc_hd__inv_2 _22101_ (.A(_01647_),
    .Y(_01663_));
 sky130_fd_sc_hd__mux2_1 _22102_ (.A0(_01660_),
    .A1(_01640_),
    .S(_01645_),
    .X(_01664_));
 sky130_fd_sc_hd__a22oi_1 _22103_ (.A1(_01663_),
    .A2(_01660_),
    .B1(_01664_),
    .B2(_01653_),
    .Y(_01665_));
 sky130_fd_sc_hd__xnor2_1 _22104_ (.A(_01195_),
    .B(_01087_),
    .Y(_01666_));
 sky130_fd_sc_hd__xnor2_1 _22105_ (.A(_01172_),
    .B(_01666_),
    .Y(_01667_));
 sky130_fd_sc_hd__mux2_1 _22106_ (.A0(_01662_),
    .A1(_01665_),
    .S(_01667_),
    .X(_01668_));
 sky130_fd_sc_hd__o21ba_1 _22107_ (.A1(_01406_),
    .A2(_01608_),
    .B1_N(_01363_),
    .X(_01669_));
 sky130_fd_sc_hd__nor2b_1 _22108_ (.A(_01637_),
    .B_N(_01611_),
    .Y(_01670_));
 sky130_fd_sc_hd__nand2_1 _22109_ (.A(_01637_),
    .B(_01605_),
    .Y(_01671_));
 sky130_fd_sc_hd__o221a_1 _22110_ (.A1(_01318_),
    .A2(_01669_),
    .B1(_01670_),
    .B2(_01590_),
    .C1(_01671_),
    .X(_01672_));
 sky130_fd_sc_hd__and3b_1 _22111_ (.A_N(_01640_),
    .B(_01660_),
    .C(_01653_),
    .X(_01673_));
 sky130_fd_sc_hd__and3_1 _22112_ (.A(_01406_),
    .B(_01318_),
    .C(_01608_),
    .X(_01674_));
 sky130_fd_sc_hd__inv_2 _22113_ (.A(_01674_),
    .Y(_01675_));
 sky130_fd_sc_hd__nor2_1 _22114_ (.A(_01637_),
    .B(_01675_),
    .Y(_01676_));
 sky130_fd_sc_hd__a21oi_1 _22115_ (.A1(_01637_),
    .A2(_01675_),
    .B1(_01612_),
    .Y(_01677_));
 sky130_fd_sc_hd__or4_1 _22116_ (.A(_01672_),
    .B(_01673_),
    .C(_01676_),
    .D(_01677_),
    .X(_01678_));
 sky130_fd_sc_hd__a311o_1 _22117_ (.A1(_01452_),
    .A2(_01547_),
    .A3(_01638_),
    .B1(_01668_),
    .C1(_01678_),
    .X(_01679_));
 sky130_fd_sc_hd__a211oi_1 _22118_ (.A1(_01653_),
    .A2(_01645_),
    .B1(_01660_),
    .C1(_01640_),
    .Y(_01680_));
 sky130_fd_sc_hd__a211o_1 _22119_ (.A1(_01640_),
    .A2(_01660_),
    .B1(_01645_),
    .C1(_01653_),
    .X(_01681_));
 sky130_fd_sc_hd__or3b_1 _22120_ (.A(_01667_),
    .B(_01680_),
    .C_N(_01681_),
    .X(_01682_));
 sky130_fd_sc_hd__a22o_1 _22121_ (.A1(_01197_),
    .A2(_01257_),
    .B1(_01679_),
    .B2(_01682_),
    .X(_01683_));
 sky130_fd_sc_hd__nand2_2 _22122_ (.A(_01258_),
    .B(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__and3_1 _22123_ (.A(net78),
    .B(net99),
    .C(net86),
    .X(_01685_));
 sky130_fd_sc_hd__nor2_1 _22124_ (.A(_01215_),
    .B(_01219_),
    .Y(_01686_));
 sky130_fd_sc_hd__or2_1 _22125_ (.A(_01063_),
    .B(_01225_),
    .X(_01687_));
 sky130_fd_sc_hd__nand2_1 _22126_ (.A(_01063_),
    .B(_01225_),
    .Y(_01688_));
 sky130_fd_sc_hd__and3_1 _22127_ (.A(_11444_),
    .B(_01687_),
    .C(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__a21oi_1 _22128_ (.A1(net96),
    .A2(_01225_),
    .B1(_11674_),
    .Y(_01690_));
 sky130_fd_sc_hd__nand2_1 _22129_ (.A(_01215_),
    .B(_01219_),
    .Y(_01691_));
 sky130_fd_sc_hd__o21ai_1 _22130_ (.A1(_01225_),
    .A2(_01686_),
    .B1(_01691_),
    .Y(_01692_));
 sky130_fd_sc_hd__mux2_1 _22131_ (.A0(_01692_),
    .A1(_01691_),
    .S(_01221_),
    .X(_01693_));
 sky130_fd_sc_hd__o31a_1 _22132_ (.A1(_01686_),
    .A2(_01689_),
    .A3(_01690_),
    .B1(_01693_),
    .X(_01694_));
 sky130_fd_sc_hd__xor2_2 _22133_ (.A(_01685_),
    .B(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__nor2_1 _22134_ (.A(_01210_),
    .B(_01227_),
    .Y(_01696_));
 sky130_fd_sc_hd__nand2_1 _22135_ (.A(_01210_),
    .B(_01227_),
    .Y(_01697_));
 sky130_fd_sc_hd__o21ai_2 _22136_ (.A1(_01205_),
    .A2(_01696_),
    .B1(_01697_),
    .Y(_01698_));
 sky130_fd_sc_hd__and2_1 _22137_ (.A(_01139_),
    .B(_01208_),
    .X(_01699_));
 sky130_fd_sc_hd__o211a_1 _22138_ (.A1(net138),
    .A2(_01076_),
    .B1(_01206_),
    .C1(_01458_),
    .X(_01700_));
 sky130_fd_sc_hd__o22ai_1 _22139_ (.A1(_01076_),
    .A2(_01206_),
    .B1(_01699_),
    .B2(_01700_),
    .Y(_01701_));
 sky130_fd_sc_hd__or2_1 _22140_ (.A(_01311_),
    .B(_01076_),
    .X(_01702_));
 sky130_fd_sc_hd__nand2_1 _22141_ (.A(_01311_),
    .B(_01076_),
    .Y(_01703_));
 sky130_fd_sc_hd__and4_1 _22142_ (.A(net133),
    .B(_01208_),
    .C(_01702_),
    .D(_01703_),
    .X(_01704_));
 sky130_fd_sc_hd__nor3_1 _22143_ (.A(net133),
    .B(_01076_),
    .C(_01208_),
    .Y(_01705_));
 sky130_fd_sc_hd__a211o_2 _22144_ (.A1(net155),
    .A2(_01701_),
    .B1(_01704_),
    .C1(_01705_),
    .X(_01706_));
 sky130_fd_sc_hd__nand2_1 _22145_ (.A(_01105_),
    .B(net127),
    .Y(_01707_));
 sky130_fd_sc_hd__nand2_1 _22146_ (.A(net132),
    .B(_01135_),
    .Y(_01708_));
 sky130_fd_sc_hd__mux2_1 _22147_ (.A0(_01707_),
    .A1(_01708_),
    .S(net149),
    .X(_01709_));
 sky130_fd_sc_hd__xnor2_1 _22148_ (.A(_01144_),
    .B(_01456_),
    .Y(_01710_));
 sky130_fd_sc_hd__xnor2_2 _22149_ (.A(_01709_),
    .B(_01710_),
    .Y(_01711_));
 sky130_fd_sc_hd__o21a_1 _22150_ (.A1(net99),
    .A2(_01223_),
    .B1(_01211_),
    .X(_01712_));
 sky130_fd_sc_hd__and4bb_1 _22151_ (.A_N(net99),
    .B_N(_01223_),
    .C(net110),
    .D(net105),
    .X(_01713_));
 sky130_fd_sc_hd__a311o_1 _22152_ (.A1(_01213_),
    .A2(net99),
    .A3(_01223_),
    .B1(_01712_),
    .C1(_01713_),
    .X(_01714_));
 sky130_fd_sc_hd__nand2_1 _22153_ (.A(net124),
    .B(_01065_),
    .Y(_01715_));
 sky130_fd_sc_hd__a221o_2 _22154_ (.A1(net114),
    .A2(_01075_),
    .B1(_01260_),
    .B2(_01715_),
    .C1(_01133_),
    .X(_01716_));
 sky130_fd_sc_hd__xnor2_1 _22155_ (.A(net90),
    .B(_01716_),
    .Y(_01717_));
 sky130_fd_sc_hd__xnor2_2 _22156_ (.A(_01714_),
    .B(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__xor2_1 _22157_ (.A(_01711_),
    .B(_01718_),
    .X(_01719_));
 sky130_fd_sc_hd__xnor2_2 _22158_ (.A(_01706_),
    .B(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__xnor2_1 _22159_ (.A(_01698_),
    .B(_01720_),
    .Y(_01721_));
 sky130_fd_sc_hd__xnor2_2 _22160_ (.A(_01695_),
    .B(_01721_),
    .Y(_01722_));
 sky130_fd_sc_hd__a21o_1 _22161_ (.A1(_01229_),
    .A2(_01242_),
    .B1(_01245_),
    .X(_01723_));
 sky130_fd_sc_hd__o21a_1 _22162_ (.A1(_01229_),
    .A2(_01242_),
    .B1(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__a21o_1 _22163_ (.A1(net105),
    .A2(net90),
    .B1(_01235_),
    .X(_01725_));
 sky130_fd_sc_hd__a21bo_1 _22164_ (.A1(_01231_),
    .A2(_01235_),
    .B1_N(_01232_),
    .X(_01726_));
 sky130_fd_sc_hd__o211a_1 _22165_ (.A1(net86),
    .A2(_01232_),
    .B1(_01725_),
    .C1(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__xnor2_1 _22166_ (.A(_01724_),
    .B(_01727_),
    .Y(_01728_));
 sky130_fd_sc_hd__xnor2_2 _22167_ (.A(_01722_),
    .B(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__nand2_1 _22168_ (.A(_01249_),
    .B(_01247_),
    .Y(_01730_));
 sky130_fd_sc_hd__o2bb2a_1 _22169_ (.A1_N(_01160_),
    .A2_N(_01730_),
    .B1(_01165_),
    .B2(_01247_),
    .X(_01731_));
 sky130_fd_sc_hd__nor2_1 _22170_ (.A(_01250_),
    .B(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__inv_2 _22171_ (.A(_01165_),
    .Y(_01733_));
 sky130_fd_sc_hd__a21oi_1 _22172_ (.A1(_01160_),
    .A2(_01733_),
    .B1(_01168_),
    .Y(_01734_));
 sky130_fd_sc_hd__a21oi_2 _22173_ (.A1(_01247_),
    .A2(_01253_),
    .B1(_01734_),
    .Y(_01735_));
 sky130_fd_sc_hd__nor2_1 _22174_ (.A(_01247_),
    .B(_01253_),
    .Y(_01736_));
 sky130_fd_sc_hd__or4_2 _22175_ (.A(_01729_),
    .B(_01732_),
    .C(_01735_),
    .D(_01736_),
    .X(_01737_));
 sky130_fd_sc_hd__o31ai_4 _22176_ (.A1(_01732_),
    .A2(_01735_),
    .A3(_01736_),
    .B1(_01729_),
    .Y(_01738_));
 sky130_fd_sc_hd__nand2_1 _22177_ (.A(_01737_),
    .B(_01738_),
    .Y(_01739_));
 sky130_fd_sc_hd__xnor2_1 _22178_ (.A(_01684_),
    .B(_01739_),
    .Y(_01740_));
 sky130_fd_sc_hd__a22o_1 _22179_ (.A1(net745),
    .A2(_12813_),
    .B1(_01740_),
    .B2(_12963_),
    .X(_00397_));
 sky130_fd_sc_hd__o21a_1 _22180_ (.A1(_01724_),
    .A2(_01722_),
    .B1(_01727_),
    .X(_01741_));
 sky130_fd_sc_hd__a21o_2 _22181_ (.A1(_01724_),
    .A2(_01722_),
    .B1(_01741_),
    .X(_01742_));
 sky130_fd_sc_hd__nor2_1 _22182_ (.A(_01698_),
    .B(_01720_),
    .Y(_01743_));
 sky130_fd_sc_hd__nand2_1 _22183_ (.A(_01698_),
    .B(_01720_),
    .Y(_01744_));
 sky130_fd_sc_hd__o21a_2 _22184_ (.A1(_01695_),
    .A2(_01743_),
    .B1(_01744_),
    .X(_01745_));
 sky130_fd_sc_hd__nand2_1 _22185_ (.A(_01711_),
    .B(_01718_),
    .Y(_01746_));
 sky130_fd_sc_hd__nor2_1 _22186_ (.A(_01711_),
    .B(_01718_),
    .Y(_01747_));
 sky130_fd_sc_hd__a21oi_2 _22187_ (.A1(_01706_),
    .A2(_01746_),
    .B1(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__o21a_1 _22188_ (.A1(net131),
    .A2(_01144_),
    .B1(_01708_),
    .X(_01749_));
 sky130_fd_sc_hd__o2bb2a_1 _22189_ (.A1_N(_01089_),
    .A2_N(_01456_),
    .B1(_01708_),
    .B2(_01144_),
    .X(_01750_));
 sky130_fd_sc_hd__o21ai_2 _22190_ (.A1(_01456_),
    .A2(_01749_),
    .B1(_01750_),
    .Y(_01751_));
 sky130_fd_sc_hd__xnor2_1 _22191_ (.A(net132),
    .B(_01144_),
    .Y(_01752_));
 sky130_fd_sc_hd__nor3_1 _22192_ (.A(net127),
    .B(_01144_),
    .C(_01456_),
    .Y(_01753_));
 sky130_fd_sc_hd__a31o_1 _22193_ (.A1(net126),
    .A2(_01456_),
    .A3(_01752_),
    .B1(_01753_),
    .X(_01754_));
 sky130_fd_sc_hd__a21oi_4 _22194_ (.A1(net149),
    .A2(_01751_),
    .B1(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hd__xor2_2 _22195_ (.A(net78),
    .B(net89),
    .X(_01756_));
 sky130_fd_sc_hd__or2b_1 _22196_ (.A(net109),
    .B_N(net119),
    .X(_01757_));
 sky130_fd_sc_hd__a221o_2 _22197_ (.A1(net109),
    .A2(_01143_),
    .B1(_01757_),
    .B2(_01291_),
    .C1(_01116_),
    .X(_01758_));
 sky130_fd_sc_hd__or2b_1 _22198_ (.A(net95),
    .B_N(net104),
    .X(_01759_));
 sky130_fd_sc_hd__xnor2_1 _22199_ (.A(net77),
    .B(net92),
    .Y(_01760_));
 sky130_fd_sc_hd__and3b_1 _22200_ (.A_N(net104),
    .B(net100),
    .C(net95),
    .X(_01761_));
 sky130_fd_sc_hd__nor2_1 _22201_ (.A(net100),
    .B(net95),
    .Y(_01762_));
 sky130_fd_sc_hd__a211o_1 _22202_ (.A1(_01759_),
    .A2(_01760_),
    .B1(_01761_),
    .C1(_01762_),
    .X(_01763_));
 sky130_fd_sc_hd__xnor2_2 _22203_ (.A(_01758_),
    .B(_01763_),
    .Y(_01764_));
 sky130_fd_sc_hd__xnor2_4 _22204_ (.A(_01756_),
    .B(_01764_),
    .Y(_01765_));
 sky130_fd_sc_hd__and3b_1 _22205_ (.A_N(net124),
    .B(net126),
    .C(net144),
    .X(_01766_));
 sky130_fd_sc_hd__a21oi_1 _22206_ (.A1(_01102_),
    .A2(_01100_),
    .B1(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__xnor2_2 _22207_ (.A(_01412_),
    .B(_01767_),
    .Y(_01768_));
 sky130_fd_sc_hd__nor2b_4 _22208_ (.A(net100),
    .B_N(net95),
    .Y(_01769_));
 sky130_fd_sc_hd__xnor2_4 _22209_ (.A(_01166_),
    .B(_01769_),
    .Y(_01770_));
 sky130_fd_sc_hd__xor2_2 _22210_ (.A(_01113_),
    .B(_01770_),
    .X(_01771_));
 sky130_fd_sc_hd__xnor2_1 _22211_ (.A(_01768_),
    .B(_01771_),
    .Y(_01772_));
 sky130_fd_sc_hd__xnor2_2 _22212_ (.A(_01765_),
    .B(_01772_),
    .Y(_01773_));
 sky130_fd_sc_hd__xnor2_2 _22213_ (.A(_01755_),
    .B(_01773_),
    .Y(_01774_));
 sky130_fd_sc_hd__nor2b_2 _22214_ (.A(net98),
    .B_N(net94),
    .Y(_01775_));
 sky130_fd_sc_hd__nor2b_1 _22215_ (.A(net90),
    .B_N(net96),
    .Y(_01776_));
 sky130_fd_sc_hd__nand2_4 _22216_ (.A(_01211_),
    .B(net102),
    .Y(_01777_));
 sky130_fd_sc_hd__nor2_1 _22217_ (.A(_01213_),
    .B(net100),
    .Y(_01778_));
 sky130_fd_sc_hd__mux2_1 _22218_ (.A0(net104),
    .A1(_01224_),
    .S(net100),
    .X(_01779_));
 sky130_fd_sc_hd__o21ai_1 _22219_ (.A1(_01223_),
    .A2(_01778_),
    .B1(_01779_),
    .Y(_01780_));
 sky130_fd_sc_hd__nand2_1 _22220_ (.A(_01716_),
    .B(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__nor2_1 _22221_ (.A(_01716_),
    .B(_01780_),
    .Y(_01782_));
 sky130_fd_sc_hd__a21oi_1 _22222_ (.A1(_01777_),
    .A2(_01781_),
    .B1(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__inv_2 _22223_ (.A(_01777_),
    .Y(_01784_));
 sky130_fd_sc_hd__nor2_1 _22224_ (.A(_01775_),
    .B(_01776_),
    .Y(_01785_));
 sky130_fd_sc_hd__o21a_1 _22225_ (.A1(_01784_),
    .A2(_01785_),
    .B1(net77),
    .X(_01786_));
 sky130_fd_sc_hd__or2_1 _22226_ (.A(_01777_),
    .B(_01785_),
    .X(_01787_));
 sky130_fd_sc_hd__nand2_1 _22227_ (.A(_01777_),
    .B(_01785_),
    .Y(_01788_));
 sky130_fd_sc_hd__and3_1 _22228_ (.A(_11444_),
    .B(_01787_),
    .C(_01788_),
    .X(_01789_));
 sky130_fd_sc_hd__and2_1 _22229_ (.A(net77),
    .B(_01785_),
    .X(_01790_));
 sky130_fd_sc_hd__o32a_1 _22230_ (.A1(_01782_),
    .A2(_01786_),
    .A3(_01789_),
    .B1(_01781_),
    .B2(_01790_),
    .X(_01791_));
 sky130_fd_sc_hd__o41a_1 _22231_ (.A1(_11674_),
    .A2(_01775_),
    .A3(_01776_),
    .A4(_01783_),
    .B1(_01791_),
    .X(_01792_));
 sky130_fd_sc_hd__and2_1 _22232_ (.A(_01774_),
    .B(_01792_),
    .X(_01793_));
 sky130_fd_sc_hd__nor2_1 _22233_ (.A(_01774_),
    .B(_01792_),
    .Y(_01794_));
 sky130_fd_sc_hd__nor2_1 _22234_ (.A(_01793_),
    .B(_01794_),
    .Y(_01795_));
 sky130_fd_sc_hd__xnor2_2 _22235_ (.A(_01748_),
    .B(_01795_),
    .Y(_01796_));
 sky130_fd_sc_hd__nor2_1 _22236_ (.A(_01685_),
    .B(_01686_),
    .Y(_01797_));
 sky130_fd_sc_hd__nor2_1 _22237_ (.A(_01643_),
    .B(net95),
    .Y(_01798_));
 sky130_fd_sc_hd__a221o_1 _22238_ (.A1(_01213_),
    .A2(net106),
    .B1(net100),
    .B2(net87),
    .C1(_01762_),
    .X(_01799_));
 sky130_fd_sc_hd__o211a_1 _22239_ (.A1(_01224_),
    .A2(_01798_),
    .B1(_01799_),
    .C1(net80),
    .X(_01800_));
 sky130_fd_sc_hd__a2bb2o_2 _22240_ (.A1_N(_01221_),
    .A2_N(_01797_),
    .B1(_01800_),
    .B2(_01691_),
    .X(_01801_));
 sky130_fd_sc_hd__xor2_2 _22241_ (.A(_01796_),
    .B(_01801_),
    .X(_01802_));
 sky130_fd_sc_hd__xor2_2 _22242_ (.A(_01745_),
    .B(_01802_),
    .X(_01803_));
 sky130_fd_sc_hd__nand2_1 _22243_ (.A(_01742_),
    .B(_01803_),
    .Y(_01804_));
 sky130_fd_sc_hd__or2_1 _22244_ (.A(_01742_),
    .B(_01803_),
    .X(_01805_));
 sky130_fd_sc_hd__nand2_2 _22245_ (.A(_01804_),
    .B(_01805_),
    .Y(_01806_));
 sky130_fd_sc_hd__or2_1 _22246_ (.A(_01684_),
    .B(_01737_),
    .X(_01807_));
 sky130_fd_sc_hd__nand2_1 _22247_ (.A(net210),
    .B(_01684_),
    .Y(_01808_));
 sky130_fd_sc_hd__a21bo_2 _22248_ (.A1(_01684_),
    .A2(_01737_),
    .B1_N(_01738_),
    .X(_01809_));
 sky130_fd_sc_hd__a32o_1 _22249_ (.A1(net210),
    .A2(_01738_),
    .A3(_01807_),
    .B1(_01808_),
    .B2(_01809_),
    .X(_01810_));
 sky130_fd_sc_hd__xor2_1 _22250_ (.A(_01806_),
    .B(_01810_),
    .X(_01811_));
 sky130_fd_sc_hd__nor2_1 _22251_ (.A(_12036_),
    .B(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__a31o_1 _22252_ (.A1(net721),
    .A2(_12034_),
    .A3(_12037_),
    .B1(_01812_),
    .X(_00398_));
 sky130_fd_sc_hd__o21a_1 _22253_ (.A1(_01803_),
    .A2(_01809_),
    .B1(_01742_),
    .X(_01813_));
 sky130_fd_sc_hd__a21oi_1 _22254_ (.A1(_01803_),
    .A2(_01809_),
    .B1(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__xnor2_2 _22255_ (.A(_01765_),
    .B(_01770_),
    .Y(_01815_));
 sky130_fd_sc_hd__xnor2_1 _22256_ (.A(_01113_),
    .B(_01768_),
    .Y(_01816_));
 sky130_fd_sc_hd__o21a_1 _22257_ (.A1(_01755_),
    .A2(_01815_),
    .B1(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__a21oi_4 _22258_ (.A1(_01755_),
    .A2(_01815_),
    .B1(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__nor2_1 _22259_ (.A(_01758_),
    .B(_01763_),
    .Y(_01819_));
 sky130_fd_sc_hd__and2b_1 _22260_ (.A_N(net91),
    .B(net87),
    .X(_01820_));
 sky130_fd_sc_hd__nor2_2 _22261_ (.A(_01166_),
    .B(net89),
    .Y(_01821_));
 sky130_fd_sc_hd__nor2_1 _22262_ (.A(_01820_),
    .B(_01821_),
    .Y(_01822_));
 sky130_fd_sc_hd__o21a_1 _22263_ (.A1(_01769_),
    .A2(_01822_),
    .B1(net77),
    .X(_01823_));
 sky130_fd_sc_hd__nand2_1 _22264_ (.A(_01066_),
    .B(net96),
    .Y(_01824_));
 sky130_fd_sc_hd__or2_1 _22265_ (.A(_01824_),
    .B(_01822_),
    .X(_01825_));
 sky130_fd_sc_hd__nand2_1 _22266_ (.A(_01824_),
    .B(_01822_),
    .Y(_01826_));
 sky130_fd_sc_hd__and3_1 _22267_ (.A(_11674_),
    .B(_01825_),
    .C(_01826_),
    .X(_01827_));
 sky130_fd_sc_hd__nand2_1 _22268_ (.A(_01758_),
    .B(_01763_),
    .Y(_01828_));
 sky130_fd_sc_hd__a21oi_1 _22269_ (.A1(_01824_),
    .A2(_01828_),
    .B1(_01819_),
    .Y(_01829_));
 sky130_fd_sc_hd__nand2_1 _22270_ (.A(net77),
    .B(_01822_),
    .Y(_01830_));
 sky130_fd_sc_hd__mux2_1 _22271_ (.A0(_01829_),
    .A1(_01828_),
    .S(_01830_),
    .X(_01831_));
 sky130_fd_sc_hd__o31a_2 _22272_ (.A1(_01819_),
    .A2(_01823_),
    .A3(_01827_),
    .B1(_01831_),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _22273_ (.A0(_01135_),
    .A1(_01412_),
    .S(_01113_),
    .X(_01833_));
 sky130_fd_sc_hd__or3b_1 _22274_ (.A(net143),
    .B(net126),
    .C_N(_01113_),
    .X(_01834_));
 sky130_fd_sc_hd__o211a_1 _22275_ (.A1(net143),
    .A2(_01412_),
    .B1(_01833_),
    .C1(_01834_),
    .X(_01835_));
 sky130_fd_sc_hd__nand2_1 _22276_ (.A(_01113_),
    .B(_01412_),
    .Y(_01836_));
 sky130_fd_sc_hd__nor2_1 _22277_ (.A(_01113_),
    .B(_01412_),
    .Y(_01837_));
 sky130_fd_sc_hd__a31o_1 _22278_ (.A1(net144),
    .A2(net126),
    .A3(_01836_),
    .B1(_01837_),
    .X(_01838_));
 sky130_fd_sc_hd__mux2_2 _22279_ (.A0(_01835_),
    .A1(_01838_),
    .S(_01408_),
    .X(_01839_));
 sky130_fd_sc_hd__and3_1 _22280_ (.A(net139),
    .B(net123),
    .C(_01217_),
    .X(_01840_));
 sky130_fd_sc_hd__a21o_1 _22281_ (.A1(_01311_),
    .A2(_01075_),
    .B1(_01840_),
    .X(_01841_));
 sky130_fd_sc_hd__xnor2_1 _22282_ (.A(_01225_),
    .B(_01328_),
    .Y(_01842_));
 sky130_fd_sc_hd__xnor2_2 _22283_ (.A(_01841_),
    .B(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__nand2_1 _22284_ (.A(net115),
    .B(_01211_),
    .Y(_01844_));
 sky130_fd_sc_hd__a21o_2 _22285_ (.A1(_01844_),
    .A2(_01550_),
    .B1(_01214_),
    .X(_01845_));
 sky130_fd_sc_hd__and2_1 _22286_ (.A(net101),
    .B(net96),
    .X(_01846_));
 sky130_fd_sc_hd__o21ai_1 _22287_ (.A1(net101),
    .A2(net86),
    .B1(net96),
    .Y(_01847_));
 sky130_fd_sc_hd__mux2_1 _22288_ (.A0(_01846_),
    .A1(_01847_),
    .S(net81),
    .X(_01848_));
 sky130_fd_sc_hd__nand2_1 _22289_ (.A(net90),
    .B(net86),
    .Y(_01849_));
 sky130_fd_sc_hd__nor2_1 _22290_ (.A(net78),
    .B(net99),
    .Y(_01850_));
 sky130_fd_sc_hd__a22o_1 _22291_ (.A1(net99),
    .A2(_01820_),
    .B1(_01849_),
    .B2(_01850_),
    .X(_01851_));
 sky130_fd_sc_hd__or2_2 _22292_ (.A(net95),
    .B(net91),
    .X(_01852_));
 sky130_fd_sc_hd__nor2_1 _22293_ (.A(net87),
    .B(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__a221o_1 _22294_ (.A1(net91),
    .A2(_01848_),
    .B1(_01851_),
    .B2(net95),
    .C1(_01853_),
    .X(_01854_));
 sky130_fd_sc_hd__xnor2_1 _22295_ (.A(_01845_),
    .B(_01854_),
    .Y(_01855_));
 sky130_fd_sc_hd__nor2_1 _22296_ (.A(_01843_),
    .B(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__nand2_1 _22297_ (.A(_01843_),
    .B(_01855_),
    .Y(_01857_));
 sky130_fd_sc_hd__or2b_1 _22298_ (.A(_01856_),
    .B_N(_01857_),
    .X(_01858_));
 sky130_fd_sc_hd__xnor2_2 _22299_ (.A(_01839_),
    .B(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__xor2_2 _22300_ (.A(_01832_),
    .B(_01859_),
    .X(_01860_));
 sky130_fd_sc_hd__xnor2_4 _22301_ (.A(_01818_),
    .B(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hd__nor2_1 _22302_ (.A(_01775_),
    .B(_01783_),
    .Y(_01862_));
 sky130_fd_sc_hd__o21a_1 _22303_ (.A1(_01776_),
    .A2(_01862_),
    .B1(net77),
    .X(_01863_));
 sky130_fd_sc_hd__nand2_1 _22304_ (.A(_01774_),
    .B(_01792_),
    .Y(_01864_));
 sky130_fd_sc_hd__o21ai_2 _22305_ (.A1(_01748_),
    .A2(_01794_),
    .B1(_01864_),
    .Y(_01865_));
 sky130_fd_sc_hd__xnor2_2 _22306_ (.A(_01863_),
    .B(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__xnor2_4 _22307_ (.A(_01861_),
    .B(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__nor2_1 _22308_ (.A(_01796_),
    .B(_01801_),
    .Y(_01868_));
 sky130_fd_sc_hd__nand2_1 _22309_ (.A(_01796_),
    .B(_01801_),
    .Y(_01869_));
 sky130_fd_sc_hd__inv_2 _22310_ (.A(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hd__nor2_1 _22311_ (.A(_01745_),
    .B(_01870_),
    .Y(_01871_));
 sky130_fd_sc_hd__nor2_1 _22312_ (.A(_01868_),
    .B(_01871_),
    .Y(_01872_));
 sky130_fd_sc_hd__xnor2_2 _22313_ (.A(_01867_),
    .B(_01872_),
    .Y(_01873_));
 sky130_fd_sc_hd__inv_2 _22314_ (.A(_01807_),
    .Y(_01874_));
 sky130_fd_sc_hd__mux2_1 _22315_ (.A0(_01738_),
    .A1(_01739_),
    .S(_01684_),
    .X(_01875_));
 sky130_fd_sc_hd__nor2_1 _22316_ (.A(_01806_),
    .B(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__inv_2 _22317_ (.A(net210),
    .Y(_01877_));
 sky130_fd_sc_hd__a211o_1 _22318_ (.A1(_01806_),
    .A2(_01874_),
    .B1(_01876_),
    .C1(_01877_),
    .X(_01878_));
 sky130_fd_sc_hd__xor2_1 _22319_ (.A(_01873_),
    .B(_01878_),
    .X(_01879_));
 sky130_fd_sc_hd__xnor2_1 _22320_ (.A(_01814_),
    .B(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__nor2_1 _22321_ (.A(_12036_),
    .B(_01880_),
    .Y(_01881_));
 sky130_fd_sc_hd__a31o_1 _22322_ (.A1(net749),
    .A2(_12034_),
    .A3(_12037_),
    .B1(_01881_),
    .X(_00399_));
 sky130_fd_sc_hd__or3_1 _22323_ (.A(_01684_),
    .B(_01737_),
    .C(_01804_),
    .X(_01882_));
 sky130_fd_sc_hd__o21ai_2 _22324_ (.A1(_01806_),
    .A2(_01875_),
    .B1(_01882_),
    .Y(_01883_));
 sky130_fd_sc_hd__or3_1 _22325_ (.A(_01805_),
    .B(_01807_),
    .C(_01873_),
    .X(_01884_));
 sky130_fd_sc_hd__a21boi_4 _22326_ (.A1(_01873_),
    .A2(_01883_),
    .B1_N(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__xor2_1 _22327_ (.A(_01742_),
    .B(_01745_),
    .X(_01886_));
 sky130_fd_sc_hd__mux2_1 _22328_ (.A0(_01868_),
    .A1(_01870_),
    .S(_01867_),
    .X(_01887_));
 sky130_fd_sc_hd__nor2_1 _22329_ (.A(_01745_),
    .B(_01867_),
    .Y(_01888_));
 sky130_fd_sc_hd__and2_1 _22330_ (.A(_01745_),
    .B(_01867_),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _22331_ (.A0(_01888_),
    .A1(_01889_),
    .S(_01742_),
    .X(_01890_));
 sky130_fd_sc_hd__a22o_1 _22332_ (.A1(_01886_),
    .A2(_01887_),
    .B1(_01890_),
    .B2(_01802_),
    .X(_01891_));
 sky130_fd_sc_hd__nand2_1 _22333_ (.A(_01867_),
    .B(_01869_),
    .Y(_01892_));
 sky130_fd_sc_hd__a2bb2o_1 _22334_ (.A1_N(_01867_),
    .A2_N(_01868_),
    .B1(_01892_),
    .B2(_01745_),
    .X(_01893_));
 sky130_fd_sc_hd__nand2_1 _22335_ (.A(_01742_),
    .B(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__o31a_1 _22336_ (.A1(_01867_),
    .A2(_01868_),
    .A3(_01871_),
    .B1(_01894_),
    .X(_01895_));
 sky130_fd_sc_hd__a21boi_2 _22337_ (.A1(_01809_),
    .A2(_01891_),
    .B1_N(_01895_),
    .Y(_01896_));
 sky130_fd_sc_hd__a21bo_1 _22338_ (.A1(_01863_),
    .A2(_01865_),
    .B1_N(_01861_),
    .X(_01897_));
 sky130_fd_sc_hd__o21a_1 _22339_ (.A1(_01863_),
    .A2(_01865_),
    .B1(_01897_),
    .X(_01898_));
 sky130_fd_sc_hd__o21a_1 _22340_ (.A1(_01839_),
    .A2(_01856_),
    .B1(_01857_),
    .X(_01899_));
 sky130_fd_sc_hd__nand2_1 _22341_ (.A(_01643_),
    .B(net91),
    .Y(_01900_));
 sky130_fd_sc_hd__a21oi_1 _22342_ (.A1(net97),
    .A2(_01900_),
    .B1(net78),
    .Y(_01901_));
 sky130_fd_sc_hd__o21ai_1 _22343_ (.A1(_01643_),
    .A2(net91),
    .B1(_01845_),
    .Y(_01902_));
 sky130_fd_sc_hd__nor2_1 _22344_ (.A(_01066_),
    .B(net91),
    .Y(_01903_));
 sky130_fd_sc_hd__o21ai_1 _22345_ (.A1(net78),
    .A2(_01903_),
    .B1(_01900_),
    .Y(_01904_));
 sky130_fd_sc_hd__o21a_1 _22346_ (.A1(_01845_),
    .A2(_01904_),
    .B1(_01230_),
    .X(_01905_));
 sky130_fd_sc_hd__a31o_1 _22347_ (.A1(net79),
    .A2(net87),
    .A3(_01902_),
    .B1(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__o21a_1 _22348_ (.A1(_11674_),
    .A2(_01845_),
    .B1(net87),
    .X(_01907_));
 sky130_fd_sc_hd__nor2_1 _22349_ (.A(_01852_),
    .B(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__a221o_1 _22350_ (.A1(_01845_),
    .A2(_01901_),
    .B1(_01906_),
    .B2(net97),
    .C1(_01908_),
    .X(_01909_));
 sky130_fd_sc_hd__nand2_1 _22351_ (.A(_01225_),
    .B(_01327_),
    .Y(_01910_));
 sky130_fd_sc_hd__a21o_1 _22352_ (.A1(_01225_),
    .A2(_01328_),
    .B1(_01311_),
    .X(_01911_));
 sky130_fd_sc_hd__o211a_1 _22353_ (.A1(_01225_),
    .A2(_01328_),
    .B1(_01911_),
    .C1(_01408_),
    .X(_01912_));
 sky130_fd_sc_hd__a21oi_1 _22354_ (.A1(net123),
    .A2(_01910_),
    .B1(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__nor2_1 _22355_ (.A(_01225_),
    .B(_01327_),
    .Y(_01914_));
 sky130_fd_sc_hd__a311o_1 _22356_ (.A1(net138),
    .A2(net123),
    .A3(_01910_),
    .B1(_01914_),
    .C1(\top0.cordic0.vec[1][9] ),
    .X(_01915_));
 sky130_fd_sc_hd__o21ai_2 _22357_ (.A1(_01217_),
    .A2(_01913_),
    .B1(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__xnor2_4 _22358_ (.A(_01062_),
    .B(_01777_),
    .Y(_01917_));
 sky130_fd_sc_hd__nor2_1 _22359_ (.A(_01217_),
    .B(net114),
    .Y(_01918_));
 sky130_fd_sc_hd__mux2_1 _22360_ (.A0(_01143_),
    .A1(_01918_),
    .S(net134),
    .X(_01919_));
 sky130_fd_sc_hd__xor2_1 _22361_ (.A(_01259_),
    .B(_01919_),
    .X(_01920_));
 sky130_fd_sc_hd__xnor2_2 _22362_ (.A(_01917_),
    .B(_01920_),
    .Y(_01921_));
 sky130_fd_sc_hd__a21o_1 _22363_ (.A1(net125),
    .A2(net120),
    .B1(_01778_),
    .X(_01922_));
 sky130_fd_sc_hd__nand2_1 _22364_ (.A(_01779_),
    .B(_01922_),
    .Y(_01923_));
 sky130_fd_sc_hd__buf_4 _22365_ (.A(_01820_),
    .X(_01924_));
 sky130_fd_sc_hd__nor2_1 _22366_ (.A(net86),
    .B(_01248_),
    .Y(_01925_));
 sky130_fd_sc_hd__nor2_1 _22367_ (.A(_01924_),
    .B(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hd__xnor2_1 _22368_ (.A(_11444_),
    .B(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__xnor2_1 _22369_ (.A(_01923_),
    .B(_01927_),
    .Y(_01928_));
 sky130_fd_sc_hd__xnor2_1 _22370_ (.A(_01921_),
    .B(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__xnor2_2 _22371_ (.A(_01916_),
    .B(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__nor2_1 _22372_ (.A(_01909_),
    .B(_01930_),
    .Y(_01931_));
 sky130_fd_sc_hd__nand2_1 _22373_ (.A(_01909_),
    .B(_01930_),
    .Y(_01932_));
 sky130_fd_sc_hd__and2b_1 _22374_ (.A_N(_01931_),
    .B(_01932_),
    .X(_01933_));
 sky130_fd_sc_hd__xnor2_2 _22375_ (.A(_01899_),
    .B(_01933_),
    .Y(_01934_));
 sky130_fd_sc_hd__o21a_1 _22376_ (.A1(_01832_),
    .A2(_01859_),
    .B1(_01818_),
    .X(_01935_));
 sky130_fd_sc_hd__a21oi_1 _22377_ (.A1(_01832_),
    .A2(_01859_),
    .B1(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__nand2_1 _22378_ (.A(net91),
    .B(_01230_),
    .Y(_01937_));
 sky130_fd_sc_hd__o21a_1 _22379_ (.A1(_01924_),
    .A2(_01829_),
    .B1(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__nor2_1 _22380_ (.A(_11674_),
    .B(_01938_),
    .Y(_01939_));
 sky130_fd_sc_hd__xnor2_1 _22381_ (.A(_01936_),
    .B(_01939_),
    .Y(_01940_));
 sky130_fd_sc_hd__xnor2_2 _22382_ (.A(_01934_),
    .B(_01940_),
    .Y(_01941_));
 sky130_fd_sc_hd__or2_1 _22383_ (.A(_01898_),
    .B(_01941_),
    .X(_01942_));
 sky130_fd_sc_hd__nand2_1 _22384_ (.A(_01898_),
    .B(_01941_),
    .Y(_01943_));
 sky130_fd_sc_hd__nand2_1 _22385_ (.A(_01942_),
    .B(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__xor2_1 _22386_ (.A(_01896_),
    .B(_01944_),
    .X(_01945_));
 sky130_fd_sc_hd__a21o_1 _22387_ (.A1(net210),
    .A2(_01885_),
    .B1(_01945_),
    .X(_01946_));
 sky130_fd_sc_hd__nand3_1 _22388_ (.A(net210),
    .B(_01885_),
    .C(_01945_),
    .Y(_01947_));
 sky130_fd_sc_hd__a32o_1 _22389_ (.A1(_12742_),
    .A2(_01946_),
    .A3(_01947_),
    .B1(_12812_),
    .B2(net712),
    .X(_00400_));
 sky130_fd_sc_hd__clkbuf_4 _22390_ (.A(_11674_),
    .X(_01948_));
 sky130_fd_sc_hd__or3_1 _22391_ (.A(_01948_),
    .B(_01934_),
    .C(_01938_),
    .X(_01949_));
 sky130_fd_sc_hd__and2b_1 _22392_ (.A_N(_01939_),
    .B(_01934_),
    .X(_01950_));
 sky130_fd_sc_hd__a21oi_1 _22393_ (.A1(_01936_),
    .A2(_01949_),
    .B1(_01950_),
    .Y(_01951_));
 sky130_fd_sc_hd__a21o_1 _22394_ (.A1(_01921_),
    .A2(_01928_),
    .B1(_01916_),
    .X(_01952_));
 sky130_fd_sc_hd__o21a_1 _22395_ (.A1(_01921_),
    .A2(_01928_),
    .B1(_01952_),
    .X(_01953_));
 sky130_fd_sc_hd__nor2_1 _22396_ (.A(\top0.cordic0.vec[1][10] ),
    .B(_01917_),
    .Y(_01954_));
 sky130_fd_sc_hd__nor2_1 _22397_ (.A(net119),
    .B(_01917_),
    .Y(_01955_));
 sky130_fd_sc_hd__o21ba_1 _22398_ (.A1(_01918_),
    .A2(_01955_),
    .B1_N(_01259_),
    .X(_01956_));
 sky130_fd_sc_hd__a221o_1 _22399_ (.A1(_01143_),
    .A2(_01259_),
    .B1(_01954_),
    .B2(net119),
    .C1(_01956_),
    .X(_01957_));
 sky130_fd_sc_hd__nand2_1 _22400_ (.A(_01217_),
    .B(_01917_),
    .Y(_01958_));
 sky130_fd_sc_hd__or2_1 _22401_ (.A(_01217_),
    .B(_01917_),
    .X(_01959_));
 sky130_fd_sc_hd__and2b_1 _22402_ (.A_N(_01259_),
    .B(_01954_),
    .X(_01960_));
 sky130_fd_sc_hd__a41o_1 _22403_ (.A1(\top0.cordic0.vec[1][10] ),
    .A2(_01259_),
    .A3(_01958_),
    .A4(_01959_),
    .B1(_01960_),
    .X(_01961_));
 sky130_fd_sc_hd__a21oi_1 _22404_ (.A1(net134),
    .A2(_01957_),
    .B1(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__nor2_1 _22405_ (.A(_01065_),
    .B(net110),
    .Y(_01963_));
 sky130_fd_sc_hd__o21a_1 _22406_ (.A1(_01112_),
    .A2(_01963_),
    .B1(net127),
    .X(_01964_));
 sky130_fd_sc_hd__xnor2_1 _22407_ (.A(_01408_),
    .B(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__xnor2_2 _22408_ (.A(_01771_),
    .B(_01965_),
    .Y(_01966_));
 sky130_fd_sc_hd__a211o_2 _22409_ (.A1(_01131_),
    .A2(_01759_),
    .B1(_01761_),
    .C1(_01762_),
    .X(_01967_));
 sky130_fd_sc_hd__o21a_1 _22410_ (.A1(net80),
    .A2(net94),
    .B1(net89),
    .X(_01968_));
 sky130_fd_sc_hd__xnor2_2 _22411_ (.A(_01967_),
    .B(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__xnor2_1 _22412_ (.A(_01966_),
    .B(_01969_),
    .Y(_01970_));
 sky130_fd_sc_hd__xnor2_1 _22413_ (.A(_01962_),
    .B(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__mux2_1 _22414_ (.A0(net86),
    .A1(net80),
    .S(_01923_),
    .X(_01972_));
 sky130_fd_sc_hd__inv_2 _22415_ (.A(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__a221o_1 _22416_ (.A1(net97),
    .A2(_01230_),
    .B1(_01779_),
    .B2(_01922_),
    .C1(_11674_),
    .X(_01974_));
 sky130_fd_sc_hd__or3b_1 _22417_ (.A(net80),
    .B(_01923_),
    .C_N(_01925_),
    .X(_01975_));
 sky130_fd_sc_hd__o211a_1 _22418_ (.A1(net93),
    .A2(_01973_),
    .B1(_01974_),
    .C1(_01975_),
    .X(_01976_));
 sky130_fd_sc_hd__xnor2_1 _22419_ (.A(_01971_),
    .B(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__xnor2_2 _22420_ (.A(_01953_),
    .B(_01977_),
    .Y(_01978_));
 sky130_fd_sc_hd__a21oi_2 _22421_ (.A1(_01899_),
    .A2(_01932_),
    .B1(_01931_),
    .Y(_01979_));
 sky130_fd_sc_hd__nand2_2 _22422_ (.A(net79),
    .B(net87),
    .Y(_01980_));
 sky130_fd_sc_hd__o2bb2a_1 _22423_ (.A1_N(net95),
    .A2_N(_01902_),
    .B1(_01845_),
    .B2(net91),
    .X(_01981_));
 sky130_fd_sc_hd__or2_2 _22424_ (.A(_01980_),
    .B(_01981_),
    .X(_01982_));
 sky130_fd_sc_hd__xor2_1 _22425_ (.A(_01979_),
    .B(_01982_),
    .X(_01983_));
 sky130_fd_sc_hd__xnor2_1 _22426_ (.A(_01978_),
    .B(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__nor2_1 _22427_ (.A(_01951_),
    .B(_01984_),
    .Y(_01985_));
 sky130_fd_sc_hd__nand2_1 _22428_ (.A(_01951_),
    .B(_01984_),
    .Y(_01986_));
 sky130_fd_sc_hd__or2b_1 _22429_ (.A(_01985_),
    .B_N(_01986_),
    .X(_01987_));
 sky130_fd_sc_hd__inv_2 _22430_ (.A(_01942_),
    .Y(_01988_));
 sky130_fd_sc_hd__nand2_1 _22431_ (.A(_01896_),
    .B(_01988_),
    .Y(_01989_));
 sky130_fd_sc_hd__nand2_1 _22432_ (.A(_01885_),
    .B(_01941_),
    .Y(_01990_));
 sky130_fd_sc_hd__o21ai_1 _22433_ (.A1(_01885_),
    .A2(_01941_),
    .B1(_01898_),
    .Y(_01991_));
 sky130_fd_sc_hd__a21oi_1 _22434_ (.A1(_01990_),
    .A2(_01991_),
    .B1(_01896_),
    .Y(_01992_));
 sky130_fd_sc_hd__a311o_1 _22435_ (.A1(_01885_),
    .A2(_01898_),
    .A3(_01941_),
    .B1(_01992_),
    .C1(_01877_),
    .X(_01993_));
 sky130_fd_sc_hd__a211o_1 _22436_ (.A1(_01896_),
    .A2(_01943_),
    .B1(_01988_),
    .C1(net210),
    .X(_01994_));
 sky130_fd_sc_hd__a2bb2o_1 _22437_ (.A1_N(_01885_),
    .A2_N(_01989_),
    .B1(_01993_),
    .B2(_01994_),
    .X(_01995_));
 sky130_fd_sc_hd__xnor2_1 _22438_ (.A(_01987_),
    .B(_01995_),
    .Y(_01996_));
 sky130_fd_sc_hd__nor2_1 _22439_ (.A(_12036_),
    .B(_01996_),
    .Y(_01997_));
 sky130_fd_sc_hd__a31o_1 _22440_ (.A1(net727),
    .A2(_12004_),
    .A3(_12740_),
    .B1(_01997_),
    .X(_00401_));
 sky130_fd_sc_hd__nor2_1 _22441_ (.A(_01944_),
    .B(_01987_),
    .Y(_01998_));
 sky130_fd_sc_hd__and3_1 _22442_ (.A(_01809_),
    .B(_01891_),
    .C(_01998_),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_1 _22443_ (.A0(_01943_),
    .A1(_01942_),
    .S(_01987_),
    .X(_02000_));
 sky130_fd_sc_hd__a21oi_1 _22444_ (.A1(_01809_),
    .A2(_01891_),
    .B1(_02000_),
    .Y(_02001_));
 sky130_fd_sc_hd__mux2_1 _22445_ (.A0(_01998_),
    .A1(_02001_),
    .S(_01895_),
    .X(_02002_));
 sky130_fd_sc_hd__o21ba_2 _22446_ (.A1(_01999_),
    .A2(_02002_),
    .B1_N(_01885_),
    .X(_02003_));
 sky130_fd_sc_hd__nand3b_1 _22447_ (.A_N(_01944_),
    .B(_01891_),
    .C(_01737_),
    .Y(_02004_));
 sky130_fd_sc_hd__a31o_1 _22448_ (.A1(_01258_),
    .A2(_01683_),
    .A3(_01738_),
    .B1(_02004_),
    .X(_02005_));
 sky130_fd_sc_hd__a21o_1 _22449_ (.A1(_01895_),
    .A2(_01943_),
    .B1(_01988_),
    .X(_02006_));
 sky130_fd_sc_hd__a31o_2 _22450_ (.A1(_01986_),
    .A2(_02005_),
    .A3(_02006_),
    .B1(_01985_),
    .X(_02007_));
 sky130_fd_sc_hd__a21o_1 _22451_ (.A1(_01979_),
    .A2(_01982_),
    .B1(_01978_),
    .X(_02008_));
 sky130_fd_sc_hd__o21ai_2 _22452_ (.A1(_01979_),
    .A2(_01982_),
    .B1(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__a21bo_1 _22453_ (.A1(_01966_),
    .A2(_01969_),
    .B1_N(_01962_),
    .X(_02010_));
 sky130_fd_sc_hd__o21ai_2 _22454_ (.A1(_01966_),
    .A2(_01969_),
    .B1(_02010_),
    .Y(_02011_));
 sky130_fd_sc_hd__mux2_1 _22455_ (.A0(_01292_),
    .A1(net114),
    .S(_01770_),
    .X(_02012_));
 sky130_fd_sc_hd__and3b_1 _22456_ (.A_N(_01770_),
    .B(_01065_),
    .C(_01135_),
    .X(_02013_));
 sky130_fd_sc_hd__a211o_1 _22457_ (.A1(_01135_),
    .A2(_01292_),
    .B1(_02012_),
    .C1(_02013_),
    .X(_02014_));
 sky130_fd_sc_hd__o21ba_1 _22458_ (.A1(_01292_),
    .A2(_01770_),
    .B1_N(_01287_),
    .X(_02015_));
 sky130_fd_sc_hd__a211o_1 _22459_ (.A1(_01292_),
    .A2(_01770_),
    .B1(_02015_),
    .C1(net109),
    .X(_02016_));
 sky130_fd_sc_hd__a21bo_2 _22460_ (.A1(net109),
    .A2(_02014_),
    .B1_N(_02016_),
    .X(_02017_));
 sky130_fd_sc_hd__nand2_1 _22461_ (.A(net111),
    .B(_01211_),
    .Y(_02018_));
 sky130_fd_sc_hd__mux2_1 _22462_ (.A0(_01224_),
    .A1(_02018_),
    .S(net125),
    .X(_02019_));
 sky130_fd_sc_hd__xnor2_2 _22463_ (.A(net88),
    .B(_01775_),
    .Y(_02020_));
 sky130_fd_sc_hd__xnor2_1 _22464_ (.A(_01312_),
    .B(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__xnor2_2 _22465_ (.A(_02019_),
    .B(_02021_),
    .Y(_02022_));
 sky130_fd_sc_hd__inv_2 _22466_ (.A(_01852_),
    .Y(_02023_));
 sky130_fd_sc_hd__o21a_1 _22467_ (.A1(_01643_),
    .A2(net92),
    .B1(_01119_),
    .X(_02024_));
 sky130_fd_sc_hd__a211o_1 _22468_ (.A1(net92),
    .A2(_01769_),
    .B1(_02023_),
    .C1(_02024_),
    .X(_02025_));
 sky130_fd_sc_hd__nand2_1 _22469_ (.A(net85),
    .B(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__or2_1 _22470_ (.A(net85),
    .B(_02025_),
    .X(_02027_));
 sky130_fd_sc_hd__and2_1 _22471_ (.A(_02026_),
    .B(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__xnor2_1 _22472_ (.A(_02022_),
    .B(_02028_),
    .Y(_02029_));
 sky130_fd_sc_hd__xnor2_2 _22473_ (.A(_02017_),
    .B(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__nor2_1 _22474_ (.A(net79),
    .B(_01166_),
    .Y(_02031_));
 sky130_fd_sc_hd__nor2_1 _22475_ (.A(_01230_),
    .B(_01967_),
    .Y(_02032_));
 sky130_fd_sc_hd__mux2_1 _22476_ (.A0(net80),
    .A1(_02031_),
    .S(_02032_),
    .X(_02033_));
 sky130_fd_sc_hd__inv_2 _22477_ (.A(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__xnor2_1 _22478_ (.A(_02030_),
    .B(_02034_),
    .Y(_02035_));
 sky130_fd_sc_hd__xnor2_2 _22479_ (.A(_02011_),
    .B(_02035_),
    .Y(_02036_));
 sky130_fd_sc_hd__a21o_1 _22480_ (.A1(_01953_),
    .A2(_01976_),
    .B1(_01971_),
    .X(_02037_));
 sky130_fd_sc_hd__o21a_1 _22481_ (.A1(_01953_),
    .A2(_01976_),
    .B1(_02037_),
    .X(_02038_));
 sky130_fd_sc_hd__nor2_1 _22482_ (.A(_01924_),
    .B(_01923_),
    .Y(_02039_));
 sky130_fd_sc_hd__o21ai_1 _22483_ (.A1(_01925_),
    .A2(_02039_),
    .B1(net80),
    .Y(_02040_));
 sky130_fd_sc_hd__nor2_1 _22484_ (.A(_02038_),
    .B(_02040_),
    .Y(_02041_));
 sky130_fd_sc_hd__nand2_1 _22485_ (.A(_02038_),
    .B(_02040_),
    .Y(_02042_));
 sky130_fd_sc_hd__and2b_1 _22486_ (.A_N(_02041_),
    .B(_02042_),
    .X(_02043_));
 sky130_fd_sc_hd__xnor2_2 _22487_ (.A(_02036_),
    .B(_02043_),
    .Y(_02044_));
 sky130_fd_sc_hd__xnor2_1 _22488_ (.A(_02009_),
    .B(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__xnor2_1 _22489_ (.A(_02007_),
    .B(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__o21ai_1 _22490_ (.A1(_01877_),
    .A2(_02003_),
    .B1(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__or3_1 _22491_ (.A(_01877_),
    .B(_02003_),
    .C(_02046_),
    .X(_02048_));
 sky130_fd_sc_hd__and3_1 _22492_ (.A(\top0.cordic0.sin[5] ),
    .B(_12004_),
    .C(_12035_),
    .X(_02049_));
 sky130_fd_sc_hd__a31o_1 _22493_ (.A1(_12742_),
    .A2(_02047_),
    .A3(_02048_),
    .B1(_02049_),
    .X(_00402_));
 sky130_fd_sc_hd__o21a_1 _22494_ (.A1(_02030_),
    .A2(_02034_),
    .B1(_02011_),
    .X(_02050_));
 sky130_fd_sc_hd__a21o_1 _22495_ (.A1(_02030_),
    .A2(_02034_),
    .B1(_02050_),
    .X(_02051_));
 sky130_fd_sc_hd__o21a_1 _22496_ (.A1(_02017_),
    .A2(_02022_),
    .B1(_02028_),
    .X(_02052_));
 sky130_fd_sc_hd__a21o_1 _22497_ (.A1(_02017_),
    .A2(_02022_),
    .B1(_02052_),
    .X(_02053_));
 sky130_fd_sc_hd__xnor2_1 _22498_ (.A(net112),
    .B(_02020_),
    .Y(_02054_));
 sky130_fd_sc_hd__nor3_1 _22499_ (.A(net107),
    .B(_01312_),
    .C(_02020_),
    .Y(_02055_));
 sky130_fd_sc_hd__or3_1 _22500_ (.A(_01213_),
    .B(net107),
    .C(_02020_),
    .X(_02056_));
 sky130_fd_sc_hd__o21a_1 _22501_ (.A1(net111),
    .A2(_02020_),
    .B1(_02018_),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_1 _22502_ (.A0(_02057_),
    .A1(_01224_),
    .S(_01312_),
    .X(_02058_));
 sky130_fd_sc_hd__a21oi_1 _22503_ (.A1(_02056_),
    .A2(_02058_),
    .B1(_01408_),
    .Y(_02059_));
 sky130_fd_sc_hd__a311o_2 _22504_ (.A1(net107),
    .A2(_01312_),
    .A3(_02054_),
    .B1(_02055_),
    .C1(_02059_),
    .X(_02060_));
 sky130_fd_sc_hd__xor2_4 _22505_ (.A(_01069_),
    .B(_01924_),
    .X(_02061_));
 sky130_fd_sc_hd__and3_1 _22506_ (.A(net119),
    .B(net104),
    .C(_01643_),
    .X(_02062_));
 sky130_fd_sc_hd__a21oi_2 _22507_ (.A1(_01217_),
    .A2(_01784_),
    .B1(_02062_),
    .Y(_02063_));
 sky130_fd_sc_hd__xnor2_4 _22508_ (.A(_02061_),
    .B(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__nor2_1 _22509_ (.A(_01230_),
    .B(_01775_),
    .Y(_02065_));
 sky130_fd_sc_hd__a22o_1 _22510_ (.A1(net111),
    .A2(net107),
    .B1(net98),
    .B2(_01230_),
    .X(_02066_));
 sky130_fd_sc_hd__o21ai_4 _22511_ (.A1(_01821_),
    .A2(_02065_),
    .B1(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__xor2_2 _22512_ (.A(_02064_),
    .B(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__xor2_2 _22513_ (.A(_02060_),
    .B(_02068_),
    .X(_02069_));
 sky130_fd_sc_hd__xnor2_1 _22514_ (.A(_02026_),
    .B(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__xnor2_1 _22515_ (.A(_02053_),
    .B(_02070_),
    .Y(_02071_));
 sky130_fd_sc_hd__nor2_1 _22516_ (.A(_01980_),
    .B(_01967_),
    .Y(_02072_));
 sky130_fd_sc_hd__nand2_1 _22517_ (.A(_02071_),
    .B(_02072_),
    .Y(_02073_));
 sky130_fd_sc_hd__nor2_1 _22518_ (.A(_02071_),
    .B(_02072_),
    .Y(_02074_));
 sky130_fd_sc_hd__inv_2 _22519_ (.A(_02074_),
    .Y(_02075_));
 sky130_fd_sc_hd__nand2_1 _22520_ (.A(_02073_),
    .B(_02075_),
    .Y(_02076_));
 sky130_fd_sc_hd__xnor2_2 _22521_ (.A(_02051_),
    .B(_02076_),
    .Y(_02077_));
 sky130_fd_sc_hd__o21ai_1 _22522_ (.A1(_02038_),
    .A2(_02040_),
    .B1(_02036_),
    .Y(_02078_));
 sky130_fd_sc_hd__nand2_2 _22523_ (.A(_02042_),
    .B(_02078_),
    .Y(_02079_));
 sky130_fd_sc_hd__nand2_1 _22524_ (.A(_02077_),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__nor2_1 _22525_ (.A(_02077_),
    .B(_02079_),
    .Y(_02081_));
 sky130_fd_sc_hd__inv_2 _22526_ (.A(_02081_),
    .Y(_02082_));
 sky130_fd_sc_hd__nand2_1 _22527_ (.A(_02080_),
    .B(_02082_),
    .Y(_02083_));
 sky130_fd_sc_hd__nor2_2 _22528_ (.A(_02009_),
    .B(_02044_),
    .Y(_02084_));
 sky130_fd_sc_hd__nand2_1 _22529_ (.A(_02009_),
    .B(_02044_),
    .Y(_02085_));
 sky130_fd_sc_hd__a21o_1 _22530_ (.A1(_02007_),
    .A2(_02085_),
    .B1(_02084_),
    .X(_02086_));
 sky130_fd_sc_hd__o21a_1 _22531_ (.A1(_02003_),
    .A2(_02084_),
    .B1(_02085_),
    .X(_02087_));
 sky130_fd_sc_hd__o221a_1 _22532_ (.A1(_02003_),
    .A2(_02085_),
    .B1(_02087_),
    .B2(_02007_),
    .C1(net210),
    .X(_02088_));
 sky130_fd_sc_hd__o21ba_1 _22533_ (.A1(net210),
    .A2(_02086_),
    .B1_N(_02088_),
    .X(_02089_));
 sky130_fd_sc_hd__a31o_1 _22534_ (.A1(_02003_),
    .A2(_02007_),
    .A3(_02084_),
    .B1(_02089_),
    .X(_02090_));
 sky130_fd_sc_hd__xnor2_1 _22535_ (.A(_02083_),
    .B(_02090_),
    .Y(_02091_));
 sky130_fd_sc_hd__nor2_1 _22536_ (.A(_12036_),
    .B(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__a31o_1 _22537_ (.A1(net726),
    .A2(_12004_),
    .A3(_12740_),
    .B1(_02092_),
    .X(_00403_));
 sky130_fd_sc_hd__o211a_1 _22538_ (.A1(_02007_),
    .A2(_02084_),
    .B1(_02085_),
    .C1(_02082_),
    .X(_02093_));
 sky130_fd_sc_hd__a21oi_1 _22539_ (.A1(_02077_),
    .A2(_02079_),
    .B1(_02093_),
    .Y(_02094_));
 sky130_fd_sc_hd__inv_2 _22540_ (.A(_02053_),
    .Y(_02095_));
 sky130_fd_sc_hd__nor2_1 _22541_ (.A(_02095_),
    .B(_02069_),
    .Y(_02096_));
 sky130_fd_sc_hd__nand2_1 _22542_ (.A(_02095_),
    .B(_02069_),
    .Y(_02097_));
 sky130_fd_sc_hd__o21ai_2 _22543_ (.A1(_02026_),
    .A2(_02096_),
    .B1(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__nor2_1 _22544_ (.A(_02064_),
    .B(_02067_),
    .Y(_02099_));
 sky130_fd_sc_hd__and3_1 _22545_ (.A(net79),
    .B(_02064_),
    .C(_02067_),
    .X(_02100_));
 sky130_fd_sc_hd__a221o_2 _22546_ (.A1(_02060_),
    .A2(_02068_),
    .B1(_02099_),
    .B2(_01948_),
    .C1(_02100_),
    .X(_02101_));
 sky130_fd_sc_hd__xnor2_1 _22547_ (.A(net77),
    .B(_01924_),
    .Y(_02102_));
 sky130_fd_sc_hd__o211ai_1 _22548_ (.A1(net119),
    .A2(net104),
    .B1(_01069_),
    .C1(_02102_),
    .Y(_02103_));
 sky130_fd_sc_hd__nor2_1 _22549_ (.A(net119),
    .B(_01069_),
    .Y(_02104_));
 sky130_fd_sc_hd__or3_1 _22550_ (.A(net104),
    .B(_02102_),
    .C(_02104_),
    .X(_02105_));
 sky130_fd_sc_hd__a21o_1 _22551_ (.A1(_01069_),
    .A2(_01616_),
    .B1(_02102_),
    .X(_02106_));
 sky130_fd_sc_hd__o211a_1 _22552_ (.A1(_01069_),
    .A2(_01616_),
    .B1(_02106_),
    .C1(_01643_),
    .X(_02107_));
 sky130_fd_sc_hd__a31o_2 _22553_ (.A1(net102),
    .A2(_02103_),
    .A3(_02105_),
    .B1(_02107_),
    .X(_02108_));
 sky130_fd_sc_hd__xnor2_1 _22554_ (.A(_01074_),
    .B(_01980_),
    .Y(_02109_));
 sky130_fd_sc_hd__mux2_1 _22555_ (.A0(_01769_),
    .A1(_01798_),
    .S(net115),
    .X(_02110_));
 sky130_fd_sc_hd__xnor2_2 _22556_ (.A(_02109_),
    .B(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__nand2_1 _22557_ (.A(net107),
    .B(net101),
    .Y(_02112_));
 sky130_fd_sc_hd__and3_1 _22558_ (.A(net107),
    .B(net100),
    .C(_01924_),
    .X(_02113_));
 sky130_fd_sc_hd__a221o_1 _22559_ (.A1(net89),
    .A2(_02031_),
    .B1(_02112_),
    .B2(net79),
    .C1(_02113_),
    .X(_02114_));
 sky130_fd_sc_hd__xor2_1 _22560_ (.A(_02111_),
    .B(_02114_),
    .X(_02115_));
 sky130_fd_sc_hd__xnor2_2 _22561_ (.A(_02108_),
    .B(_02115_),
    .Y(_02116_));
 sky130_fd_sc_hd__nand2_1 _22562_ (.A(net80),
    .B(_02067_),
    .Y(_02117_));
 sky130_fd_sc_hd__xor2_1 _22563_ (.A(_02116_),
    .B(_02117_),
    .X(_02118_));
 sky130_fd_sc_hd__xnor2_2 _22564_ (.A(_02101_),
    .B(_02118_),
    .Y(_02119_));
 sky130_fd_sc_hd__nor2_1 _22565_ (.A(_01948_),
    .B(_02025_),
    .Y(_02120_));
 sky130_fd_sc_hd__xnor2_1 _22566_ (.A(_02119_),
    .B(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__xnor2_1 _22567_ (.A(_02098_),
    .B(_02121_),
    .Y(_02122_));
 sky130_fd_sc_hd__a21oi_2 _22568_ (.A1(_02051_),
    .A2(_02073_),
    .B1(_02074_),
    .Y(_02123_));
 sky130_fd_sc_hd__nand2_1 _22569_ (.A(_02122_),
    .B(_02123_),
    .Y(_02124_));
 sky130_fd_sc_hd__or2_1 _22570_ (.A(_02122_),
    .B(_02123_),
    .X(_02125_));
 sky130_fd_sc_hd__and2_1 _22571_ (.A(_02124_),
    .B(_02125_),
    .X(_02126_));
 sky130_fd_sc_hd__xnor2_1 _22572_ (.A(_02094_),
    .B(_02126_),
    .Y(_02127_));
 sky130_fd_sc_hd__mux2_1 _22573_ (.A0(_02045_),
    .A1(_02085_),
    .S(_02007_),
    .X(_02128_));
 sky130_fd_sc_hd__nand2_1 _22574_ (.A(_02007_),
    .B(_02084_),
    .Y(_02129_));
 sky130_fd_sc_hd__mux2_1 _22575_ (.A0(_02128_),
    .A1(_02129_),
    .S(_02083_),
    .X(_02130_));
 sky130_fd_sc_hd__or2b_1 _22576_ (.A(_02130_),
    .B_N(_02003_),
    .X(_02131_));
 sky130_fd_sc_hd__nand2_1 _22577_ (.A(net211),
    .B(_02131_),
    .Y(_02132_));
 sky130_fd_sc_hd__xor2_1 _22578_ (.A(_02127_),
    .B(_02132_),
    .X(_02133_));
 sky130_fd_sc_hd__a22o_1 _22579_ (.A1(net769),
    .A2(_12813_),
    .B1(_02133_),
    .B2(_12963_),
    .X(_00404_));
 sky130_fd_sc_hd__inv_2 _22580_ (.A(_02123_),
    .Y(_02134_));
 sky130_fd_sc_hd__a22o_1 _22581_ (.A1(_02079_),
    .A2(_02134_),
    .B1(_02124_),
    .B2(_02086_),
    .X(_02135_));
 sky130_fd_sc_hd__a21oi_1 _22582_ (.A1(_02080_),
    .A2(_02123_),
    .B1(_02122_),
    .Y(_02136_));
 sky130_fd_sc_hd__a31o_1 _22583_ (.A1(_02079_),
    .A2(_02086_),
    .A3(_02124_),
    .B1(_02136_),
    .X(_02137_));
 sky130_fd_sc_hd__a21oi_2 _22584_ (.A1(_02077_),
    .A2(_02135_),
    .B1(_02137_),
    .Y(_02138_));
 sky130_fd_sc_hd__a21bo_1 _22585_ (.A1(_02101_),
    .A2(_02116_),
    .B1_N(_02117_),
    .X(_02139_));
 sky130_fd_sc_hd__o21a_2 _22586_ (.A1(_02101_),
    .A2(_02116_),
    .B1(_02139_),
    .X(_02140_));
 sky130_fd_sc_hd__a21bo_1 _22587_ (.A1(_02111_),
    .A2(_02114_),
    .B1_N(_02108_),
    .X(_02141_));
 sky130_fd_sc_hd__o21a_1 _22588_ (.A1(_02111_),
    .A2(_02114_),
    .B1(_02141_),
    .X(_02142_));
 sky130_fd_sc_hd__inv_2 _22589_ (.A(_02142_),
    .Y(_02143_));
 sky130_fd_sc_hd__or2_1 _22590_ (.A(_02112_),
    .B(_01924_),
    .X(_02144_));
 sky130_fd_sc_hd__nand2_1 _22591_ (.A(net79),
    .B(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__nor2_1 _22592_ (.A(net95),
    .B(_01980_),
    .Y(_02146_));
 sky130_fd_sc_hd__nor2_1 _22593_ (.A(\top0.cordic0.vec[1][13] ),
    .B(_01980_),
    .Y(_02147_));
 sky130_fd_sc_hd__o21ba_1 _22594_ (.A1(_01798_),
    .A2(_02147_),
    .B1_N(_01074_),
    .X(_02148_));
 sky130_fd_sc_hd__a221o_1 _22595_ (.A1(_01074_),
    .A2(_01769_),
    .B1(_02146_),
    .B2(net100),
    .C1(_02148_),
    .X(_02149_));
 sky130_fd_sc_hd__and2_1 _22596_ (.A(net103),
    .B(_01980_),
    .X(_02150_));
 sky130_fd_sc_hd__o21a_1 _22597_ (.A1(_02147_),
    .A2(_02150_),
    .B1(net98),
    .X(_02151_));
 sky130_fd_sc_hd__mux2_1 _22598_ (.A0(_02146_),
    .A1(_02151_),
    .S(_01074_),
    .X(_02152_));
 sky130_fd_sc_hd__a21oi_2 _22599_ (.A1(net114),
    .A2(_02149_),
    .B1(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__a31o_1 _22600_ (.A1(net101),
    .A2(net97),
    .A3(net87),
    .B1(_11674_),
    .X(_02154_));
 sky130_fd_sc_hd__or3_1 _22601_ (.A(_01213_),
    .B(_01063_),
    .C(net92),
    .X(_02155_));
 sky130_fd_sc_hd__or3_1 _22602_ (.A(net112),
    .B(net95),
    .C(_01166_),
    .X(_02156_));
 sky130_fd_sc_hd__nand2_1 _22603_ (.A(_02155_),
    .B(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__xnor2_1 _22604_ (.A(net79),
    .B(_01115_),
    .Y(_02158_));
 sky130_fd_sc_hd__xnor2_1 _22605_ (.A(_02157_),
    .B(_02158_),
    .Y(_02159_));
 sky130_fd_sc_hd__or2b_1 _22606_ (.A(_02154_),
    .B_N(_02159_),
    .X(_02160_));
 sky130_fd_sc_hd__or2b_1 _22607_ (.A(_02159_),
    .B_N(_02154_),
    .X(_02161_));
 sky130_fd_sc_hd__nand2_1 _22608_ (.A(_02160_),
    .B(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hd__xor2_2 _22609_ (.A(_02153_),
    .B(_02162_),
    .X(_02163_));
 sky130_fd_sc_hd__xor2_1 _22610_ (.A(_02145_),
    .B(_02163_),
    .X(_02164_));
 sky130_fd_sc_hd__xnor2_2 _22611_ (.A(_02143_),
    .B(_02164_),
    .Y(_02165_));
 sky130_fd_sc_hd__or2_1 _22612_ (.A(_01948_),
    .B(_02067_),
    .X(_02166_));
 sky130_fd_sc_hd__xnor2_1 _22613_ (.A(_02165_),
    .B(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__xnor2_2 _22614_ (.A(_02140_),
    .B(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__a21o_1 _22615_ (.A1(_02098_),
    .A2(_02119_),
    .B1(_02120_),
    .X(_02169_));
 sky130_fd_sc_hd__o21ai_2 _22616_ (.A1(_02098_),
    .A2(_02119_),
    .B1(_02169_),
    .Y(_02170_));
 sky130_fd_sc_hd__nor2_2 _22617_ (.A(_02168_),
    .B(_02170_),
    .Y(_02171_));
 sky130_fd_sc_hd__inv_2 _22618_ (.A(_02171_),
    .Y(_02172_));
 sky130_fd_sc_hd__nand2_1 _22619_ (.A(_02168_),
    .B(_02170_),
    .Y(_02173_));
 sky130_fd_sc_hd__and2_1 _22620_ (.A(_02172_),
    .B(_02173_),
    .X(_02174_));
 sky130_fd_sc_hd__xor2_2 _22621_ (.A(_02138_),
    .B(_02174_),
    .X(_02175_));
 sky130_fd_sc_hd__nand3b_1 _22622_ (.A_N(_02130_),
    .B(_02127_),
    .C(_02003_),
    .Y(_02176_));
 sky130_fd_sc_hd__or3b_1 _22623_ (.A(_01877_),
    .B(_02175_),
    .C_N(_02176_),
    .X(_02177_));
 sky130_fd_sc_hd__a21bo_1 _22624_ (.A1(net211),
    .A2(_02176_),
    .B1_N(_02175_),
    .X(_02178_));
 sky130_fd_sc_hd__a21oi_1 _22625_ (.A1(_02177_),
    .A2(_02178_),
    .B1(_12740_),
    .Y(_02179_));
 sky130_fd_sc_hd__a31o_1 _22626_ (.A1(net724),
    .A2(_12004_),
    .A3(_12740_),
    .B1(_02179_),
    .X(_00405_));
 sky130_fd_sc_hd__or2_2 _22627_ (.A(_02175_),
    .B(_02176_),
    .X(_02180_));
 sky130_fd_sc_hd__nand2_1 _22628_ (.A(net211),
    .B(_02180_),
    .Y(_02181_));
 sky130_fd_sc_hd__or2b_1 _22629_ (.A(_02094_),
    .B_N(_02124_),
    .X(_02182_));
 sky130_fd_sc_hd__and2_1 _22630_ (.A(_02125_),
    .B(_02173_),
    .X(_02183_));
 sky130_fd_sc_hd__a21o_1 _22631_ (.A1(_02182_),
    .A2(_02183_),
    .B1(_02171_),
    .X(_02184_));
 sky130_fd_sc_hd__a21bo_1 _22632_ (.A1(_02140_),
    .A2(_02165_),
    .B1_N(_02166_),
    .X(_02185_));
 sky130_fd_sc_hd__o21ai_2 _22633_ (.A1(_02140_),
    .A2(_02165_),
    .B1(_02185_),
    .Y(_02186_));
 sky130_fd_sc_hd__a21o_1 _22634_ (.A1(_01213_),
    .A2(_01063_),
    .B1(net78),
    .X(_02187_));
 sky130_fd_sc_hd__a211o_1 _22635_ (.A1(_01221_),
    .A2(_02187_),
    .B1(_01166_),
    .C1(_01118_),
    .X(_02188_));
 sky130_fd_sc_hd__a21o_1 _22636_ (.A1(_01063_),
    .A2(_01118_),
    .B1(_01776_),
    .X(_02189_));
 sky130_fd_sc_hd__a22o_1 _22637_ (.A1(_01118_),
    .A2(_01776_),
    .B1(_02189_),
    .B2(net77),
    .X(_02190_));
 sky130_fd_sc_hd__nand2_1 _22638_ (.A(net110),
    .B(_02190_),
    .Y(_02191_));
 sky130_fd_sc_hd__o311a_2 _22639_ (.A1(_11674_),
    .A2(net93),
    .A3(_01115_),
    .B1(_02188_),
    .C1(_02191_),
    .X(_02192_));
 sky130_fd_sc_hd__mux2_1 _22640_ (.A0(_01924_),
    .A1(_01821_),
    .S(net107),
    .X(_02193_));
 sky130_fd_sc_hd__xnor2_2 _22641_ (.A(_01643_),
    .B(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__nand2_1 _22642_ (.A(net79),
    .B(_01248_),
    .Y(_02195_));
 sky130_fd_sc_hd__or2_1 _22643_ (.A(_02194_),
    .B(_02195_),
    .X(_02196_));
 sky130_fd_sc_hd__nand2_1 _22644_ (.A(_02194_),
    .B(_02195_),
    .Y(_02197_));
 sky130_fd_sc_hd__and2_1 _22645_ (.A(_02196_),
    .B(_02197_),
    .X(_02198_));
 sky130_fd_sc_hd__xnor2_2 _22646_ (.A(_02192_),
    .B(_02198_),
    .Y(_02199_));
 sky130_fd_sc_hd__mux2_1 _22647_ (.A0(_02161_),
    .A1(_02160_),
    .S(_02153_),
    .X(_02200_));
 sky130_fd_sc_hd__xor2_1 _22648_ (.A(_02199_),
    .B(_02200_),
    .X(_02201_));
 sky130_fd_sc_hd__inv_2 _22649_ (.A(_02201_),
    .Y(_02202_));
 sky130_fd_sc_hd__o21a_1 _22650_ (.A1(_02143_),
    .A2(_02163_),
    .B1(_01948_),
    .X(_02203_));
 sky130_fd_sc_hd__a31o_1 _22651_ (.A1(_02144_),
    .A2(_02143_),
    .A3(_02163_),
    .B1(_02203_),
    .X(_02204_));
 sky130_fd_sc_hd__and2_1 _22652_ (.A(_02202_),
    .B(_02204_),
    .X(_02205_));
 sky130_fd_sc_hd__nor2_1 _22653_ (.A(_02202_),
    .B(_02204_),
    .Y(_02206_));
 sky130_fd_sc_hd__or2_2 _22654_ (.A(_02205_),
    .B(_02206_),
    .X(_02207_));
 sky130_fd_sc_hd__or2_1 _22655_ (.A(_02186_),
    .B(_02207_),
    .X(_02208_));
 sky130_fd_sc_hd__nand2_1 _22656_ (.A(_02186_),
    .B(_02207_),
    .Y(_02209_));
 sky130_fd_sc_hd__nand2_1 _22657_ (.A(_02208_),
    .B(_02209_),
    .Y(_02210_));
 sky130_fd_sc_hd__xnor2_1 _22658_ (.A(_02184_),
    .B(_02210_),
    .Y(_02211_));
 sky130_fd_sc_hd__xnor2_1 _22659_ (.A(_02181_),
    .B(_02211_),
    .Y(_02212_));
 sky130_fd_sc_hd__a22o_1 _22660_ (.A1(net720),
    .A2(_12813_),
    .B1(_02212_),
    .B2(_12742_),
    .X(_00406_));
 sky130_fd_sc_hd__a21o_1 _22661_ (.A1(_02159_),
    .A2(_02199_),
    .B1(_02154_),
    .X(_02213_));
 sky130_fd_sc_hd__or2_1 _22662_ (.A(_02159_),
    .B(_02199_),
    .X(_02214_));
 sky130_fd_sc_hd__a22o_1 _22663_ (.A1(_02153_),
    .A2(_02213_),
    .B1(_02214_),
    .B2(_02154_),
    .X(_02215_));
 sky130_fd_sc_hd__o21ai_1 _22664_ (.A1(net101),
    .A2(net90),
    .B1(net86),
    .Y(_02216_));
 sky130_fd_sc_hd__nand2_1 _22665_ (.A(net99),
    .B(net90),
    .Y(_02217_));
 sky130_fd_sc_hd__a22o_1 _22666_ (.A1(_01211_),
    .A2(_02216_),
    .B1(_02217_),
    .B2(_01230_),
    .X(_02218_));
 sky130_fd_sc_hd__xnor2_2 _22667_ (.A(_01223_),
    .B(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__mux2_1 _22668_ (.A0(_02197_),
    .A1(_02196_),
    .S(_02192_),
    .X(_02220_));
 sky130_fd_sc_hd__xor2_1 _22669_ (.A(_02219_),
    .B(_02220_),
    .X(_02221_));
 sky130_fd_sc_hd__o32a_1 _22670_ (.A1(_01643_),
    .A2(_01063_),
    .A3(_01980_),
    .B1(_02215_),
    .B2(_02221_),
    .X(_02222_));
 sky130_fd_sc_hd__a21boi_2 _22671_ (.A1(_02215_),
    .A2(_02221_),
    .B1_N(_02222_),
    .Y(_02223_));
 sky130_fd_sc_hd__xnor2_2 _22672_ (.A(_02206_),
    .B(_02223_),
    .Y(_02224_));
 sky130_fd_sc_hd__inv_2 _22673_ (.A(_02207_),
    .Y(_02225_));
 sky130_fd_sc_hd__o31a_1 _22674_ (.A1(_02175_),
    .A2(_02176_),
    .A3(_02225_),
    .B1(_02184_),
    .X(_02226_));
 sky130_fd_sc_hd__a21oi_1 _22675_ (.A1(_02180_),
    .A2(_02225_),
    .B1(_02226_),
    .Y(_02227_));
 sky130_fd_sc_hd__a21oi_1 _22676_ (.A1(_02182_),
    .A2(_02183_),
    .B1(_02171_),
    .Y(_02228_));
 sky130_fd_sc_hd__or3b_1 _22677_ (.A(_02207_),
    .B(_02228_),
    .C_N(_02180_),
    .X(_02229_));
 sky130_fd_sc_hd__o211a_1 _22678_ (.A1(_02186_),
    .A2(_02227_),
    .B1(_02229_),
    .C1(net210),
    .X(_02230_));
 sky130_fd_sc_hd__inv_2 _22679_ (.A(_02209_),
    .Y(_02231_));
 sky130_fd_sc_hd__a211oi_1 _22680_ (.A1(_02228_),
    .A2(_02208_),
    .B1(_02231_),
    .C1(net210),
    .Y(_02232_));
 sky130_fd_sc_hd__o32a_1 _22681_ (.A1(_02180_),
    .A2(_02184_),
    .A3(_02209_),
    .B1(_02230_),
    .B2(_02232_),
    .X(_02233_));
 sky130_fd_sc_hd__xnor2_1 _22682_ (.A(_02224_),
    .B(_02233_),
    .Y(_02234_));
 sky130_fd_sc_hd__and3_1 _22683_ (.A(\top0.cordic0.sin[10] ),
    .B(_12004_),
    .C(_12036_),
    .X(_02235_));
 sky130_fd_sc_hd__a21o_1 _22684_ (.A1(_12963_),
    .A2(_02234_),
    .B1(_02235_),
    .X(_00407_));
 sky130_fd_sc_hd__o211a_1 _22685_ (.A1(_02138_),
    .A2(_02171_),
    .B1(_02173_),
    .C1(_02209_),
    .X(_02236_));
 sky130_fd_sc_hd__o21ai_1 _22686_ (.A1(_02223_),
    .A2(_02236_),
    .B1(_02206_),
    .Y(_02237_));
 sky130_fd_sc_hd__a221o_1 _22687_ (.A1(_02077_),
    .A2(_02135_),
    .B1(_02168_),
    .B2(_02170_),
    .C1(_02137_),
    .X(_02238_));
 sky130_fd_sc_hd__a21o_1 _22688_ (.A1(_02172_),
    .A2(_02238_),
    .B1(_02231_),
    .X(_02239_));
 sky130_fd_sc_hd__a21bo_1 _22689_ (.A1(_02208_),
    .A2(_02239_),
    .B1_N(_02223_),
    .X(_02240_));
 sky130_fd_sc_hd__nand2_1 _22690_ (.A(_02237_),
    .B(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__a22oi_1 _22691_ (.A1(net100),
    .A2(_01924_),
    .B1(_01821_),
    .B2(_01762_),
    .Y(_02242_));
 sky130_fd_sc_hd__a211o_1 _22692_ (.A1(net97),
    .A2(net87),
    .B1(net91),
    .C1(net79),
    .X(_02243_));
 sky130_fd_sc_hd__o32a_1 _22693_ (.A1(net78),
    .A2(net99),
    .A3(net91),
    .B1(_01221_),
    .B2(_01937_),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_1 _22694_ (.A0(net90),
    .A1(_01849_),
    .S(_01948_),
    .X(_02245_));
 sky130_fd_sc_hd__nor2_1 _22695_ (.A(_01643_),
    .B(_01248_),
    .Y(_02246_));
 sky130_fd_sc_hd__mux2_1 _22696_ (.A0(_01924_),
    .A1(_02246_),
    .S(_01948_),
    .X(_02247_));
 sky130_fd_sc_hd__nand2_1 _22697_ (.A(net104),
    .B(_02247_),
    .Y(_02248_));
 sky130_fd_sc_hd__o221a_1 _22698_ (.A1(net104),
    .A2(_02244_),
    .B1(_02245_),
    .B2(_01063_),
    .C1(_02248_),
    .X(_02249_));
 sky130_fd_sc_hd__o211a_1 _22699_ (.A1(_01948_),
    .A2(_02242_),
    .B1(_02243_),
    .C1(_02249_),
    .X(_02250_));
 sky130_fd_sc_hd__a21oi_1 _22700_ (.A1(_02194_),
    .A2(_02219_),
    .B1(net79),
    .Y(_02251_));
 sky130_fd_sc_hd__nor2_1 _22701_ (.A(_02194_),
    .B(_02219_),
    .Y(_02252_));
 sky130_fd_sc_hd__o22ai_2 _22702_ (.A1(_02192_),
    .A2(_02251_),
    .B1(_02252_),
    .B2(_02195_),
    .Y(_02253_));
 sky130_fd_sc_hd__o2bb2a_1 _22703_ (.A1_N(_02250_),
    .A2_N(_02253_),
    .B1(_01948_),
    .B2(_01248_),
    .X(_02254_));
 sky130_fd_sc_hd__o21ai_2 _22704_ (.A1(_02250_),
    .A2(_02253_),
    .B1(_02254_),
    .Y(_02255_));
 sky130_fd_sc_hd__xor2_1 _22705_ (.A(_02222_),
    .B(_02255_),
    .X(_02256_));
 sky130_fd_sc_hd__xnor2_1 _22706_ (.A(_02241_),
    .B(_02256_),
    .Y(_02257_));
 sky130_fd_sc_hd__nand2_1 _22707_ (.A(_02231_),
    .B(_02224_),
    .Y(_02258_));
 sky130_fd_sc_hd__or3_1 _22708_ (.A(_02186_),
    .B(_02207_),
    .C(_02224_),
    .X(_02259_));
 sky130_fd_sc_hd__a21o_1 _22709_ (.A1(_02258_),
    .A2(_02259_),
    .B1(_02171_),
    .X(_02260_));
 sky130_fd_sc_hd__or3b_1 _22710_ (.A(_02210_),
    .B(_02224_),
    .C_N(_02183_),
    .X(_02261_));
 sky130_fd_sc_hd__mux2_1 _22711_ (.A0(_02260_),
    .A1(_02261_),
    .S(_02182_),
    .X(_02262_));
 sky130_fd_sc_hd__o21a_1 _22712_ (.A1(_02125_),
    .A2(_02171_),
    .B1(_02173_),
    .X(_02263_));
 sky130_fd_sc_hd__o21a_1 _22713_ (.A1(_02186_),
    .A2(_02263_),
    .B1(_02172_),
    .X(_02264_));
 sky130_fd_sc_hd__or2_1 _22714_ (.A(_02258_),
    .B(_02263_),
    .X(_02265_));
 sky130_fd_sc_hd__o31a_1 _22715_ (.A1(_02207_),
    .A2(_02224_),
    .A3(_02264_),
    .B1(_02265_),
    .X(_02266_));
 sky130_fd_sc_hd__a21oi_1 _22716_ (.A1(_02262_),
    .A2(_02266_),
    .B1(_02180_),
    .Y(_02267_));
 sky130_fd_sc_hd__or2_1 _22717_ (.A(_01877_),
    .B(_02267_),
    .X(_02268_));
 sky130_fd_sc_hd__xnor2_1 _22718_ (.A(_02257_),
    .B(_02268_),
    .Y(_02269_));
 sky130_fd_sc_hd__nor2_1 _22719_ (.A(_12036_),
    .B(_02269_),
    .Y(_02270_));
 sky130_fd_sc_hd__a31o_1 _22720_ (.A1(net733),
    .A2(_12004_),
    .A3(_12740_),
    .B1(_02270_),
    .X(_00408_));
 sky130_fd_sc_hd__a21o_1 _22721_ (.A1(_02237_),
    .A2(_02240_),
    .B1(_02255_),
    .X(_02271_));
 sky130_fd_sc_hd__a22o_1 _22722_ (.A1(_02237_),
    .A2(_02255_),
    .B1(_02271_),
    .B2(_02222_),
    .X(_02272_));
 sky130_fd_sc_hd__o32a_1 _22723_ (.A1(net104),
    .A2(net100),
    .A3(_01852_),
    .B1(_01167_),
    .B2(net78),
    .X(_02273_));
 sky130_fd_sc_hd__o22a_1 _22724_ (.A1(_01248_),
    .A2(_02112_),
    .B1(_02023_),
    .B2(_01948_),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _22725_ (.A0(_02273_),
    .A1(_02274_),
    .S(_01230_),
    .X(_02275_));
 sky130_fd_sc_hd__xnor2_1 _22726_ (.A(_02254_),
    .B(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__xnor2_1 _22727_ (.A(_02272_),
    .B(_02276_),
    .Y(_02277_));
 sky130_fd_sc_hd__a21oi_1 _22728_ (.A1(_02257_),
    .A2(_02267_),
    .B1(_01877_),
    .Y(_02278_));
 sky130_fd_sc_hd__xnor2_1 _22729_ (.A(_02277_),
    .B(_02278_),
    .Y(_02279_));
 sky130_fd_sc_hd__and3_1 _22730_ (.A(\top0.cordic0.sin[12] ),
    .B(_12004_),
    .C(_12036_),
    .X(_02280_));
 sky130_fd_sc_hd__a21o_1 _22731_ (.A1(_12963_),
    .A2(_02279_),
    .B1(_02280_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _22732_ (.A0(_01877_),
    .A1(_02278_),
    .S(_02277_),
    .X(_02281_));
 sky130_fd_sc_hd__a22o_1 _22733_ (.A1(net740),
    .A2(_12813_),
    .B1(_02281_),
    .B2(_12742_),
    .X(_00410_));
 sky130_fd_sc_hd__o21a_1 _22734_ (.A1(net915),
    .A2(_11431_),
    .B1(net178),
    .X(_00411_));
 sky130_fd_sc_hd__clkbuf_4 _22735_ (.A(_08900_),
    .X(_02282_));
 sky130_fd_sc_hd__nor2_1 _22736_ (.A(_02282_),
    .B(_12012_),
    .Y(_02283_));
 sky130_fd_sc_hd__o2bb2a_1 _22737_ (.A1_N(\top0.state[1] ),
    .A2_N(net206),
    .B1(\top0.start_svm ),
    .B2(_02283_),
    .X(_00412_));
 sky130_fd_sc_hd__nor2_1 _22738_ (.A(net197),
    .B(_11526_),
    .Y(_02284_));
 sky130_fd_sc_hd__mux2_1 _22739_ (.A0(net197),
    .A1(_02284_),
    .S(net174),
    .X(_02285_));
 sky130_fd_sc_hd__clkbuf_1 _22740_ (.A(_02285_),
    .X(_00413_));
 sky130_fd_sc_hd__nand2_1 _22741_ (.A(net174),
    .B(net197),
    .Y(_02286_));
 sky130_fd_sc_hd__xnor2_1 _22742_ (.A(net191),
    .B(_02286_),
    .Y(_00414_));
 sky130_fd_sc_hd__nor2_1 _22743_ (.A(_11954_),
    .B(_11629_),
    .Y(_02287_));
 sky130_fd_sc_hd__xnor2_1 _22744_ (.A(_11654_),
    .B(_02287_),
    .Y(_00415_));
 sky130_fd_sc_hd__nand2_1 _22745_ (.A(net176),
    .B(_11558_),
    .Y(_02288_));
 sky130_fd_sc_hd__xnor2_1 _22746_ (.A(net186),
    .B(_02288_),
    .Y(_00416_));
 sky130_fd_sc_hd__and2_1 _22747_ (.A(net186),
    .B(_11558_),
    .X(_02289_));
 sky130_fd_sc_hd__o21ai_1 _22748_ (.A1(_11413_),
    .A2(_02289_),
    .B1(net176),
    .Y(_02290_));
 sky130_fd_sc_hd__a22o_1 _22749_ (.A1(_11997_),
    .A2(_02289_),
    .B1(_02290_),
    .B2(net180),
    .X(_00417_));
 sky130_fd_sc_hd__nand2_1 _22750_ (.A(_11785_),
    .B(_12034_),
    .Y(_00418_));
 sky130_fd_sc_hd__o21a_2 _22751_ (.A1(net549),
    .A2(_07704_),
    .B1(_05443_),
    .X(_02291_));
 sky130_fd_sc_hd__clkbuf_4 _22752_ (.A(_02291_),
    .X(_02292_));
 sky130_fd_sc_hd__and4b_1 _22753_ (.A_N(net549),
    .B(_05442_),
    .C(net13),
    .D(net545),
    .X(_02293_));
 sky130_fd_sc_hd__buf_2 _22754_ (.A(_02293_),
    .X(_02294_));
 sky130_fd_sc_hd__clkbuf_4 _22755_ (.A(_02294_),
    .X(_02295_));
 sky130_fd_sc_hd__a22o_1 _22756_ (.A1(net991),
    .A2(_02292_),
    .B1(_02295_),
    .B2(\top0.pid_q.curr_int[0] ),
    .X(_00419_));
 sky130_fd_sc_hd__a22o_1 _22757_ (.A1(\top0.pid_q.prev_int[1] ),
    .A2(_02292_),
    .B1(_02295_),
    .B2(\top0.pid_q.curr_int[1] ),
    .X(_00420_));
 sky130_fd_sc_hd__a22o_1 _22758_ (.A1(net995),
    .A2(_02292_),
    .B1(_02295_),
    .B2(\top0.pid_q.curr_int[2] ),
    .X(_00421_));
 sky130_fd_sc_hd__a22o_1 _22759_ (.A1(net977),
    .A2(_02292_),
    .B1(_02295_),
    .B2(\top0.pid_q.curr_int[3] ),
    .X(_00422_));
 sky130_fd_sc_hd__a22o_1 _22760_ (.A1(net982),
    .A2(_02292_),
    .B1(_02295_),
    .B2(\top0.pid_q.curr_int[4] ),
    .X(_00423_));
 sky130_fd_sc_hd__a22o_1 _22761_ (.A1(\top0.pid_q.prev_int[5] ),
    .A2(_02292_),
    .B1(_02295_),
    .B2(\top0.pid_q.curr_int[5] ),
    .X(_00424_));
 sky130_fd_sc_hd__a22o_1 _22762_ (.A1(\top0.pid_q.prev_int[6] ),
    .A2(_02292_),
    .B1(_02295_),
    .B2(\top0.pid_q.curr_int[6] ),
    .X(_00425_));
 sky130_fd_sc_hd__a22o_1 _22763_ (.A1(net976),
    .A2(_02292_),
    .B1(_02295_),
    .B2(\top0.pid_q.curr_int[7] ),
    .X(_00426_));
 sky130_fd_sc_hd__a22o_1 _22764_ (.A1(\top0.pid_q.prev_int[8] ),
    .A2(_02292_),
    .B1(_02295_),
    .B2(net924),
    .X(_00427_));
 sky130_fd_sc_hd__a22o_1 _22765_ (.A1(net970),
    .A2(_02292_),
    .B1(_02295_),
    .B2(\top0.pid_q.curr_int[9] ),
    .X(_00428_));
 sky130_fd_sc_hd__a22o_1 _22766_ (.A1(net988),
    .A2(_02291_),
    .B1(_02294_),
    .B2(\top0.pid_q.curr_int[10] ),
    .X(_00429_));
 sky130_fd_sc_hd__a22o_1 _22767_ (.A1(net914),
    .A2(_02291_),
    .B1(_02294_),
    .B2(\top0.pid_q.curr_int[11] ),
    .X(_00430_));
 sky130_fd_sc_hd__a22o_1 _22768_ (.A1(\top0.pid_q.prev_int[12] ),
    .A2(_02291_),
    .B1(_02294_),
    .B2(\top0.pid_q.curr_int[12] ),
    .X(_00431_));
 sky130_fd_sc_hd__a22o_1 _22769_ (.A1(\top0.pid_q.prev_int[13] ),
    .A2(_02291_),
    .B1(_02294_),
    .B2(\top0.pid_q.curr_int[13] ),
    .X(_00432_));
 sky130_fd_sc_hd__a22o_1 _22770_ (.A1(\top0.pid_q.prev_int[14] ),
    .A2(_02291_),
    .B1(_02294_),
    .B2(\top0.pid_q.curr_int[14] ),
    .X(_00433_));
 sky130_fd_sc_hd__a22o_1 _22771_ (.A1(\top0.pid_q.prev_int[15] ),
    .A2(_02291_),
    .B1(_02294_),
    .B2(net772),
    .X(_00434_));
 sky130_fd_sc_hd__nor2_1 _22772_ (.A(_07115_),
    .B(_06276_),
    .Y(_02296_));
 sky130_fd_sc_hd__clkbuf_4 _22773_ (.A(_02296_),
    .X(_02297_));
 sky130_fd_sc_hd__inv_2 _22774_ (.A(\top0.svm0.counter[0] ),
    .Y(_02298_));
 sky130_fd_sc_hd__or4_1 _22775_ (.A(_02298_),
    .B(\top0.svm0.counter[1] ),
    .C(\top0.svm0.counter[2] ),
    .D(\top0.svm0.counter[3] ),
    .X(_02299_));
 sky130_fd_sc_hd__or4_1 _22776_ (.A(\top0.svm0.counter[5] ),
    .B(\top0.svm0.counter[6] ),
    .C(\top0.svm0.counter[8] ),
    .D(\top0.svm0.rising ),
    .X(_02300_));
 sky130_fd_sc_hd__or4_1 _22777_ (.A(\top0.svm0.counter[9] ),
    .B(net169),
    .C(\top0.svm0.counter[11] ),
    .D(\top0.svm0.counter[12] ),
    .X(_02301_));
 sky130_fd_sc_hd__or2_1 _22778_ (.A(_02300_),
    .B(_02301_),
    .X(_02302_));
 sky130_fd_sc_hd__or4_1 _22779_ (.A(\top0.svm0.counter[4] ),
    .B(net170),
    .C(_02299_),
    .D(_02302_),
    .X(_02303_));
 sky130_fd_sc_hd__or4_1 _22780_ (.A(\top0.svm0.counter[13] ),
    .B(\top0.svm0.counter[14] ),
    .C(\top0.svm0.counter[15] ),
    .D(_02303_),
    .X(_02304_));
 sky130_fd_sc_hd__nand2_1 _22781_ (.A(_02296_),
    .B(_02304_),
    .Y(_02305_));
 sky130_fd_sc_hd__clkbuf_4 _22782_ (.A(_07113_),
    .X(_02306_));
 sky130_fd_sc_hd__o21ai_1 _22783_ (.A1(net171),
    .A2(_02306_),
    .B1(_02305_),
    .Y(_02307_));
 sky130_fd_sc_hd__a22o_1 _22784_ (.A1(_02297_),
    .A2(_02305_),
    .B1(_02307_),
    .B2(\top0.svm0.out_valid ),
    .X(_00435_));
 sky130_fd_sc_hd__inv_4 _22785_ (.A(\top0.svm0.state[0] ),
    .Y(_02308_));
 sky130_fd_sc_hd__clkbuf_4 _22786_ (.A(_07115_),
    .X(_02309_));
 sky130_fd_sc_hd__o211a_1 _22787_ (.A1(\top0.svm0.state[1] ),
    .A2(\top0.start_svm ),
    .B1(_02308_),
    .C1(_02309_),
    .X(_00436_));
 sky130_fd_sc_hd__or2_1 _22788_ (.A(_05719_),
    .B(_05717_),
    .X(_02310_));
 sky130_fd_sc_hd__clkbuf_1 _22789_ (.A(_02310_),
    .X(_00437_));
 sky130_fd_sc_hd__a21o_1 _22790_ (.A1(_02297_),
    .A2(_02304_),
    .B1(_06381_),
    .X(_00438_));
 sky130_fd_sc_hd__xor2_1 _22791_ (.A(\top0.svm0.counter[12] ),
    .B(\top0.svm0.tA[12] ),
    .X(_02311_));
 sky130_fd_sc_hd__xor2_1 _22792_ (.A(net168),
    .B(\top0.svm0.tA[14] ),
    .X(_02312_));
 sky130_fd_sc_hd__inv_2 _22793_ (.A(\top0.svm0.counter[15] ),
    .Y(_02313_));
 sky130_fd_sc_hd__nor2_1 _22794_ (.A(_02313_),
    .B(\top0.svm0.tA[15] ),
    .Y(_02314_));
 sky130_fd_sc_hd__nand2_1 _22795_ (.A(_02313_),
    .B(\top0.svm0.tA[15] ),
    .Y(_02315_));
 sky130_fd_sc_hd__inv_2 _22796_ (.A(_02315_),
    .Y(_02316_));
 sky130_fd_sc_hd__inv_2 _22797_ (.A(\top0.svm0.counter[13] ),
    .Y(_02317_));
 sky130_fd_sc_hd__and2_1 _22798_ (.A(_02317_),
    .B(\top0.svm0.tA[13] ),
    .X(_02318_));
 sky130_fd_sc_hd__or2_1 _22799_ (.A(_02317_),
    .B(\top0.svm0.tA[13] ),
    .X(_02319_));
 sky130_fd_sc_hd__or4b_1 _22800_ (.A(_02314_),
    .B(_02316_),
    .C(_02318_),
    .D_N(_02319_),
    .X(_02320_));
 sky130_fd_sc_hd__or3_1 _22801_ (.A(_02311_),
    .B(_02312_),
    .C(_02320_),
    .X(_02321_));
 sky130_fd_sc_hd__inv_2 _22802_ (.A(\top0.svm0.tA[4] ),
    .Y(_02322_));
 sky130_fd_sc_hd__inv_2 _22803_ (.A(\top0.svm0.tA[5] ),
    .Y(_02323_));
 sky130_fd_sc_hd__inv_2 _22804_ (.A(\top0.svm0.counter[6] ),
    .Y(_02324_));
 sky130_fd_sc_hd__nor2_1 _22805_ (.A(_02324_),
    .B(\top0.svm0.tA[6] ),
    .Y(_02325_));
 sky130_fd_sc_hd__and2_1 _22806_ (.A(_02324_),
    .B(\top0.svm0.tA[6] ),
    .X(_02326_));
 sky130_fd_sc_hd__or2_1 _22807_ (.A(_02325_),
    .B(_02326_),
    .X(_02327_));
 sky130_fd_sc_hd__and2b_1 _22808_ (.A_N(net170),
    .B(\top0.svm0.tA[7] ),
    .X(_02328_));
 sky130_fd_sc_hd__and2b_1 _22809_ (.A_N(\top0.svm0.tA[7] ),
    .B(net170),
    .X(_02329_));
 sky130_fd_sc_hd__a2111o_1 _22810_ (.A1(\top0.svm0.counter[5] ),
    .A2(_02323_),
    .B1(_02327_),
    .C1(_02328_),
    .D1(_02329_),
    .X(_02330_));
 sky130_fd_sc_hd__inv_2 _22811_ (.A(\top0.svm0.counter[5] ),
    .Y(_02331_));
 sky130_fd_sc_hd__inv_2 _22812_ (.A(\top0.svm0.counter[4] ),
    .Y(_02332_));
 sky130_fd_sc_hd__a22o_1 _22813_ (.A1(_02331_),
    .A2(\top0.svm0.tA[5] ),
    .B1(\top0.svm0.tA[4] ),
    .B2(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__nand2_1 _22814_ (.A(\top0.svm0.counter[8] ),
    .B(\top0.svm0.tA[8] ),
    .Y(_02334_));
 sky130_fd_sc_hd__or2_1 _22815_ (.A(\top0.svm0.counter[8] ),
    .B(\top0.svm0.tA[8] ),
    .X(_02335_));
 sky130_fd_sc_hd__or2_1 _22816_ (.A(\top0.svm0.counter[9] ),
    .B(\top0.svm0.tA[9] ),
    .X(_02336_));
 sky130_fd_sc_hd__nand2_1 _22817_ (.A(\top0.svm0.counter[9] ),
    .B(\top0.svm0.tA[9] ),
    .Y(_02337_));
 sky130_fd_sc_hd__a22o_1 _22818_ (.A1(_02334_),
    .A2(_02335_),
    .B1(_02336_),
    .B2(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__inv_2 _22819_ (.A(\top0.svm0.counter[3] ),
    .Y(_02339_));
 sky130_fd_sc_hd__nor2_1 _22820_ (.A(_02339_),
    .B(\top0.svm0.tA[3] ),
    .Y(_02340_));
 sky130_fd_sc_hd__and2_1 _22821_ (.A(_02339_),
    .B(\top0.svm0.tA[3] ),
    .X(_02341_));
 sky130_fd_sc_hd__and2b_1 _22822_ (.A_N(\top0.svm0.counter[10] ),
    .B(\top0.svm0.tA[10] ),
    .X(_02342_));
 sky130_fd_sc_hd__or2b_1 _22823_ (.A(\top0.svm0.tA[10] ),
    .B_N(net169),
    .X(_02343_));
 sky130_fd_sc_hd__or4b_1 _22824_ (.A(_02340_),
    .B(_02341_),
    .C(_02342_),
    .D_N(_02343_),
    .X(_02344_));
 sky130_fd_sc_hd__inv_2 _22825_ (.A(\top0.svm0.counter[11] ),
    .Y(_02345_));
 sky130_fd_sc_hd__nor2_1 _22826_ (.A(_02345_),
    .B(\top0.svm0.tA[11] ),
    .Y(_02346_));
 sky130_fd_sc_hd__inv_2 _22827_ (.A(\top0.svm0.counter[2] ),
    .Y(_02347_));
 sky130_fd_sc_hd__and2_1 _22828_ (.A(_02347_),
    .B(\top0.svm0.tA[2] ),
    .X(_02348_));
 sky130_fd_sc_hd__nor2_1 _22829_ (.A(_02347_),
    .B(\top0.svm0.tA[2] ),
    .Y(_02349_));
 sky130_fd_sc_hd__and2_1 _22830_ (.A(_02345_),
    .B(\top0.svm0.tA[11] ),
    .X(_02350_));
 sky130_fd_sc_hd__or4_1 _22831_ (.A(_02346_),
    .B(_02348_),
    .C(_02349_),
    .D(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__inv_2 _22832_ (.A(\top0.svm0.counter[1] ),
    .Y(_02352_));
 sky130_fd_sc_hd__nor2_1 _22833_ (.A(_02352_),
    .B(\top0.svm0.tA[1] ),
    .Y(_02353_));
 sky130_fd_sc_hd__a21o_1 _22834_ (.A1(_02298_),
    .A2(\top0.svm0.tA[0] ),
    .B1(_02353_),
    .X(_02354_));
 sky130_fd_sc_hd__nor2_1 _22835_ (.A(_02298_),
    .B(\top0.svm0.tA[0] ),
    .Y(_02355_));
 sky130_fd_sc_hd__nand2_1 _22836_ (.A(_02352_),
    .B(\top0.svm0.tA[1] ),
    .Y(_02356_));
 sky130_fd_sc_hd__or3b_1 _22837_ (.A(_02354_),
    .B(_02355_),
    .C_N(_02356_),
    .X(_02357_));
 sky130_fd_sc_hd__or4_1 _22838_ (.A(_02338_),
    .B(_02344_),
    .C(_02351_),
    .D(_02357_),
    .X(_02358_));
 sky130_fd_sc_hd__a2111o_1 _22839_ (.A1(\top0.svm0.counter[4] ),
    .A2(_02322_),
    .B1(_02330_),
    .C1(_02333_),
    .D1(_02358_),
    .X(_02359_));
 sky130_fd_sc_hd__inv_2 _22840_ (.A(\top0.svm0.counter[9] ),
    .Y(_02360_));
 sky130_fd_sc_hd__a2111oi_1 _22841_ (.A1(\top0.svm0.counter[5] ),
    .A2(_02323_),
    .B1(_02327_),
    .C1(_02328_),
    .D1(_02329_),
    .Y(_02361_));
 sky130_fd_sc_hd__a2111oi_1 _22842_ (.A1(\top0.svm0.counter[4] ),
    .A2(_02322_),
    .B1(_02330_),
    .C1(_02340_),
    .D1(_02333_),
    .Y(_02362_));
 sky130_fd_sc_hd__a211o_1 _22843_ (.A1(_02356_),
    .A2(_02355_),
    .B1(_02353_),
    .C1(_02349_),
    .X(_02363_));
 sky130_fd_sc_hd__or3b_1 _22844_ (.A(_02341_),
    .B(_02348_),
    .C_N(_02363_),
    .X(_02364_));
 sky130_fd_sc_hd__o21ba_1 _22845_ (.A1(_02326_),
    .A2(_02328_),
    .B1_N(_02329_),
    .X(_02365_));
 sky130_fd_sc_hd__a221o_1 _22846_ (.A1(_02361_),
    .A2(_02333_),
    .B1(_02362_),
    .B2(_02364_),
    .C1(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__inv_2 _22847_ (.A(\top0.svm0.counter[8] ),
    .Y(_02367_));
 sky130_fd_sc_hd__o21a_1 _22848_ (.A1(\top0.svm0.tA[8] ),
    .A2(_02366_),
    .B1(_02367_),
    .X(_02368_));
 sky130_fd_sc_hd__and2_1 _22849_ (.A(\top0.svm0.tA[8] ),
    .B(_02366_),
    .X(_02369_));
 sky130_fd_sc_hd__o22a_1 _22850_ (.A1(_02360_),
    .A2(\top0.svm0.tA[9] ),
    .B1(_02368_),
    .B2(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__a21o_1 _22851_ (.A1(_02360_),
    .A2(\top0.svm0.tA[9] ),
    .B1(_02370_),
    .X(_02371_));
 sky130_fd_sc_hd__a21oi_1 _22852_ (.A1(_02371_),
    .A2(_02343_),
    .B1(_02342_),
    .Y(_02372_));
 sky130_fd_sc_hd__o21ba_1 _22853_ (.A1(_02346_),
    .A2(_02372_),
    .B1_N(_02350_),
    .X(_02373_));
 sky130_fd_sc_hd__inv_2 _22854_ (.A(\top0.svm0.counter[12] ),
    .Y(_02374_));
 sky130_fd_sc_hd__a31o_1 _22855_ (.A1(_02374_),
    .A2(\top0.svm0.tA[12] ),
    .A3(_02319_),
    .B1(_02318_),
    .X(_02375_));
 sky130_fd_sc_hd__nand2_1 _22856_ (.A(\top0.svm0.tA[14] ),
    .B(_02375_),
    .Y(_02376_));
 sky130_fd_sc_hd__nor2_1 _22857_ (.A(\top0.svm0.tA[14] ),
    .B(_02375_),
    .Y(_02377_));
 sky130_fd_sc_hd__a211o_1 _22858_ (.A1(net168),
    .A2(_02376_),
    .B1(_02377_),
    .C1(_02314_),
    .X(_02378_));
 sky130_fd_sc_hd__o211a_1 _22859_ (.A1(_02321_),
    .A2(_02373_),
    .B1(_02378_),
    .C1(_02315_),
    .X(_02379_));
 sky130_fd_sc_hd__o21bai_1 _22860_ (.A1(_02321_),
    .A2(_02359_),
    .B1_N(_02379_),
    .Y(_02380_));
 sky130_fd_sc_hd__a32o_1 _22861_ (.A1(\top0.svm0.calc_ready ),
    .A2(_02297_),
    .A3(_02380_),
    .B1(net704),
    .B2(_02309_),
    .X(_00439_));
 sky130_fd_sc_hd__inv_2 _22862_ (.A(\top0.svm0.tB[10] ),
    .Y(_02381_));
 sky130_fd_sc_hd__o211a_1 _22863_ (.A1(_02352_),
    .A2(\top0.svm0.tB[1] ),
    .B1(\top0.svm0.tB[0] ),
    .C1(_02298_),
    .X(_02382_));
 sky130_fd_sc_hd__a221o_1 _22864_ (.A1(_02352_),
    .A2(\top0.svm0.tB[1] ),
    .B1(\top0.svm0.tB[2] ),
    .B2(_02347_),
    .C1(_02382_),
    .X(_02383_));
 sky130_fd_sc_hd__o21a_1 _22865_ (.A1(_02347_),
    .A2(\top0.svm0.tB[2] ),
    .B1(_02383_),
    .X(_02384_));
 sky130_fd_sc_hd__a21o_1 _22866_ (.A1(\top0.svm0.tB[3] ),
    .A2(_02384_),
    .B1(_02339_),
    .X(_02385_));
 sky130_fd_sc_hd__o221a_1 _22867_ (.A1(_02332_),
    .A2(\top0.svm0.tB[4] ),
    .B1(_02384_),
    .B2(\top0.svm0.tB[3] ),
    .C1(_02385_),
    .X(_02386_));
 sky130_fd_sc_hd__a21o_1 _22868_ (.A1(_02332_),
    .A2(\top0.svm0.tB[4] ),
    .B1(_02386_),
    .X(_02387_));
 sky130_fd_sc_hd__o21a_1 _22869_ (.A1(\top0.svm0.tB[5] ),
    .A2(_02387_),
    .B1(_02331_),
    .X(_02388_));
 sky130_fd_sc_hd__a221o_1 _22870_ (.A1(_02324_),
    .A2(\top0.svm0.tB[6] ),
    .B1(\top0.svm0.tB[5] ),
    .B2(_02387_),
    .C1(_02388_),
    .X(_02389_));
 sky130_fd_sc_hd__o21a_1 _22871_ (.A1(_02324_),
    .A2(\top0.svm0.tB[6] ),
    .B1(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__o21ba_1 _22872_ (.A1(\top0.svm0.tB[7] ),
    .A2(_02390_),
    .B1_N(net170),
    .X(_02391_));
 sky130_fd_sc_hd__and2_1 _22873_ (.A(\top0.svm0.tB[7] ),
    .B(_02390_),
    .X(_02392_));
 sky130_fd_sc_hd__o22a_1 _22874_ (.A1(_02367_),
    .A2(\top0.svm0.tB[8] ),
    .B1(_02391_),
    .B2(_02392_),
    .X(_02393_));
 sky130_fd_sc_hd__a21o_1 _22875_ (.A1(_02367_),
    .A2(\top0.svm0.tB[8] ),
    .B1(_02393_),
    .X(_02394_));
 sky130_fd_sc_hd__o21a_1 _22876_ (.A1(\top0.svm0.tB[9] ),
    .A2(_02394_),
    .B1(_02360_),
    .X(_02395_));
 sky130_fd_sc_hd__a21oi_1 _22877_ (.A1(\top0.svm0.tB[9] ),
    .A2(_02394_),
    .B1(_02395_),
    .Y(_02396_));
 sky130_fd_sc_hd__a21o_1 _22878_ (.A1(net169),
    .A2(_02381_),
    .B1(_02396_),
    .X(_02397_));
 sky130_fd_sc_hd__o21ai_1 _22879_ (.A1(net169),
    .A2(_02381_),
    .B1(_02397_),
    .Y(_02398_));
 sky130_fd_sc_hd__o21a_1 _22880_ (.A1(\top0.svm0.tB[11] ),
    .A2(_02398_),
    .B1(_02345_),
    .X(_02399_));
 sky130_fd_sc_hd__and2_1 _22881_ (.A(\top0.svm0.tB[11] ),
    .B(_02398_),
    .X(_02400_));
 sky130_fd_sc_hd__o22a_1 _22882_ (.A1(_02374_),
    .A2(\top0.svm0.tB[12] ),
    .B1(_02399_),
    .B2(_02400_),
    .X(_02401_));
 sky130_fd_sc_hd__and2_1 _22883_ (.A(_02374_),
    .B(\top0.svm0.tB[12] ),
    .X(_02402_));
 sky130_fd_sc_hd__o22a_1 _22884_ (.A1(_02317_),
    .A2(\top0.svm0.tB[13] ),
    .B1(_02401_),
    .B2(_02402_),
    .X(_02403_));
 sky130_fd_sc_hd__a21o_1 _22885_ (.A1(_02317_),
    .A2(\top0.svm0.tB[13] ),
    .B1(_02403_),
    .X(_02404_));
 sky130_fd_sc_hd__inv_2 _22886_ (.A(net168),
    .Y(_02405_));
 sky130_fd_sc_hd__o21a_1 _22887_ (.A1(\top0.svm0.tB[14] ),
    .A2(_02404_),
    .B1(_02405_),
    .X(_02406_));
 sky130_fd_sc_hd__a221o_1 _22888_ (.A1(_02313_),
    .A2(\top0.svm0.tB[15] ),
    .B1(\top0.svm0.tB[14] ),
    .B2(_02404_),
    .C1(_02406_),
    .X(_02407_));
 sky130_fd_sc_hd__o21ai_1 _22889_ (.A1(_02313_),
    .A2(\top0.svm0.tB[15] ),
    .B1(_02407_),
    .Y(_02408_));
 sky130_fd_sc_hd__a32o_1 _22890_ (.A1(\top0.svm0.calc_ready ),
    .A2(_02297_),
    .A3(_02408_),
    .B1(net708),
    .B2(_02309_),
    .X(_00440_));
 sky130_fd_sc_hd__inv_2 _22891_ (.A(\top0.svm0.tC[10] ),
    .Y(_02409_));
 sky130_fd_sc_hd__o211a_1 _22892_ (.A1(_02352_),
    .A2(\top0.svm0.tC[1] ),
    .B1(\top0.svm0.tC[0] ),
    .C1(_02298_),
    .X(_02410_));
 sky130_fd_sc_hd__a221o_1 _22893_ (.A1(_02352_),
    .A2(\top0.svm0.tC[1] ),
    .B1(\top0.svm0.tC[2] ),
    .B2(_02347_),
    .C1(_02410_),
    .X(_02411_));
 sky130_fd_sc_hd__o21a_1 _22894_ (.A1(_02347_),
    .A2(\top0.svm0.tC[2] ),
    .B1(_02411_),
    .X(_02412_));
 sky130_fd_sc_hd__a21o_1 _22895_ (.A1(\top0.svm0.tC[3] ),
    .A2(_02412_),
    .B1(_02339_),
    .X(_02413_));
 sky130_fd_sc_hd__o221a_1 _22896_ (.A1(_02332_),
    .A2(\top0.svm0.tC[4] ),
    .B1(_02412_),
    .B2(\top0.svm0.tC[3] ),
    .C1(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__a21o_1 _22897_ (.A1(_02332_),
    .A2(\top0.svm0.tC[4] ),
    .B1(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__o21a_1 _22898_ (.A1(\top0.svm0.tC[5] ),
    .A2(_02415_),
    .B1(_02331_),
    .X(_02416_));
 sky130_fd_sc_hd__a221o_1 _22899_ (.A1(_02324_),
    .A2(\top0.svm0.tC[6] ),
    .B1(\top0.svm0.tC[5] ),
    .B2(_02415_),
    .C1(_02416_),
    .X(_02417_));
 sky130_fd_sc_hd__o21a_1 _22900_ (.A1(_02324_),
    .A2(\top0.svm0.tC[6] ),
    .B1(_02417_),
    .X(_02418_));
 sky130_fd_sc_hd__o21ba_1 _22901_ (.A1(\top0.svm0.tC[7] ),
    .A2(_02418_),
    .B1_N(\top0.svm0.counter[7] ),
    .X(_02419_));
 sky130_fd_sc_hd__and2_1 _22902_ (.A(\top0.svm0.tC[7] ),
    .B(_02418_),
    .X(_02420_));
 sky130_fd_sc_hd__o22a_1 _22903_ (.A1(_02367_),
    .A2(\top0.svm0.tC[8] ),
    .B1(_02419_),
    .B2(_02420_),
    .X(_02421_));
 sky130_fd_sc_hd__a21o_1 _22904_ (.A1(_02367_),
    .A2(\top0.svm0.tC[8] ),
    .B1(_02421_),
    .X(_02422_));
 sky130_fd_sc_hd__o21a_1 _22905_ (.A1(\top0.svm0.tC[9] ),
    .A2(_02422_),
    .B1(_02360_),
    .X(_02423_));
 sky130_fd_sc_hd__a21oi_1 _22906_ (.A1(\top0.svm0.tC[9] ),
    .A2(_02422_),
    .B1(_02423_),
    .Y(_02424_));
 sky130_fd_sc_hd__a21oi_1 _22907_ (.A1(net169),
    .A2(_02409_),
    .B1(_02424_),
    .Y(_02425_));
 sky130_fd_sc_hd__nor2_1 _22908_ (.A(net169),
    .B(_02409_),
    .Y(_02426_));
 sky130_fd_sc_hd__o22a_1 _22909_ (.A1(_02345_),
    .A2(\top0.svm0.tC[11] ),
    .B1(_02425_),
    .B2(_02426_),
    .X(_02427_));
 sky130_fd_sc_hd__a221o_1 _22910_ (.A1(_02374_),
    .A2(\top0.svm0.tC[12] ),
    .B1(\top0.svm0.tC[11] ),
    .B2(_02345_),
    .C1(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__o221a_1 _22911_ (.A1(_02317_),
    .A2(\top0.svm0.tC[13] ),
    .B1(\top0.svm0.tC[12] ),
    .B2(_02374_),
    .C1(_02428_),
    .X(_02429_));
 sky130_fd_sc_hd__a221o_1 _22912_ (.A1(_02405_),
    .A2(\top0.svm0.tC[14] ),
    .B1(\top0.svm0.tC[13] ),
    .B2(_02317_),
    .C1(_02429_),
    .X(_02430_));
 sky130_fd_sc_hd__or2_1 _22913_ (.A(_02405_),
    .B(\top0.svm0.tC[14] ),
    .X(_02431_));
 sky130_fd_sc_hd__a22o_1 _22914_ (.A1(_02313_),
    .A2(\top0.svm0.tC[15] ),
    .B1(_02430_),
    .B2(_02431_),
    .X(_02432_));
 sky130_fd_sc_hd__o21ai_1 _22915_ (.A1(_02313_),
    .A2(\top0.svm0.tC[15] ),
    .B1(_02432_),
    .Y(_02433_));
 sky130_fd_sc_hd__a32o_1 _22916_ (.A1(\top0.svm0.calc_ready ),
    .A2(_02297_),
    .A3(_02433_),
    .B1(net706),
    .B2(_02309_),
    .X(_00441_));
 sky130_fd_sc_hd__o21a_1 _22917_ (.A1(net555),
    .A2(_06277_),
    .B1(net172),
    .X(_02434_));
 sky130_fd_sc_hd__nor2_1 _22918_ (.A(_02298_),
    .B(_02434_),
    .Y(_02435_));
 sky130_fd_sc_hd__a31o_1 _22919_ (.A1(_02298_),
    .A2(net555),
    .A3(_02297_),
    .B1(_02435_),
    .X(_00442_));
 sky130_fd_sc_hd__nand2_1 _22920_ (.A(\top0.svm0.counter[0] ),
    .B(net555),
    .Y(_02436_));
 sky130_fd_sc_hd__xor2_1 _22921_ (.A(\top0.svm0.delta[1] ),
    .B(_02436_),
    .X(_02437_));
 sky130_fd_sc_hd__a21o_1 _22922_ (.A1(_02306_),
    .A2(_02437_),
    .B1(_02309_),
    .X(_02438_));
 sky130_fd_sc_hd__nand2_1 _22923_ (.A(net171),
    .B(_02306_),
    .Y(_02439_));
 sky130_fd_sc_hd__buf_2 _22924_ (.A(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__nor2_1 _22925_ (.A(_02440_),
    .B(_02437_),
    .Y(_02441_));
 sky130_fd_sc_hd__mux2_1 _22926_ (.A0(_02438_),
    .A1(_02441_),
    .S(_02352_),
    .X(_02442_));
 sky130_fd_sc_hd__clkbuf_1 _22927_ (.A(_02442_),
    .X(_00443_));
 sky130_fd_sc_hd__inv_2 _22928_ (.A(\top0.svm0.delta[2] ),
    .Y(_02443_));
 sky130_fd_sc_hd__nand2_1 _22929_ (.A(\top0.svm0.counter[1] ),
    .B(\top0.svm0.delta[1] ),
    .Y(_02444_));
 sky130_fd_sc_hd__o211ai_2 _22930_ (.A1(\top0.svm0.counter[1] ),
    .A2(\top0.svm0.delta[1] ),
    .B1(net555),
    .C1(\top0.svm0.counter[0] ),
    .Y(_02445_));
 sky130_fd_sc_hd__and3_1 _22931_ (.A(_02443_),
    .B(_02444_),
    .C(_02445_),
    .X(_02446_));
 sky130_fd_sc_hd__a21o_1 _22932_ (.A1(_02444_),
    .A2(_02445_),
    .B1(_02443_),
    .X(_02447_));
 sky130_fd_sc_hd__or2b_1 _22933_ (.A(_02446_),
    .B_N(_02447_),
    .X(_02448_));
 sky130_fd_sc_hd__a21o_1 _22934_ (.A1(_02306_),
    .A2(_02448_),
    .B1(_02309_),
    .X(_02449_));
 sky130_fd_sc_hd__nor2_1 _22935_ (.A(_02440_),
    .B(_02448_),
    .Y(_02450_));
 sky130_fd_sc_hd__mux2_1 _22936_ (.A0(_02449_),
    .A1(_02450_),
    .S(_02347_),
    .X(_02451_));
 sky130_fd_sc_hd__clkbuf_1 _22937_ (.A(_02451_),
    .X(_00444_));
 sky130_fd_sc_hd__a31o_1 _22938_ (.A1(_02443_),
    .A2(_02444_),
    .A3(_02445_),
    .B1(_02347_),
    .X(_02452_));
 sky130_fd_sc_hd__nand2_1 _22939_ (.A(_02447_),
    .B(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__xnor2_1 _22940_ (.A(\top0.svm0.delta[3] ),
    .B(_02453_),
    .Y(_02454_));
 sky130_fd_sc_hd__a21o_1 _22941_ (.A1(_02306_),
    .A2(_02454_),
    .B1(_02309_),
    .X(_02455_));
 sky130_fd_sc_hd__nor2_1 _22942_ (.A(_02440_),
    .B(_02454_),
    .Y(_02456_));
 sky130_fd_sc_hd__mux2_1 _22943_ (.A0(_02455_),
    .A1(_02456_),
    .S(_02339_),
    .X(_02457_));
 sky130_fd_sc_hd__clkbuf_1 _22944_ (.A(_02457_),
    .X(_00445_));
 sky130_fd_sc_hd__inv_2 _22945_ (.A(\top0.svm0.delta[4] ),
    .Y(_02458_));
 sky130_fd_sc_hd__inv_2 _22946_ (.A(\top0.svm0.delta[3] ),
    .Y(_02459_));
 sky130_fd_sc_hd__a31o_1 _22947_ (.A1(_02459_),
    .A2(_02447_),
    .A3(_02452_),
    .B1(_02339_),
    .X(_02460_));
 sky130_fd_sc_hd__a21boi_2 _22948_ (.A1(\top0.svm0.delta[3] ),
    .A2(_02453_),
    .B1_N(_02460_),
    .Y(_02461_));
 sky130_fd_sc_hd__xnor2_1 _22949_ (.A(_02458_),
    .B(_02461_),
    .Y(_02462_));
 sky130_fd_sc_hd__a21o_1 _22950_ (.A1(_02306_),
    .A2(_02462_),
    .B1(_02309_),
    .X(_02463_));
 sky130_fd_sc_hd__nor2_1 _22951_ (.A(_02440_),
    .B(_02462_),
    .Y(_02464_));
 sky130_fd_sc_hd__mux2_1 _22952_ (.A0(_02463_),
    .A1(_02464_),
    .S(_02332_),
    .X(_02465_));
 sky130_fd_sc_hd__clkbuf_1 _22953_ (.A(_02465_),
    .X(_00446_));
 sky130_fd_sc_hd__inv_2 _22954_ (.A(\top0.svm0.delta[5] ),
    .Y(_02466_));
 sky130_fd_sc_hd__o21a_1 _22955_ (.A1(_02458_),
    .A2(_02461_),
    .B1(_02332_),
    .X(_02467_));
 sky130_fd_sc_hd__a21o_1 _22956_ (.A1(_02458_),
    .A2(_02461_),
    .B1(_02467_),
    .X(_02468_));
 sky130_fd_sc_hd__xnor2_1 _22957_ (.A(_02466_),
    .B(_02468_),
    .Y(_02469_));
 sky130_fd_sc_hd__a21o_1 _22958_ (.A1(_02306_),
    .A2(_02469_),
    .B1(_02309_),
    .X(_02470_));
 sky130_fd_sc_hd__nor2_1 _22959_ (.A(_02440_),
    .B(_02469_),
    .Y(_02471_));
 sky130_fd_sc_hd__mux2_1 _22960_ (.A0(_02470_),
    .A1(_02471_),
    .S(_02331_),
    .X(_02472_));
 sky130_fd_sc_hd__clkbuf_1 _22961_ (.A(_02472_),
    .X(_00447_));
 sky130_fd_sc_hd__o21a_1 _22962_ (.A1(_02466_),
    .A2(_02468_),
    .B1(_02331_),
    .X(_02473_));
 sky130_fd_sc_hd__a21o_1 _22963_ (.A1(_02466_),
    .A2(_02468_),
    .B1(_02473_),
    .X(_02474_));
 sky130_fd_sc_hd__xnor2_1 _22964_ (.A(\top0.svm0.delta[6] ),
    .B(_02474_),
    .Y(_02475_));
 sky130_fd_sc_hd__o21a_1 _22965_ (.A1(_06277_),
    .A2(_02475_),
    .B1(net172),
    .X(_02476_));
 sky130_fd_sc_hd__nor2_1 _22966_ (.A(_02324_),
    .B(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__a31o_1 _22967_ (.A1(_02324_),
    .A2(_02297_),
    .A3(_02475_),
    .B1(_02477_),
    .X(_00448_));
 sky130_fd_sc_hd__inv_2 _22968_ (.A(\top0.svm0.delta[6] ),
    .Y(_02478_));
 sky130_fd_sc_hd__a21o_1 _22969_ (.A1(_02478_),
    .A2(_02474_),
    .B1(_02324_),
    .X(_02479_));
 sky130_fd_sc_hd__o21a_1 _22970_ (.A1(_02478_),
    .A2(_02474_),
    .B1(_02479_),
    .X(_02480_));
 sky130_fd_sc_hd__xnor2_1 _22971_ (.A(\top0.svm0.delta[7] ),
    .B(_02480_),
    .Y(_02481_));
 sky130_fd_sc_hd__o21ai_1 _22972_ (.A1(_06277_),
    .A2(_02481_),
    .B1(net172),
    .Y(_02482_));
 sky130_fd_sc_hd__clkbuf_4 _22973_ (.A(_02440_),
    .X(_02483_));
 sky130_fd_sc_hd__nor2_1 _22974_ (.A(net170),
    .B(_02483_),
    .Y(_02484_));
 sky130_fd_sc_hd__a22o_1 _22975_ (.A1(net170),
    .A2(_02482_),
    .B1(_02484_),
    .B2(_02481_),
    .X(_00449_));
 sky130_fd_sc_hd__inv_2 _22976_ (.A(\top0.svm0.delta[7] ),
    .Y(_02485_));
 sky130_fd_sc_hd__o21ba_1 _22977_ (.A1(_02485_),
    .A2(_02480_),
    .B1_N(net170),
    .X(_02486_));
 sky130_fd_sc_hd__a21o_1 _22978_ (.A1(_02485_),
    .A2(_02480_),
    .B1(_02486_),
    .X(_02487_));
 sky130_fd_sc_hd__xnor2_1 _22979_ (.A(\top0.svm0.delta[8] ),
    .B(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__o21ai_1 _22980_ (.A1(_06277_),
    .A2(_02488_),
    .B1(net172),
    .Y(_02489_));
 sky130_fd_sc_hd__nor2_1 _22981_ (.A(\top0.svm0.counter[8] ),
    .B(_02483_),
    .Y(_02490_));
 sky130_fd_sc_hd__a22o_1 _22982_ (.A1(\top0.svm0.counter[8] ),
    .A2(_02489_),
    .B1(_02490_),
    .B2(_02488_),
    .X(_00450_));
 sky130_fd_sc_hd__inv_2 _22983_ (.A(\top0.svm0.delta[8] ),
    .Y(_02491_));
 sky130_fd_sc_hd__o21a_1 _22984_ (.A1(_02491_),
    .A2(_02487_),
    .B1(_02367_),
    .X(_02492_));
 sky130_fd_sc_hd__a21o_1 _22985_ (.A1(_02491_),
    .A2(_02487_),
    .B1(_02492_),
    .X(_02493_));
 sky130_fd_sc_hd__xnor2_1 _22986_ (.A(\top0.svm0.delta[9] ),
    .B(_02493_),
    .Y(_02494_));
 sky130_fd_sc_hd__o21ai_1 _22987_ (.A1(_06277_),
    .A2(_02494_),
    .B1(net172),
    .Y(_02495_));
 sky130_fd_sc_hd__nor2_1 _22988_ (.A(\top0.svm0.counter[9] ),
    .B(_02483_),
    .Y(_02496_));
 sky130_fd_sc_hd__a22o_1 _22989_ (.A1(\top0.svm0.counter[9] ),
    .A2(_02495_),
    .B1(_02496_),
    .B2(_02494_),
    .X(_00451_));
 sky130_fd_sc_hd__inv_2 _22990_ (.A(\top0.svm0.delta[9] ),
    .Y(_02497_));
 sky130_fd_sc_hd__o21a_1 _22991_ (.A1(_02497_),
    .A2(_02493_),
    .B1(_02360_),
    .X(_02498_));
 sky130_fd_sc_hd__a21oi_2 _22992_ (.A1(_02497_),
    .A2(_02493_),
    .B1(_02498_),
    .Y(_02499_));
 sky130_fd_sc_hd__xor2_1 _22993_ (.A(\top0.svm0.delta[10] ),
    .B(_02499_),
    .X(_02500_));
 sky130_fd_sc_hd__o21ai_1 _22994_ (.A1(_06277_),
    .A2(_02500_),
    .B1(net172),
    .Y(_02501_));
 sky130_fd_sc_hd__nor2_1 _22995_ (.A(net169),
    .B(_02483_),
    .Y(_02502_));
 sky130_fd_sc_hd__a22o_1 _22996_ (.A1(net169),
    .A2(_02501_),
    .B1(_02502_),
    .B2(_02500_),
    .X(_00452_));
 sky130_fd_sc_hd__a21o_1 _22997_ (.A1(\top0.svm0.delta[10] ),
    .A2(_02499_),
    .B1(net169),
    .X(_02503_));
 sky130_fd_sc_hd__o21ai_2 _22998_ (.A1(\top0.svm0.delta[10] ),
    .A2(_02499_),
    .B1(_02503_),
    .Y(_02504_));
 sky130_fd_sc_hd__xnor2_1 _22999_ (.A(\top0.svm0.delta[11] ),
    .B(_02504_),
    .Y(_02505_));
 sky130_fd_sc_hd__o21a_1 _23000_ (.A1(_06277_),
    .A2(_02505_),
    .B1(net171),
    .X(_02506_));
 sky130_fd_sc_hd__nor2_1 _23001_ (.A(_02345_),
    .B(_02506_),
    .Y(_02507_));
 sky130_fd_sc_hd__a31o_1 _23002_ (.A1(_02345_),
    .A2(_02297_),
    .A3(_02505_),
    .B1(_02507_),
    .X(_00453_));
 sky130_fd_sc_hd__inv_2 _23003_ (.A(\top0.svm0.delta[11] ),
    .Y(_02508_));
 sky130_fd_sc_hd__a21o_1 _23004_ (.A1(_02508_),
    .A2(_02504_),
    .B1(_02345_),
    .X(_02509_));
 sky130_fd_sc_hd__o21a_1 _23005_ (.A1(_02508_),
    .A2(_02504_),
    .B1(_02509_),
    .X(_02510_));
 sky130_fd_sc_hd__xnor2_1 _23006_ (.A(\top0.svm0.delta[12] ),
    .B(_02510_),
    .Y(_02511_));
 sky130_fd_sc_hd__o21a_1 _23007_ (.A1(_06277_),
    .A2(_02511_),
    .B1(net171),
    .X(_02512_));
 sky130_fd_sc_hd__nor2_1 _23008_ (.A(_02374_),
    .B(_02512_),
    .Y(_02513_));
 sky130_fd_sc_hd__a31o_1 _23009_ (.A1(_02374_),
    .A2(_02297_),
    .A3(_02511_),
    .B1(_02513_),
    .X(_00454_));
 sky130_fd_sc_hd__inv_2 _23010_ (.A(\top0.svm0.delta[12] ),
    .Y(_02514_));
 sky130_fd_sc_hd__o21a_1 _23011_ (.A1(_02514_),
    .A2(_02510_),
    .B1(_02374_),
    .X(_02515_));
 sky130_fd_sc_hd__a21o_1 _23012_ (.A1(_02514_),
    .A2(_02510_),
    .B1(_02515_),
    .X(_02516_));
 sky130_fd_sc_hd__xor2_1 _23013_ (.A(\top0.svm0.delta[13] ),
    .B(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__or3_1 _23014_ (.A(\top0.svm0.counter[13] ),
    .B(_02439_),
    .C(_02517_),
    .X(_02518_));
 sky130_fd_sc_hd__o21ai_1 _23015_ (.A1(net172),
    .A2(_02317_),
    .B1(_02518_),
    .Y(_02519_));
 sky130_fd_sc_hd__a31o_1 _23016_ (.A1(\top0.svm0.counter[13] ),
    .A2(_02306_),
    .A3(_02517_),
    .B1(_02519_),
    .X(_00455_));
 sky130_fd_sc_hd__nor2_1 _23017_ (.A(\top0.svm0.counter[13] ),
    .B(\top0.svm0.delta[13] ),
    .Y(_02520_));
 sky130_fd_sc_hd__nand2_1 _23018_ (.A(\top0.svm0.counter[13] ),
    .B(\top0.svm0.delta[13] ),
    .Y(_02521_));
 sky130_fd_sc_hd__o21ai_2 _23019_ (.A1(_02516_),
    .A2(_02520_),
    .B1(_02521_),
    .Y(_02522_));
 sky130_fd_sc_hd__xor2_1 _23020_ (.A(\top0.svm0.delta[14] ),
    .B(_02522_),
    .X(_02523_));
 sky130_fd_sc_hd__o21ai_1 _23021_ (.A1(_06277_),
    .A2(_02523_),
    .B1(net172),
    .Y(_02524_));
 sky130_fd_sc_hd__nor2_1 _23022_ (.A(net168),
    .B(_02483_),
    .Y(_02525_));
 sky130_fd_sc_hd__a22o_1 _23023_ (.A1(net168),
    .A2(_02524_),
    .B1(_02525_),
    .B2(_02523_),
    .X(_00456_));
 sky130_fd_sc_hd__and2_1 _23024_ (.A(net168),
    .B(\top0.svm0.delta[14] ),
    .X(_02526_));
 sky130_fd_sc_hd__xnor2_1 _23025_ (.A(\top0.svm0.counter[15] ),
    .B(\top0.svm0.delta[15] ),
    .Y(_02527_));
 sky130_fd_sc_hd__or3_1 _23026_ (.A(_02439_),
    .B(_02526_),
    .C(_02527_),
    .X(_02528_));
 sky130_fd_sc_hd__o2111ai_1 _23027_ (.A1(net168),
    .A2(\top0.svm0.delta[14] ),
    .B1(_02297_),
    .C1(_02522_),
    .D1(_02527_),
    .Y(_02529_));
 sky130_fd_sc_hd__nor2_1 _23028_ (.A(net168),
    .B(\top0.svm0.delta[14] ),
    .Y(_02530_));
 sky130_fd_sc_hd__mux2_1 _23029_ (.A0(_02530_),
    .A1(_02526_),
    .S(\top0.svm0.delta[15] ),
    .X(_02531_));
 sky130_fd_sc_hd__mux2_1 _23030_ (.A0(_02526_),
    .A1(_02530_),
    .S(\top0.svm0.delta[15] ),
    .X(_02532_));
 sky130_fd_sc_hd__nor2_1 _23031_ (.A(_07115_),
    .B(\top0.svm0.counter[15] ),
    .Y(_02533_));
 sky130_fd_sc_hd__a22o_1 _23032_ (.A1(\top0.svm0.counter[15] ),
    .A2(_02531_),
    .B1(_02532_),
    .B2(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__a22oi_1 _23033_ (.A1(_02309_),
    .A2(\top0.svm0.counter[15] ),
    .B1(_02306_),
    .B2(_02534_),
    .Y(_02535_));
 sky130_fd_sc_hd__o211ai_1 _23034_ (.A1(_02522_),
    .A2(_02528_),
    .B1(_02529_),
    .C1(_02535_),
    .Y(_00457_));
 sky130_fd_sc_hd__nand2_1 _23035_ (.A(net21),
    .B(\top0.svm0.counter[15] ),
    .Y(_02536_));
 sky130_fd_sc_hd__or2_1 _23036_ (.A(net20),
    .B(\top0.svm0.counter[15] ),
    .X(_02537_));
 sky130_fd_sc_hd__or3_1 _23037_ (.A(net65),
    .B(net63),
    .C(net61),
    .X(_02538_));
 sky130_fd_sc_hd__or2_1 _23038_ (.A(net57),
    .B(_02538_),
    .X(_02539_));
 sky130_fd_sc_hd__or4_2 _23039_ (.A(net54),
    .B(net52),
    .C(net49),
    .D(_02539_),
    .X(_02540_));
 sky130_fd_sc_hd__or4_1 _23040_ (.A(net46),
    .B(net44),
    .C(\top0.periodTop_r[9] ),
    .D(_02540_),
    .X(_02541_));
 sky130_fd_sc_hd__or2_1 _23041_ (.A(net40),
    .B(_02541_),
    .X(_02542_));
 sky130_fd_sc_hd__or4_2 _23042_ (.A(net36),
    .B(net34),
    .C(net32),
    .D(_02542_),
    .X(_02543_));
 sky130_fd_sc_hd__nand2_1 _23043_ (.A(net168),
    .B(_02543_),
    .Y(_02544_));
 sky130_fd_sc_hd__or2_1 _23044_ (.A(net168),
    .B(_02543_),
    .X(_02545_));
 sky130_fd_sc_hd__a21o_1 _23045_ (.A1(_02544_),
    .A2(_02545_),
    .B1(_06217_),
    .X(_02546_));
 sky130_fd_sc_hd__or3b_1 _23046_ (.A(net26),
    .B(\top0.svm0.counter[14] ),
    .C_N(_02543_),
    .X(_02547_));
 sky130_fd_sc_hd__a22o_1 _23047_ (.A1(_02536_),
    .A2(_02537_),
    .B1(_02546_),
    .B2(_02547_),
    .X(_02548_));
 sky130_fd_sc_hd__or4b_1 _23048_ (.A(\top0.svm0.counter[15] ),
    .B(_06777_),
    .C(_02543_),
    .D_N(\top0.svm0.counter[14] ),
    .X(_02549_));
 sky130_fd_sc_hd__nor2_1 _23049_ (.A(net36),
    .B(_02542_),
    .Y(_02550_));
 sky130_fd_sc_hd__xnor2_1 _23050_ (.A(\top0.svm0.counter[12] ),
    .B(_02550_),
    .Y(_02551_));
 sky130_fd_sc_hd__or3_1 _23051_ (.A(net34),
    .B(\top0.svm0.counter[12] ),
    .C(_02550_),
    .X(_02552_));
 sky130_fd_sc_hd__o21a_1 _23052_ (.A1(_05500_),
    .A2(_02551_),
    .B1(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__xnor2_1 _23053_ (.A(net32),
    .B(\top0.svm0.counter[13] ),
    .Y(_02554_));
 sky130_fd_sc_hd__a31o_1 _23054_ (.A1(_05500_),
    .A2(\top0.svm0.counter[12] ),
    .A3(_02550_),
    .B1(_02554_),
    .X(_02555_));
 sky130_fd_sc_hd__a21bo_1 _23055_ (.A1(_02553_),
    .A2(_02554_),
    .B1_N(_02555_),
    .X(_02556_));
 sky130_fd_sc_hd__nor2_1 _23056_ (.A(\top0.periodTop_r[4] ),
    .B(_02539_),
    .Y(_02557_));
 sky130_fd_sc_hd__xnor2_1 _23057_ (.A(\top0.svm0.counter[5] ),
    .B(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__or3_1 _23058_ (.A(net52),
    .B(\top0.svm0.counter[5] ),
    .C(_02557_),
    .X(_02559_));
 sky130_fd_sc_hd__o21a_1 _23059_ (.A1(_05541_),
    .A2(_02558_),
    .B1(_02559_),
    .X(_02560_));
 sky130_fd_sc_hd__xnor2_1 _23060_ (.A(net49),
    .B(\top0.svm0.counter[6] ),
    .Y(_02561_));
 sky130_fd_sc_hd__a31o_1 _23061_ (.A1(_05541_),
    .A2(\top0.svm0.counter[5] ),
    .A3(_02557_),
    .B1(_02561_),
    .X(_02562_));
 sky130_fd_sc_hd__a21bo_1 _23062_ (.A1(_02560_),
    .A2(_02561_),
    .B1_N(_02562_),
    .X(_02563_));
 sky130_fd_sc_hd__xor2_1 _23063_ (.A(net42),
    .B(\top0.svm0.counter[9] ),
    .X(_02564_));
 sky130_fd_sc_hd__xor2_1 _23064_ (.A(net170),
    .B(_02540_),
    .X(_02565_));
 sky130_fd_sc_hd__nand2_1 _23065_ (.A(_05565_),
    .B(\top0.svm0.counter[8] ),
    .Y(_02566_));
 sky130_fd_sc_hd__nor2_1 _23066_ (.A(net46),
    .B(_02540_),
    .Y(_02567_));
 sky130_fd_sc_hd__nand2_1 _23067_ (.A(net44),
    .B(_02367_),
    .Y(_02568_));
 sky130_fd_sc_hd__o221a_1 _23068_ (.A1(_05573_),
    .A2(_02565_),
    .B1(_02566_),
    .B2(_02567_),
    .C1(_02568_),
    .X(_02569_));
 sky130_fd_sc_hd__or3b_1 _23069_ (.A(net170),
    .B(_02564_),
    .C_N(_02540_),
    .X(_02570_));
 sky130_fd_sc_hd__or3b_1 _23070_ (.A(_02540_),
    .B(_02566_),
    .C_N(_02564_),
    .X(_02571_));
 sky130_fd_sc_hd__a21o_1 _23071_ (.A1(_02570_),
    .A2(_02571_),
    .B1(net46),
    .X(_02572_));
 sky130_fd_sc_hd__o21a_1 _23072_ (.A1(_02564_),
    .A2(_02569_),
    .B1(_02572_),
    .X(_02573_));
 sky130_fd_sc_hd__xor2_1 _23073_ (.A(net61),
    .B(\top0.svm0.counter[2] ),
    .X(_02574_));
 sky130_fd_sc_hd__xor2_1 _23074_ (.A(net63),
    .B(\top0.svm0.counter[1] ),
    .X(_02575_));
 sky130_fd_sc_hd__or4_1 _23075_ (.A(\top0.svm0.counter[0] ),
    .B(_05805_),
    .C(_02574_),
    .D(_02575_),
    .X(_02576_));
 sky130_fd_sc_hd__or3_1 _23076_ (.A(_05607_),
    .B(\top0.svm0.counter[1] ),
    .C(_02574_),
    .X(_02577_));
 sky130_fd_sc_hd__or3b_1 _23077_ (.A(net64),
    .B(_02352_),
    .C_N(_02574_),
    .X(_02578_));
 sky130_fd_sc_hd__a211o_1 _23078_ (.A1(_02577_),
    .A2(_02578_),
    .B1(_02298_),
    .C1(net65),
    .X(_02579_));
 sky130_fd_sc_hd__xnor2_1 _23079_ (.A(_02339_),
    .B(_02538_),
    .Y(_02580_));
 sky130_fd_sc_hd__nor2_1 _23080_ (.A(_05735_),
    .B(_02580_),
    .Y(_02581_));
 sky130_fd_sc_hd__and3_1 _23081_ (.A(_05735_),
    .B(_02339_),
    .C(_02538_),
    .X(_02582_));
 sky130_fd_sc_hd__xnor2_1 _23082_ (.A(\top0.periodTop_r[4] ),
    .B(\top0.svm0.counter[4] ),
    .Y(_02583_));
 sky130_fd_sc_hd__o21ai_1 _23083_ (.A1(_02581_),
    .A2(_02582_),
    .B1(_02583_),
    .Y(_02584_));
 sky130_fd_sc_hd__or3_1 _23084_ (.A(_02339_),
    .B(_02539_),
    .C(_02583_),
    .X(_02585_));
 sky130_fd_sc_hd__a22oi_1 _23085_ (.A1(net170),
    .A2(_02567_),
    .B1(_02568_),
    .B2(_02566_),
    .Y(_02586_));
 sky130_fd_sc_hd__a221o_1 _23086_ (.A1(_02576_),
    .A2(_02579_),
    .B1(_02584_),
    .B2(_02585_),
    .C1(_02586_),
    .X(_02587_));
 sky130_fd_sc_hd__xor2_1 _23087_ (.A(net36),
    .B(\top0.svm0.counter[11] ),
    .X(_02588_));
 sky130_fd_sc_hd__xnor2_1 _23088_ (.A(_02542_),
    .B(_02588_),
    .Y(_02589_));
 sky130_fd_sc_hd__xor2_1 _23089_ (.A(net40),
    .B(net169),
    .X(_02590_));
 sky130_fd_sc_hd__xnor2_1 _23090_ (.A(_02541_),
    .B(_02590_),
    .Y(_02591_));
 sky130_fd_sc_hd__or4_1 _23091_ (.A(_02573_),
    .B(_02587_),
    .C(_02589_),
    .D(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__a2111oi_1 _23092_ (.A1(_02548_),
    .A2(_02549_),
    .B1(_02556_),
    .C1(_02563_),
    .D1(_02592_),
    .Y(_02593_));
 sky130_fd_sc_hd__a21o_1 _23093_ (.A1(\top0.svm0.rising ),
    .A2(net9),
    .B1(_02305_),
    .X(_02594_));
 sky130_fd_sc_hd__o21a_2 _23094_ (.A1(net171),
    .A2(_07114_),
    .B1(_02594_),
    .X(_02595_));
 sky130_fd_sc_hd__buf_2 _23095_ (.A(_02595_),
    .X(_02596_));
 sky130_fd_sc_hd__o21ai_1 _23096_ (.A1(net555),
    .A2(_02483_),
    .B1(_02596_),
    .Y(_02597_));
 sky130_fd_sc_hd__and3_2 _23097_ (.A(net171),
    .B(_02306_),
    .C(_02594_),
    .X(_02598_));
 sky130_fd_sc_hd__and3b_1 _23098_ (.A_N(\top0.svm0.delta[1] ),
    .B(net555),
    .C(_02598_),
    .X(_02599_));
 sky130_fd_sc_hd__a21o_1 _23099_ (.A1(\top0.svm0.delta[1] ),
    .A2(_02597_),
    .B1(_02599_),
    .X(_00458_));
 sky130_fd_sc_hd__o31ai_1 _23100_ (.A1(\top0.svm0.delta[1] ),
    .A2(net555),
    .A3(_02440_),
    .B1(_02596_),
    .Y(_02600_));
 sky130_fd_sc_hd__o211a_1 _23101_ (.A1(\top0.svm0.delta[1] ),
    .A2(net555),
    .B1(_02443_),
    .C1(_02598_),
    .X(_02601_));
 sky130_fd_sc_hd__a21o_1 _23102_ (.A1(net896),
    .A2(_02600_),
    .B1(_02601_),
    .X(_00459_));
 sky130_fd_sc_hd__o31a_1 _23103_ (.A1(\top0.svm0.delta[1] ),
    .A2(net555),
    .A3(\top0.svm0.delta[2] ),
    .B1(_02595_),
    .X(_02602_));
 sky130_fd_sc_hd__xnor2_1 _23104_ (.A(\top0.svm0.delta[3] ),
    .B(_02602_),
    .Y(_02603_));
 sky130_fd_sc_hd__nor2_1 _23105_ (.A(_07117_),
    .B(_02603_),
    .Y(_00460_));
 sky130_fd_sc_hd__or4_2 _23106_ (.A(\top0.svm0.delta[1] ),
    .B(net555),
    .C(\top0.svm0.delta[2] ),
    .D(\top0.svm0.delta[3] ),
    .X(_02604_));
 sky130_fd_sc_hd__or2_1 _23107_ (.A(_02440_),
    .B(_02604_),
    .X(_02605_));
 sky130_fd_sc_hd__a21oi_1 _23108_ (.A1(_02596_),
    .A2(_02605_),
    .B1(_02458_),
    .Y(_02606_));
 sky130_fd_sc_hd__a31o_1 _23109_ (.A1(_02458_),
    .A2(_02598_),
    .A3(_02604_),
    .B1(_02606_),
    .X(_00461_));
 sky130_fd_sc_hd__o21a_1 _23110_ (.A1(\top0.svm0.delta[4] ),
    .A2(_02604_),
    .B1(_02595_),
    .X(_02607_));
 sky130_fd_sc_hd__xnor2_1 _23111_ (.A(\top0.svm0.delta[5] ),
    .B(_02607_),
    .Y(_02608_));
 sky130_fd_sc_hd__nor2_1 _23112_ (.A(_07117_),
    .B(_02608_),
    .Y(_00462_));
 sky130_fd_sc_hd__or3_1 _23113_ (.A(\top0.svm0.delta[4] ),
    .B(\top0.svm0.delta[5] ),
    .C(_02604_),
    .X(_02609_));
 sky130_fd_sc_hd__o21ai_1 _23114_ (.A1(_02483_),
    .A2(_02609_),
    .B1(_02596_),
    .Y(_02610_));
 sky130_fd_sc_hd__and3_1 _23115_ (.A(_02478_),
    .B(_02598_),
    .C(_02609_),
    .X(_02611_));
 sky130_fd_sc_hd__a21o_1 _23116_ (.A1(net955),
    .A2(_02610_),
    .B1(_02611_),
    .X(_00463_));
 sky130_fd_sc_hd__or2_1 _23117_ (.A(\top0.svm0.delta[6] ),
    .B(_02609_),
    .X(_02612_));
 sky130_fd_sc_hd__o21ai_1 _23118_ (.A1(_02483_),
    .A2(_02612_),
    .B1(_02596_),
    .Y(_02613_));
 sky130_fd_sc_hd__and3_1 _23119_ (.A(_02485_),
    .B(_02598_),
    .C(_02612_),
    .X(_02614_));
 sky130_fd_sc_hd__a21o_1 _23120_ (.A1(net933),
    .A2(_02613_),
    .B1(_02614_),
    .X(_00464_));
 sky130_fd_sc_hd__o21a_1 _23121_ (.A1(\top0.svm0.delta[7] ),
    .A2(_02612_),
    .B1(_02595_),
    .X(_02615_));
 sky130_fd_sc_hd__xnor2_1 _23122_ (.A(\top0.svm0.delta[8] ),
    .B(_02615_),
    .Y(_02616_));
 sky130_fd_sc_hd__nor2_1 _23123_ (.A(_07117_),
    .B(_02616_),
    .Y(_00465_));
 sky130_fd_sc_hd__o31a_1 _23124_ (.A1(\top0.svm0.delta[7] ),
    .A2(\top0.svm0.delta[8] ),
    .A3(_02612_),
    .B1(_02595_),
    .X(_02617_));
 sky130_fd_sc_hd__xnor2_1 _23125_ (.A(\top0.svm0.delta[9] ),
    .B(_02617_),
    .Y(_02618_));
 sky130_fd_sc_hd__nor2_1 _23126_ (.A(_07117_),
    .B(_02618_),
    .Y(_00466_));
 sky130_fd_sc_hd__or4_1 _23127_ (.A(\top0.svm0.delta[7] ),
    .B(\top0.svm0.delta[8] ),
    .C(\top0.svm0.delta[9] ),
    .D(_02612_),
    .X(_02619_));
 sky130_fd_sc_hd__nand2_1 _23128_ (.A(_02596_),
    .B(_02619_),
    .Y(_02620_));
 sky130_fd_sc_hd__xor2_1 _23129_ (.A(\top0.svm0.delta[10] ),
    .B(_02620_),
    .X(_02621_));
 sky130_fd_sc_hd__nor2_1 _23130_ (.A(_07117_),
    .B(_02621_),
    .Y(_00467_));
 sky130_fd_sc_hd__or2_1 _23131_ (.A(\top0.svm0.delta[10] ),
    .B(_02619_),
    .X(_02622_));
 sky130_fd_sc_hd__o21ai_1 _23132_ (.A1(_02483_),
    .A2(_02622_),
    .B1(_02596_),
    .Y(_02623_));
 sky130_fd_sc_hd__and3_1 _23133_ (.A(_02508_),
    .B(_02598_),
    .C(_02622_),
    .X(_02624_));
 sky130_fd_sc_hd__a21o_1 _23134_ (.A1(net959),
    .A2(_02623_),
    .B1(_02624_),
    .X(_00468_));
 sky130_fd_sc_hd__or2_1 _23135_ (.A(\top0.svm0.delta[11] ),
    .B(_02622_),
    .X(_02625_));
 sky130_fd_sc_hd__o21ai_1 _23136_ (.A1(_02483_),
    .A2(_02625_),
    .B1(_02596_),
    .Y(_02626_));
 sky130_fd_sc_hd__and3_1 _23137_ (.A(_02514_),
    .B(_02598_),
    .C(_02625_),
    .X(_02627_));
 sky130_fd_sc_hd__a21o_1 _23138_ (.A1(net972),
    .A2(_02626_),
    .B1(_02627_),
    .X(_00469_));
 sky130_fd_sc_hd__or2_1 _23139_ (.A(\top0.svm0.delta[12] ),
    .B(_02625_),
    .X(_02628_));
 sky130_fd_sc_hd__and2_1 _23140_ (.A(_02598_),
    .B(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__o21ai_1 _23141_ (.A1(_02440_),
    .A2(_02628_),
    .B1(_02596_),
    .Y(_02630_));
 sky130_fd_sc_hd__mux2_1 _23142_ (.A0(_02629_),
    .A1(_02630_),
    .S(\top0.svm0.delta[13] ),
    .X(_02631_));
 sky130_fd_sc_hd__clkbuf_1 _23143_ (.A(_02631_),
    .X(_00470_));
 sky130_fd_sc_hd__or2_1 _23144_ (.A(\top0.svm0.delta[13] ),
    .B(_02628_),
    .X(_02632_));
 sky130_fd_sc_hd__and2_1 _23145_ (.A(_02598_),
    .B(_02632_),
    .X(_02633_));
 sky130_fd_sc_hd__o21ai_1 _23146_ (.A1(_02440_),
    .A2(_02632_),
    .B1(_02596_),
    .Y(_02634_));
 sky130_fd_sc_hd__mux2_1 _23147_ (.A0(_02633_),
    .A1(_02634_),
    .S(\top0.svm0.delta[14] ),
    .X(_02635_));
 sky130_fd_sc_hd__clkbuf_1 _23148_ (.A(_02635_),
    .X(_00471_));
 sky130_fd_sc_hd__o21ai_1 _23149_ (.A1(\top0.svm0.delta[14] ),
    .A2(_02632_),
    .B1(_02595_),
    .Y(_02636_));
 sky130_fd_sc_hd__nand2_1 _23150_ (.A(\top0.svm0.delta[15] ),
    .B(_02636_),
    .Y(_02637_));
 sky130_fd_sc_hd__or2_1 _23151_ (.A(\top0.svm0.delta[15] ),
    .B(_02636_),
    .X(_02638_));
 sky130_fd_sc_hd__a21oi_1 _23152_ (.A1(_02637_),
    .A2(_02638_),
    .B1(_07117_),
    .Y(_00472_));
 sky130_fd_sc_hd__nand2_1 _23153_ (.A(net171),
    .B(_02305_),
    .Y(_02639_));
 sky130_fd_sc_hd__a21bo_1 _23154_ (.A1(net171),
    .A2(net9),
    .B1_N(\top0.svm0.rising ),
    .X(_02640_));
 sky130_fd_sc_hd__nand2_1 _23155_ (.A(_02639_),
    .B(_02640_),
    .Y(_00473_));
 sky130_fd_sc_hd__o21a_1 _23156_ (.A1(net902),
    .A2(_06381_),
    .B1(_02639_),
    .X(_00474_));
 sky130_fd_sc_hd__clkbuf_4 _23157_ (.A(_05717_),
    .X(_02641_));
 sky130_fd_sc_hd__inv_2 _23158_ (.A(\top0.svm0.state[1] ),
    .Y(_02642_));
 sky130_fd_sc_hd__mux2_1 _23159_ (.A0(_07115_),
    .A1(_02308_),
    .S(_02642_),
    .X(_02643_));
 sky130_fd_sc_hd__buf_6 _23160_ (.A(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__clkbuf_4 _23161_ (.A(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__a22o_1 _23162_ (.A1(_02641_),
    .A2(_06275_),
    .B1(_02645_),
    .B2(net830),
    .X(_00475_));
 sky130_fd_sc_hd__a22o_1 _23163_ (.A1(_02641_),
    .A2(_06380_),
    .B1(_02645_),
    .B2(net795),
    .X(_00476_));
 sky130_fd_sc_hd__a22o_1 _23164_ (.A1(_02641_),
    .A2(_06473_),
    .B1(_02645_),
    .B2(net783),
    .X(_00477_));
 sky130_fd_sc_hd__a22o_1 _23165_ (.A1(_02641_),
    .A2(_06546_),
    .B1(_02645_),
    .B2(net811),
    .X(_00478_));
 sky130_fd_sc_hd__a22o_1 _23166_ (.A1(_02641_),
    .A2(_06612_),
    .B1(_02645_),
    .B2(net883),
    .X(_00479_));
 sky130_fd_sc_hd__a22o_1 _23167_ (.A1(_02641_),
    .A2(_06682_),
    .B1(_02645_),
    .B2(net894),
    .X(_00480_));
 sky130_fd_sc_hd__a22o_1 _23168_ (.A1(_02641_),
    .A2(_06748_),
    .B1(_02645_),
    .B2(net780),
    .X(_00481_));
 sky130_fd_sc_hd__a22o_1 _23169_ (.A1(_02641_),
    .A2(_06799_),
    .B1(_02645_),
    .B2(net788),
    .X(_00482_));
 sky130_fd_sc_hd__a22o_1 _23170_ (.A1(_02641_),
    .A2(_06860_),
    .B1(_02645_),
    .B2(net930),
    .X(_00483_));
 sky130_fd_sc_hd__a22o_1 _23171_ (.A1(_02641_),
    .A2(_06907_),
    .B1(_02645_),
    .B2(net989),
    .X(_00484_));
 sky130_fd_sc_hd__a22o_1 _23172_ (.A1(_05717_),
    .A2(_06945_),
    .B1(_02644_),
    .B2(net781),
    .X(_00485_));
 sky130_fd_sc_hd__a22o_1 _23173_ (.A1(_05717_),
    .A2(_06971_),
    .B1(_02644_),
    .B2(net806),
    .X(_00486_));
 sky130_fd_sc_hd__a22o_1 _23174_ (.A1(_05717_),
    .A2(_07000_),
    .B1(_02644_),
    .B2(net882),
    .X(_00487_));
 sky130_fd_sc_hd__a22o_1 _23175_ (.A1(_05717_),
    .A2(_07028_),
    .B1(_02644_),
    .B2(net777),
    .X(_00488_));
 sky130_fd_sc_hd__a22o_1 _23176_ (.A1(_05717_),
    .A2(_07034_),
    .B1(_02644_),
    .B2(net908),
    .X(_00489_));
 sky130_fd_sc_hd__a22o_1 _23177_ (.A1(_05717_),
    .A2(_07038_),
    .B1(_02644_),
    .B2(net800),
    .X(_00490_));
 sky130_fd_sc_hd__clkbuf_4 _23178_ (.A(_05719_),
    .X(_02646_));
 sky130_fd_sc_hd__mux2_1 _23179_ (.A0(_07115_),
    .A1(_02642_),
    .S(_02308_),
    .X(_02647_));
 sky130_fd_sc_hd__buf_6 _23180_ (.A(_02647_),
    .X(_02648_));
 sky130_fd_sc_hd__clkbuf_4 _23181_ (.A(_02648_),
    .X(_02649_));
 sky130_fd_sc_hd__a22o_1 _23182_ (.A1(_02646_),
    .A2(_06275_),
    .B1(_02649_),
    .B2(net729),
    .X(_00491_));
 sky130_fd_sc_hd__a22o_1 _23183_ (.A1(_02646_),
    .A2(_06380_),
    .B1(_02649_),
    .B2(net831),
    .X(_00492_));
 sky130_fd_sc_hd__a22o_1 _23184_ (.A1(_02646_),
    .A2(_06473_),
    .B1(_02649_),
    .B2(net835),
    .X(_00493_));
 sky130_fd_sc_hd__a22o_1 _23185_ (.A1(_02646_),
    .A2(_06546_),
    .B1(_02649_),
    .B2(net837),
    .X(_00494_));
 sky130_fd_sc_hd__a22o_1 _23186_ (.A1(_02646_),
    .A2(_06612_),
    .B1(_02649_),
    .B2(net823),
    .X(_00495_));
 sky130_fd_sc_hd__a22o_1 _23187_ (.A1(_02646_),
    .A2(_06682_),
    .B1(_02649_),
    .B2(net821),
    .X(_00496_));
 sky130_fd_sc_hd__a22o_1 _23188_ (.A1(_02646_),
    .A2(_06748_),
    .B1(_02649_),
    .B2(net834),
    .X(_00497_));
 sky130_fd_sc_hd__a22o_1 _23189_ (.A1(_02646_),
    .A2(_06799_),
    .B1(_02649_),
    .B2(net776),
    .X(_00498_));
 sky130_fd_sc_hd__a22o_1 _23190_ (.A1(_02646_),
    .A2(_06860_),
    .B1(_02649_),
    .B2(net814),
    .X(_00499_));
 sky130_fd_sc_hd__a22o_1 _23191_ (.A1(_02646_),
    .A2(_06907_),
    .B1(_02649_),
    .B2(net797),
    .X(_00500_));
 sky130_fd_sc_hd__a22o_1 _23192_ (.A1(_05719_),
    .A2(_06945_),
    .B1(_02648_),
    .B2(net774),
    .X(_00501_));
 sky130_fd_sc_hd__a22o_1 _23193_ (.A1(_05719_),
    .A2(_06971_),
    .B1(_02648_),
    .B2(net790),
    .X(_00502_));
 sky130_fd_sc_hd__a22o_1 _23194_ (.A1(_05719_),
    .A2(_07000_),
    .B1(_02648_),
    .B2(net809),
    .X(_00503_));
 sky130_fd_sc_hd__a22o_1 _23195_ (.A1(_05719_),
    .A2(_07028_),
    .B1(_02648_),
    .B2(net804),
    .X(_00504_));
 sky130_fd_sc_hd__a22o_1 _23196_ (.A1(_05719_),
    .A2(_07034_),
    .B1(_02648_),
    .B2(net838),
    .X(_00505_));
 sky130_fd_sc_hd__a22o_1 _23197_ (.A1(_05719_),
    .A2(_07038_),
    .B1(_02648_),
    .B2(net839),
    .X(_00506_));
 sky130_fd_sc_hd__mux4_2 _23198_ (.A0(net243),
    .A1(net237),
    .A2(net233),
    .A3(net228),
    .S0(net204),
    .S1(net196),
    .X(_02650_));
 sky130_fd_sc_hd__mux4_1 _23199_ (.A0(net260),
    .A1(net254),
    .A2(net251),
    .A3(net245),
    .S0(net204),
    .S1(net196),
    .X(_02651_));
 sky130_fd_sc_hd__mux2_1 _23200_ (.A0(_02650_),
    .A1(_02651_),
    .S(_11572_),
    .X(_02652_));
 sky130_fd_sc_hd__mux4_1 _23201_ (.A0(net297),
    .A1(net291),
    .A2(net272),
    .A3(net266),
    .S0(net197),
    .S1(net188),
    .X(_02653_));
 sky130_fd_sc_hd__mux4_1 _23202_ (.A0(net306),
    .A1(net300),
    .A2(net286),
    .A3(net277),
    .S0(net197),
    .S1(net188),
    .X(_02654_));
 sky130_fd_sc_hd__mux2_1 _23203_ (.A0(_02653_),
    .A1(_02654_),
    .S(_11409_),
    .X(_02655_));
 sky130_fd_sc_hd__mux2_1 _23204_ (.A0(_02652_),
    .A1(_02655_),
    .S(_11420_),
    .X(_02656_));
 sky130_fd_sc_hd__mux2_2 _23205_ (.A0(net223),
    .A1(net217),
    .S(net203),
    .X(_02657_));
 sky130_fd_sc_hd__mux2_1 _23206_ (.A0(_02657_),
    .A1(net217),
    .S(_11775_),
    .X(_02658_));
 sky130_fd_sc_hd__mux2_1 _23207_ (.A0(_02656_),
    .A1(_02658_),
    .S(net179),
    .X(_02659_));
 sky130_fd_sc_hd__buf_2 _23208_ (.A(_02659_),
    .X(_02660_));
 sky130_fd_sc_hd__o21a_1 _23209_ (.A1(_11526_),
    .A2(_02660_),
    .B1(net174),
    .X(_02661_));
 sky130_fd_sc_hd__nor2_1 _23210_ (.A(_01320_),
    .B(_02661_),
    .Y(_02662_));
 sky130_fd_sc_hd__a31o_1 _23211_ (.A1(_01320_),
    .A2(net1013),
    .A3(_02660_),
    .B1(_02662_),
    .X(_00507_));
 sky130_fd_sc_hd__mux4_2 _23212_ (.A0(net237),
    .A1(net233),
    .A2(net228),
    .A3(net223),
    .S0(net204),
    .S1(net196),
    .X(_02663_));
 sky130_fd_sc_hd__mux4_2 _23213_ (.A0(net254),
    .A1(net250),
    .A2(net244),
    .A3(net243),
    .S0(net198),
    .S1(net192),
    .X(_02664_));
 sky130_fd_sc_hd__mux4_1 _23214_ (.A0(net279),
    .A1(net272),
    .A2(net266),
    .A3(net260),
    .S0(net198),
    .S1(net191),
    .X(_02665_));
 sky130_fd_sc_hd__mux4_1 _23215_ (.A0(net301),
    .A1(net297),
    .A2(net292),
    .A3(net286),
    .S0(net198),
    .S1(net191),
    .X(_02666_));
 sky130_fd_sc_hd__mux4_1 _23216_ (.A0(_02663_),
    .A1(_02664_),
    .A2(_02665_),
    .A3(_02666_),
    .S0(_11572_),
    .S1(_11576_),
    .X(_02667_));
 sky130_fd_sc_hd__nand2_1 _23217_ (.A(net179),
    .B(net215),
    .Y(_02668_));
 sky130_fd_sc_hd__a21bo_2 _23218_ (.A1(_11425_),
    .A2(_02667_),
    .B1_N(_02668_),
    .X(_02669_));
 sky130_fd_sc_hd__nor2_1 _23219_ (.A(_01320_),
    .B(_11515_),
    .Y(_02670_));
 sky130_fd_sc_hd__nor2_1 _23220_ (.A(net165),
    .B(_11519_),
    .Y(_02671_));
 sky130_fd_sc_hd__o21a_1 _23221_ (.A1(_02670_),
    .A2(_02671_),
    .B1(_02660_),
    .X(_02672_));
 sky130_fd_sc_hd__xnor2_1 _23222_ (.A(_02669_),
    .B(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hd__a21o_1 _23223_ (.A1(_11650_),
    .A2(_02673_),
    .B1(net1020),
    .X(_02674_));
 sky130_fd_sc_hd__or3_1 _23224_ (.A(net160),
    .B(_11784_),
    .C(_02673_),
    .X(_02675_));
 sky130_fd_sc_hd__a21bo_1 _23225_ (.A1(net161),
    .A2(_02674_),
    .B1_N(_02675_),
    .X(_00508_));
 sky130_fd_sc_hd__or3b_1 _23226_ (.A(_01267_),
    .B(_02669_),
    .C_N(_02660_),
    .X(_02676_));
 sky130_fd_sc_hd__nand2_1 _23227_ (.A(net161),
    .B(_02669_),
    .Y(_02677_));
 sky130_fd_sc_hd__mux2_1 _23228_ (.A0(_02676_),
    .A1(_02677_),
    .S(net1016),
    .X(_02678_));
 sky130_fd_sc_hd__a21boi_2 _23229_ (.A1(_11425_),
    .A2(_02667_),
    .B1_N(_02668_),
    .Y(_02679_));
 sky130_fd_sc_hd__or3b_1 _23230_ (.A(_02679_),
    .B(_01320_),
    .C_N(_02659_),
    .X(_02680_));
 sky130_fd_sc_hd__or3b_1 _23231_ (.A(_01320_),
    .B(_02669_),
    .C_N(_02659_),
    .X(_02681_));
 sky130_fd_sc_hd__mux2_1 _23232_ (.A0(_02680_),
    .A1(_02681_),
    .S(_11511_),
    .X(_02682_));
 sky130_fd_sc_hd__nor2_1 _23233_ (.A(_01320_),
    .B(_01267_),
    .Y(_02683_));
 sky130_fd_sc_hd__nand2_1 _23234_ (.A(_02683_),
    .B(_02660_),
    .Y(_02684_));
 sky130_fd_sc_hd__or3_1 _23235_ (.A(_01267_),
    .B(_02660_),
    .C(_02679_),
    .X(_02685_));
 sky130_fd_sc_hd__nand4_2 _23236_ (.A(_02678_),
    .B(_02682_),
    .C(_02684_),
    .D(_02685_),
    .Y(_02686_));
 sky130_fd_sc_hd__mux4_2 _23237_ (.A0(net233),
    .A1(net228),
    .A2(net223),
    .A3(net220),
    .S0(net203),
    .S1(net196),
    .X(_02687_));
 sky130_fd_sc_hd__mux4_2 _23238_ (.A0(net249),
    .A1(net244),
    .A2(net243),
    .A3(net237),
    .S0(net198),
    .S1(net192),
    .X(_02688_));
 sky130_fd_sc_hd__mux4_1 _23239_ (.A0(net272),
    .A1(net266),
    .A2(net260),
    .A3(net254),
    .S0(net198),
    .S1(net192),
    .X(_02689_));
 sky130_fd_sc_hd__mux4_1 _23240_ (.A0(net297),
    .A1(net291),
    .A2(net286),
    .A3(net279),
    .S0(net198),
    .S1(net192),
    .X(_02690_));
 sky130_fd_sc_hd__mux4_1 _23241_ (.A0(_02687_),
    .A1(_02688_),
    .A2(_02689_),
    .A3(_02690_),
    .S0(_11572_),
    .S1(_11420_),
    .X(_02691_));
 sky130_fd_sc_hd__a21bo_1 _23242_ (.A1(_11425_),
    .A2(_02691_),
    .B1_N(_02668_),
    .X(_02692_));
 sky130_fd_sc_hd__nor2_1 _23243_ (.A(_02660_),
    .B(_02669_),
    .Y(_02693_));
 sky130_fd_sc_hd__a211o_1 _23244_ (.A1(_11484_),
    .A2(_11504_),
    .B1(_11509_),
    .C1(_02693_),
    .X(_02694_));
 sky130_fd_sc_hd__xnor2_2 _23245_ (.A(_02692_),
    .B(_02694_),
    .Y(_02695_));
 sky130_fd_sc_hd__xnor2_1 _23246_ (.A(_02686_),
    .B(_02695_),
    .Y(_02696_));
 sky130_fd_sc_hd__nor2_1 _23247_ (.A(_11857_),
    .B(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__a21o_1 _23248_ (.A1(_11649_),
    .A2(_02696_),
    .B1(_11954_),
    .X(_02698_));
 sky130_fd_sc_hd__mux2_1 _23249_ (.A0(_02697_),
    .A1(_02698_),
    .S(net156),
    .X(_02699_));
 sky130_fd_sc_hd__clkbuf_1 _23250_ (.A(_02699_),
    .X(_00509_));
 sky130_fd_sc_hd__a21oi_1 _23251_ (.A1(_11511_),
    .A2(_02660_),
    .B1(_02677_),
    .Y(_02700_));
 sky130_fd_sc_hd__or2_1 _23252_ (.A(net155),
    .B(_02700_),
    .X(_02701_));
 sky130_fd_sc_hd__and3_1 _23253_ (.A(net165),
    .B(net1016),
    .C(_02669_),
    .X(_02702_));
 sky130_fd_sc_hd__and3_1 _23254_ (.A(net161),
    .B(_11511_),
    .C(_02679_),
    .X(_02703_));
 sky130_fd_sc_hd__a31o_1 _23255_ (.A1(net165),
    .A2(_11511_),
    .A3(_02679_),
    .B1(_02683_),
    .X(_02704_));
 sky130_fd_sc_hd__o31a_1 _23256_ (.A1(_02702_),
    .A2(_02703_),
    .A3(_02704_),
    .B1(_02660_),
    .X(_02705_));
 sky130_fd_sc_hd__or2_1 _23257_ (.A(net155),
    .B(_02695_),
    .X(_02706_));
 sky130_fd_sc_hd__o221a_1 _23258_ (.A1(_02686_),
    .A2(_02695_),
    .B1(_02701_),
    .B2(_02705_),
    .C1(_02706_),
    .X(_02707_));
 sky130_fd_sc_hd__and2b_1 _23259_ (.A_N(_02692_),
    .B(_02693_),
    .X(_02708_));
 sky130_fd_sc_hd__mux4_1 _23260_ (.A0(net268),
    .A1(net259),
    .A2(net254),
    .A3(net251),
    .S0(net204),
    .S1(net196),
    .X(_02709_));
 sky130_fd_sc_hd__mux4_1 _23261_ (.A0(net291),
    .A1(net286),
    .A2(net278),
    .A3(net272),
    .S0(net198),
    .S1(net192),
    .X(_02710_));
 sky130_fd_sc_hd__mux2_1 _23262_ (.A0(net228),
    .A1(net223),
    .S(net203),
    .X(_02711_));
 sky130_fd_sc_hd__a22o_1 _23263_ (.A1(net215),
    .A2(_11633_),
    .B1(_02711_),
    .B2(_11409_),
    .X(_02712_));
 sky130_fd_sc_hd__mux4_2 _23264_ (.A0(net244),
    .A1(net243),
    .A2(net237),
    .A3(net233),
    .S0(net204),
    .S1(net196),
    .X(_02713_));
 sky130_fd_sc_hd__mux4_1 _23265_ (.A0(_02709_),
    .A1(_02710_),
    .A2(_02712_),
    .A3(_02713_),
    .S0(_11572_),
    .S1(net182),
    .X(_02714_));
 sky130_fd_sc_hd__o21a_1 _23266_ (.A1(net180),
    .A2(_02289_),
    .B1(net215),
    .X(_02715_));
 sky130_fd_sc_hd__a21oi_1 _23267_ (.A1(_11425_),
    .A2(_02714_),
    .B1(_02715_),
    .Y(_02716_));
 sky130_fd_sc_hd__o21ai_1 _23268_ (.A1(net1016),
    .A2(_02708_),
    .B1(_02716_),
    .Y(_02717_));
 sky130_fd_sc_hd__or3_1 _23269_ (.A(net1016),
    .B(_02716_),
    .C(_02708_),
    .X(_02718_));
 sky130_fd_sc_hd__and2_1 _23270_ (.A(_02717_),
    .B(_02718_),
    .X(_02719_));
 sky130_fd_sc_hd__and2_1 _23271_ (.A(_02707_),
    .B(_02719_),
    .X(_02720_));
 sky130_fd_sc_hd__or2_1 _23272_ (.A(_02707_),
    .B(_02719_),
    .X(_02721_));
 sky130_fd_sc_hd__and2b_1 _23273_ (.A_N(_02720_),
    .B(_02721_),
    .X(_02722_));
 sky130_fd_sc_hd__o21ai_1 _23274_ (.A1(net1014),
    .A2(_02722_),
    .B1(net176),
    .Y(_02723_));
 sky130_fd_sc_hd__nor2_1 _23275_ (.A(net150),
    .B(_11857_),
    .Y(_02724_));
 sky130_fd_sc_hd__a22o_1 _23276_ (.A1(net150),
    .A2(_02723_),
    .B1(_02724_),
    .B2(_02722_),
    .X(_00510_));
 sky130_fd_sc_hd__a21oi_2 _23277_ (.A1(net150),
    .A2(_02721_),
    .B1(_02720_),
    .Y(_02725_));
 sky130_fd_sc_hd__mux4_1 _23278_ (.A0(net286),
    .A1(net278),
    .A2(net272),
    .A3(net265),
    .S0(net204),
    .S1(net196),
    .X(_02726_));
 sky130_fd_sc_hd__mux2_1 _23279_ (.A0(_02651_),
    .A1(_02726_),
    .S(_11572_),
    .X(_02727_));
 sky130_fd_sc_hd__or2_1 _23280_ (.A(net182),
    .B(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__a221o_1 _23281_ (.A1(_11572_),
    .A2(_02650_),
    .B1(_02657_),
    .B2(_11574_),
    .C1(_11576_),
    .X(_02729_));
 sky130_fd_sc_hd__a32o_1 _23282_ (.A1(_11425_),
    .A2(_02728_),
    .A3(_02729_),
    .B1(net215),
    .B2(_11580_),
    .X(_02730_));
 sky130_fd_sc_hd__a211o_1 _23283_ (.A1(_11425_),
    .A2(_02714_),
    .B1(_02715_),
    .C1(_02692_),
    .X(_02731_));
 sky130_fd_sc_hd__nor3_1 _23284_ (.A(_02660_),
    .B(_02669_),
    .C(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__a211o_1 _23285_ (.A1(_11484_),
    .A2(_11504_),
    .B1(_11509_),
    .C1(_02732_),
    .X(_02733_));
 sky130_fd_sc_hd__xor2_2 _23286_ (.A(_02730_),
    .B(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__xnor2_1 _23287_ (.A(_02725_),
    .B(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__a21o_1 _23288_ (.A1(_11649_),
    .A2(_02735_),
    .B1(_11954_),
    .X(_02736_));
 sky130_fd_sc_hd__nor2_1 _23289_ (.A(_11784_),
    .B(_02735_),
    .Y(_02737_));
 sky130_fd_sc_hd__mux2_1 _23290_ (.A0(_02736_),
    .A1(_02737_),
    .S(_01102_),
    .X(_02738_));
 sky130_fd_sc_hd__clkbuf_1 _23291_ (.A(_02738_),
    .X(_00511_));
 sky130_fd_sc_hd__nor2_1 _23292_ (.A(_11788_),
    .B(_11427_),
    .Y(_02739_));
 sky130_fd_sc_hd__mux4_1 _23293_ (.A0(_02663_),
    .A1(_02665_),
    .A2(_02739_),
    .A3(_02664_),
    .S0(_11576_),
    .S1(net188),
    .X(_02740_));
 sky130_fd_sc_hd__a22o_2 _23294_ (.A1(net220),
    .A2(_11594_),
    .B1(_02740_),
    .B2(_11425_),
    .X(_02741_));
 sky130_fd_sc_hd__or4_1 _23295_ (.A(_02659_),
    .B(_02669_),
    .C(_02730_),
    .D(_02731_),
    .X(_02742_));
 sky130_fd_sc_hd__nand2_1 _23296_ (.A(_11512_),
    .B(_02742_),
    .Y(_02743_));
 sky130_fd_sc_hd__xnor2_2 _23297_ (.A(_02741_),
    .B(_02743_),
    .Y(_02744_));
 sky130_fd_sc_hd__o21a_1 _23298_ (.A1(_02725_),
    .A2(_02734_),
    .B1(_01102_),
    .X(_02745_));
 sky130_fd_sc_hd__a21oi_1 _23299_ (.A1(_02725_),
    .A2(_02734_),
    .B1(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__xnor2_1 _23300_ (.A(_02744_),
    .B(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__a21o_1 _23301_ (.A1(_11650_),
    .A2(_02747_),
    .B1(net1020),
    .X(_02748_));
 sky130_fd_sc_hd__or3_1 _23302_ (.A(net138),
    .B(_11784_),
    .C(_02747_),
    .X(_02749_));
 sky130_fd_sc_hd__a21bo_1 _23303_ (.A1(net138),
    .A2(_02748_),
    .B1_N(_02749_),
    .X(_00512_));
 sky130_fd_sc_hd__o22a_1 _23304_ (.A1(_11573_),
    .A2(net215),
    .B1(_11613_),
    .B2(_02687_),
    .X(_02750_));
 sky130_fd_sc_hd__mux2_1 _23305_ (.A0(_02688_),
    .A1(_02689_),
    .S(_11573_),
    .X(_02751_));
 sky130_fd_sc_hd__or2_1 _23306_ (.A(_11448_),
    .B(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__o221a_2 _23307_ (.A1(_11425_),
    .A2(net215),
    .B1(_02750_),
    .B2(_11576_),
    .C1(_02752_),
    .X(_02753_));
 sky130_fd_sc_hd__o21a_1 _23308_ (.A1(_02741_),
    .A2(_02742_),
    .B1(_11512_),
    .X(_02754_));
 sky130_fd_sc_hd__xor2_2 _23309_ (.A(_02753_),
    .B(_02754_),
    .X(_02755_));
 sky130_fd_sc_hd__o2111a_1 _23310_ (.A1(net140),
    .A2(_02744_),
    .B1(_02707_),
    .C1(net144),
    .D1(_02719_),
    .X(_02756_));
 sky130_fd_sc_hd__xnor2_1 _23311_ (.A(_11512_),
    .B(_02741_),
    .Y(_02757_));
 sky130_fd_sc_hd__a21oi_1 _23312_ (.A1(_01311_),
    .A2(_02757_),
    .B1(_02734_),
    .Y(_02758_));
 sky130_fd_sc_hd__o21a_1 _23313_ (.A1(net150),
    .A2(_02719_),
    .B1(_02758_),
    .X(_02759_));
 sky130_fd_sc_hd__a31o_1 _23314_ (.A1(net150),
    .A2(_02717_),
    .A3(_02718_),
    .B1(net145),
    .X(_02760_));
 sky130_fd_sc_hd__a22o_1 _23315_ (.A1(net140),
    .A2(_02744_),
    .B1(_02758_),
    .B2(_02760_),
    .X(_02761_));
 sky130_fd_sc_hd__a21o_1 _23316_ (.A1(_02707_),
    .A2(_02759_),
    .B1(_02761_),
    .X(_02762_));
 sky130_fd_sc_hd__o221a_1 _23317_ (.A1(_02707_),
    .A2(_02719_),
    .B1(_02744_),
    .B2(net140),
    .C1(_01123_),
    .X(_02763_));
 sky130_fd_sc_hd__or3_2 _23318_ (.A(_02756_),
    .B(_02762_),
    .C(_02763_),
    .X(_02764_));
 sky130_fd_sc_hd__xnor2_1 _23319_ (.A(_02755_),
    .B(_02764_),
    .Y(_02765_));
 sky130_fd_sc_hd__a21o_1 _23320_ (.A1(_11649_),
    .A2(_02765_),
    .B1(_11954_),
    .X(_02766_));
 sky130_fd_sc_hd__nor2_1 _23321_ (.A(_11784_),
    .B(_02765_),
    .Y(_02767_));
 sky130_fd_sc_hd__mux2_1 _23322_ (.A0(_02766_),
    .A1(_02767_),
    .S(_01105_),
    .X(_02768_));
 sky130_fd_sc_hd__clkbuf_1 _23323_ (.A(_02768_),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _23324_ (.A0(_02709_),
    .A1(_02713_),
    .S(net187),
    .X(_02769_));
 sky130_fd_sc_hd__a22o_1 _23325_ (.A1(_11876_),
    .A2(_02712_),
    .B1(_02769_),
    .B2(_11612_),
    .X(_02770_));
 sky130_fd_sc_hd__a22oi_4 _23326_ (.A1(net216),
    .A2(_11631_),
    .B1(_02770_),
    .B2(_11426_),
    .Y(_02771_));
 sky130_fd_sc_hd__nor3_1 _23327_ (.A(_02741_),
    .B(_02742_),
    .C(_02753_),
    .Y(_02772_));
 sky130_fd_sc_hd__nor2_1 _23328_ (.A(net1016),
    .B(_02772_),
    .Y(_02773_));
 sky130_fd_sc_hd__xnor2_2 _23329_ (.A(_02771_),
    .B(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__o21a_1 _23330_ (.A1(_02755_),
    .A2(_02764_),
    .B1(net133),
    .X(_02775_));
 sky130_fd_sc_hd__a21oi_1 _23331_ (.A1(_02755_),
    .A2(_02764_),
    .B1(_02775_),
    .Y(_02776_));
 sky130_fd_sc_hd__xnor2_1 _23332_ (.A(_02774_),
    .B(_02776_),
    .Y(_02777_));
 sky130_fd_sc_hd__o21a_1 _23333_ (.A1(_11526_),
    .A2(_02777_),
    .B1(net176),
    .X(_02778_));
 sky130_fd_sc_hd__nor2_1 _23334_ (.A(_01135_),
    .B(_02778_),
    .Y(_02779_));
 sky130_fd_sc_hd__a31o_1 _23335_ (.A1(_01135_),
    .A2(net1013),
    .A3(_02777_),
    .B1(_02779_),
    .X(_00514_));
 sky130_fd_sc_hd__and2_1 _23336_ (.A(net128),
    .B(_02774_),
    .X(_02780_));
 sky130_fd_sc_hd__or2_1 _23337_ (.A(_02755_),
    .B(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__or2_1 _23338_ (.A(net134),
    .B(_02780_),
    .X(_02782_));
 sky130_fd_sc_hd__a2111o_1 _23339_ (.A1(_02781_),
    .A2(_02782_),
    .B1(_02756_),
    .C1(_02762_),
    .D1(_02763_),
    .X(_02783_));
 sky130_fd_sc_hd__or3_1 _23340_ (.A(net134),
    .B(_02755_),
    .C(_02780_),
    .X(_02784_));
 sky130_fd_sc_hd__o211a_1 _23341_ (.A1(net128),
    .A2(_02774_),
    .B1(_02783_),
    .C1(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__a22o_1 _23342_ (.A1(net217),
    .A2(_11657_),
    .B1(_11658_),
    .B2(_02657_),
    .X(_02786_));
 sky130_fd_sc_hd__a21bo_1 _23343_ (.A1(net182),
    .A2(_02786_),
    .B1_N(_02668_),
    .X(_02787_));
 sky130_fd_sc_hd__a21o_2 _23344_ (.A1(_11560_),
    .A2(_02652_),
    .B1(_02787_),
    .X(_02788_));
 sky130_fd_sc_hd__nand2_1 _23345_ (.A(_02771_),
    .B(_02772_),
    .Y(_02789_));
 sky130_fd_sc_hd__nand2_2 _23346_ (.A(_11512_),
    .B(_02789_),
    .Y(_02790_));
 sky130_fd_sc_hd__xor2_4 _23347_ (.A(_02788_),
    .B(_02790_),
    .X(_02791_));
 sky130_fd_sc_hd__xnor2_1 _23348_ (.A(_02785_),
    .B(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__o21a_1 _23349_ (.A1(_11526_),
    .A2(_02792_),
    .B1(net176),
    .X(_02793_));
 sky130_fd_sc_hd__nor2_1 _23350_ (.A(_01408_),
    .B(_02793_),
    .Y(_02794_));
 sky130_fd_sc_hd__a31o_1 _23351_ (.A1(_01408_),
    .A2(_11548_),
    .A3(_02792_),
    .B1(_02794_),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _23352_ (.A0(_02663_),
    .A1(_02664_),
    .S(_11654_),
    .X(_02795_));
 sky130_fd_sc_hd__mux2_2 _23353_ (.A0(net216),
    .A1(_02795_),
    .S(_11560_),
    .X(_02796_));
 sky130_fd_sc_hd__or2_1 _23354_ (.A(_02788_),
    .B(_02789_),
    .X(_02797_));
 sky130_fd_sc_hd__nand2_1 _23355_ (.A(_11513_),
    .B(_02797_),
    .Y(_02798_));
 sky130_fd_sc_hd__xnor2_1 _23356_ (.A(_02796_),
    .B(_02798_),
    .Y(_02799_));
 sky130_fd_sc_hd__inv_2 _23357_ (.A(_02785_),
    .Y(_02800_));
 sky130_fd_sc_hd__o21a_1 _23358_ (.A1(_02800_),
    .A2(_02791_),
    .B1(_01408_),
    .X(_02801_));
 sky130_fd_sc_hd__a21oi_1 _23359_ (.A1(_02800_),
    .A2(_02791_),
    .B1(_02801_),
    .Y(_02802_));
 sky130_fd_sc_hd__xnor2_1 _23360_ (.A(_02799_),
    .B(_02802_),
    .Y(_02803_));
 sky130_fd_sc_hd__a21o_1 _23361_ (.A1(_11650_),
    .A2(_02803_),
    .B1(net1020),
    .X(_02804_));
 sky130_fd_sc_hd__or3_1 _23362_ (.A(net120),
    .B(_11783_),
    .C(_02803_),
    .X(_02805_));
 sky130_fd_sc_hd__a21bo_1 _23363_ (.A1(net120),
    .A2(_02804_),
    .B1_N(_02805_),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _23364_ (.A0(_02687_),
    .A1(_02688_),
    .S(_11654_),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_1 _23365_ (.A0(net216),
    .A1(_02806_),
    .S(_11560_),
    .X(_02807_));
 sky130_fd_sc_hd__o21ai_1 _23366_ (.A1(_02796_),
    .A2(_02797_),
    .B1(_11513_),
    .Y(_02808_));
 sky130_fd_sc_hd__xnor2_2 _23367_ (.A(_02807_),
    .B(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__inv_2 _23368_ (.A(_02809_),
    .Y(_02810_));
 sky130_fd_sc_hd__nand2_1 _23369_ (.A(_11518_),
    .B(_02796_),
    .Y(_02811_));
 sky130_fd_sc_hd__or2_1 _23370_ (.A(_11518_),
    .B(_02796_),
    .X(_02812_));
 sky130_fd_sc_hd__a31o_1 _23371_ (.A1(_01217_),
    .A2(_02811_),
    .A3(_02812_),
    .B1(_01408_),
    .X(_02813_));
 sky130_fd_sc_hd__a2bb2o_1 _23372_ (.A1_N(_02791_),
    .A2_N(_02813_),
    .B1(_02799_),
    .B2(net120),
    .X(_02814_));
 sky130_fd_sc_hd__inv_2 _23373_ (.A(_02814_),
    .Y(_02815_));
 sky130_fd_sc_hd__xnor2_1 _23374_ (.A(net125),
    .B(_02791_),
    .Y(_02816_));
 sky130_fd_sc_hd__o211ai_1 _23375_ (.A1(net120),
    .A2(_02799_),
    .B1(_02816_),
    .C1(_02785_),
    .Y(_02817_));
 sky130_fd_sc_hd__nand2_1 _23376_ (.A(_02815_),
    .B(_02817_),
    .Y(_02818_));
 sky130_fd_sc_hd__xnor2_1 _23377_ (.A(_02810_),
    .B(_02818_),
    .Y(_02819_));
 sky130_fd_sc_hd__o21ai_1 _23378_ (.A1(net1014),
    .A2(_02819_),
    .B1(net178),
    .Y(_02820_));
 sky130_fd_sc_hd__nor2_1 _23379_ (.A(net116),
    .B(_11857_),
    .Y(_02821_));
 sky130_fd_sc_hd__a22o_1 _23380_ (.A1(net116),
    .A2(_02820_),
    .B1(_02821_),
    .B2(_02819_),
    .X(_00517_));
 sky130_fd_sc_hd__a2bb2o_1 _23381_ (.A1_N(_11789_),
    .A2_N(_11629_),
    .B1(_02712_),
    .B2(_11560_),
    .X(_02822_));
 sky130_fd_sc_hd__a22o_1 _23382_ (.A1(net215),
    .A2(_11448_),
    .B1(_11730_),
    .B2(_02713_),
    .X(_02823_));
 sky130_fd_sc_hd__a21o_1 _23383_ (.A1(net187),
    .A2(_02822_),
    .B1(_02823_),
    .X(_02824_));
 sky130_fd_sc_hd__or3_1 _23384_ (.A(_02796_),
    .B(_02797_),
    .C(_02807_),
    .X(_02825_));
 sky130_fd_sc_hd__nand2_1 _23385_ (.A(_11513_),
    .B(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__xnor2_2 _23386_ (.A(_02824_),
    .B(_02826_),
    .Y(_02827_));
 sky130_fd_sc_hd__o21a_1 _23387_ (.A1(_02809_),
    .A2(_02818_),
    .B1(net116),
    .X(_02828_));
 sky130_fd_sc_hd__a21o_1 _23388_ (.A1(_02809_),
    .A2(_02818_),
    .B1(_02828_),
    .X(_02829_));
 sky130_fd_sc_hd__xnor2_1 _23389_ (.A(_02827_),
    .B(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__a21oi_1 _23390_ (.A1(_11650_),
    .A2(_02830_),
    .B1(net1020),
    .Y(_02831_));
 sky130_fd_sc_hd__or3_1 _23391_ (.A(net111),
    .B(_11784_),
    .C(_02830_),
    .X(_02832_));
 sky130_fd_sc_hd__o21ai_1 _23392_ (.A1(_01213_),
    .A2(_02831_),
    .B1(_02832_),
    .Y(_00518_));
 sky130_fd_sc_hd__o22a_1 _23393_ (.A1(_11632_),
    .A2(net216),
    .B1(_11715_),
    .B2(_02657_),
    .X(_02833_));
 sky130_fd_sc_hd__or2_1 _23394_ (.A(_11714_),
    .B(_02650_),
    .X(_02834_));
 sky130_fd_sc_hd__o221a_2 _23395_ (.A1(net215),
    .A2(_11560_),
    .B1(_02833_),
    .B2(_11654_),
    .C1(_02834_),
    .X(_02835_));
 sky130_fd_sc_hd__or2_1 _23396_ (.A(_02824_),
    .B(_02825_),
    .X(_02836_));
 sky130_fd_sc_hd__nand2_1 _23397_ (.A(_11513_),
    .B(_02836_),
    .Y(_02837_));
 sky130_fd_sc_hd__xor2_2 _23398_ (.A(_02835_),
    .B(_02837_),
    .X(_02838_));
 sky130_fd_sc_hd__nand2_1 _23399_ (.A(net112),
    .B(_02827_),
    .Y(_02839_));
 sky130_fd_sc_hd__o2111a_1 _23400_ (.A1(_01065_),
    .A2(_02810_),
    .B1(_02815_),
    .C1(_02817_),
    .D1(_02839_),
    .X(_02840_));
 sky130_fd_sc_hd__nor2_1 _23401_ (.A(net111),
    .B(_02827_),
    .Y(_02841_));
 sky130_fd_sc_hd__a311o_1 _23402_ (.A1(_01065_),
    .A2(_02810_),
    .A3(_02839_),
    .B1(_02840_),
    .C1(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__xor2_1 _23403_ (.A(_02838_),
    .B(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__o21ai_1 _23404_ (.A1(net1014),
    .A2(_02843_),
    .B1(net178),
    .Y(_02844_));
 sky130_fd_sc_hd__nor2_1 _23405_ (.A(net108),
    .B(_11857_),
    .Y(_02845_));
 sky130_fd_sc_hd__a22o_1 _23406_ (.A1(net107),
    .A2(_02844_),
    .B1(_02845_),
    .B2(_02843_),
    .X(_00519_));
 sky130_fd_sc_hd__or2_1 _23407_ (.A(_02835_),
    .B(_02836_),
    .X(_02846_));
 sky130_fd_sc_hd__nand2_1 _23408_ (.A(_11514_),
    .B(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__mux2_1 _23409_ (.A0(net216),
    .A1(_02663_),
    .S(_11730_),
    .X(_02848_));
 sky130_fd_sc_hd__xnor2_2 _23410_ (.A(_02847_),
    .B(_02848_),
    .Y(_02849_));
 sky130_fd_sc_hd__o21a_1 _23411_ (.A1(_02838_),
    .A2(_02842_),
    .B1(_01211_),
    .X(_02850_));
 sky130_fd_sc_hd__a21o_1 _23412_ (.A1(_02838_),
    .A2(_02842_),
    .B1(_02850_),
    .X(_02851_));
 sky130_fd_sc_hd__xnor2_1 _23413_ (.A(_02849_),
    .B(_02851_),
    .Y(_02852_));
 sky130_fd_sc_hd__o21ai_1 _23414_ (.A1(_11439_),
    .A2(_02852_),
    .B1(net176),
    .Y(_02853_));
 sky130_fd_sc_hd__nor2_1 _23415_ (.A(net103),
    .B(_11857_),
    .Y(_02854_));
 sky130_fd_sc_hd__a22o_1 _23416_ (.A1(net103),
    .A2(_02853_),
    .B1(_02854_),
    .B2(_02852_),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _23417_ (.A0(net215),
    .A1(_02687_),
    .S(_11730_),
    .X(_02855_));
 sky130_fd_sc_hd__or2_1 _23418_ (.A(_02846_),
    .B(_02848_),
    .X(_02856_));
 sky130_fd_sc_hd__nand2_1 _23419_ (.A(_11514_),
    .B(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__xnor2_2 _23420_ (.A(_02855_),
    .B(_02857_),
    .Y(_02858_));
 sky130_fd_sc_hd__nand2_1 _23421_ (.A(net103),
    .B(_02849_),
    .Y(_02859_));
 sky130_fd_sc_hd__nor2_1 _23422_ (.A(net103),
    .B(_02849_),
    .Y(_02860_));
 sky130_fd_sc_hd__a21o_1 _23423_ (.A1(_02851_),
    .A2(_02859_),
    .B1(_02860_),
    .X(_02861_));
 sky130_fd_sc_hd__xor2_1 _23424_ (.A(_02858_),
    .B(_02861_),
    .X(_02862_));
 sky130_fd_sc_hd__a21o_1 _23425_ (.A1(_11650_),
    .A2(_02862_),
    .B1(_11954_),
    .X(_02863_));
 sky130_fd_sc_hd__or3_1 _23426_ (.A(net98),
    .B(_11783_),
    .C(_02862_),
    .X(_02864_));
 sky130_fd_sc_hd__a21bo_1 _23427_ (.A1(net98),
    .A2(_02863_),
    .B1_N(_02864_),
    .X(_00521_));
 sky130_fd_sc_hd__a22o_1 _23428_ (.A1(net215),
    .A2(_11760_),
    .B1(_02712_),
    .B2(_11730_),
    .X(_02865_));
 sky130_fd_sc_hd__or2_1 _23429_ (.A(_02855_),
    .B(_02856_),
    .X(_02866_));
 sky130_fd_sc_hd__nand2_1 _23430_ (.A(_11515_),
    .B(_02866_),
    .Y(_02867_));
 sky130_fd_sc_hd__xnor2_2 _23431_ (.A(_02865_),
    .B(_02867_),
    .Y(_02868_));
 sky130_fd_sc_hd__a21bo_1 _23432_ (.A1(\top0.cordic0.vec[1][14] ),
    .A2(_02858_),
    .B1_N(_02861_),
    .X(_02869_));
 sky130_fd_sc_hd__or2_1 _23433_ (.A(\top0.cordic0.vec[1][14] ),
    .B(_02858_),
    .X(_02870_));
 sky130_fd_sc_hd__nand2_1 _23434_ (.A(_02869_),
    .B(_02870_),
    .Y(_02871_));
 sky130_fd_sc_hd__xor2_1 _23435_ (.A(_02868_),
    .B(_02871_),
    .X(_02872_));
 sky130_fd_sc_hd__a21o_1 _23436_ (.A1(_11649_),
    .A2(_02872_),
    .B1(_11954_),
    .X(_02873_));
 sky130_fd_sc_hd__nor2_1 _23437_ (.A(_11784_),
    .B(_02872_),
    .Y(_02874_));
 sky130_fd_sc_hd__mux2_1 _23438_ (.A0(_02873_),
    .A1(_02874_),
    .S(_01166_),
    .X(_02875_));
 sky130_fd_sc_hd__clkbuf_1 _23439_ (.A(_02875_),
    .X(_00522_));
 sky130_fd_sc_hd__o211a_1 _23440_ (.A1(net94),
    .A2(_02868_),
    .B1(_02869_),
    .C1(_02870_),
    .X(_02876_));
 sky130_fd_sc_hd__a21o_1 _23441_ (.A1(\top0.cordic0.vec[1][15] ),
    .A2(_02868_),
    .B1(_02876_),
    .X(_02877_));
 sky130_fd_sc_hd__mux2_2 _23442_ (.A0(_02657_),
    .A1(net217),
    .S(_11776_),
    .X(_02878_));
 sky130_fd_sc_hd__nor2_1 _23443_ (.A(_02865_),
    .B(_02866_),
    .Y(_02879_));
 sky130_fd_sc_hd__or2_1 _23444_ (.A(_11519_),
    .B(_02879_),
    .X(_02880_));
 sky130_fd_sc_hd__xnor2_1 _23445_ (.A(_02878_),
    .B(_02880_),
    .Y(_02881_));
 sky130_fd_sc_hd__xnor2_1 _23446_ (.A(_02877_),
    .B(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__a21o_1 _23447_ (.A1(_11650_),
    .A2(_02882_),
    .B1(_11954_),
    .X(_02883_));
 sky130_fd_sc_hd__or3_1 _23448_ (.A(net88),
    .B(_11783_),
    .C(_02882_),
    .X(_02884_));
 sky130_fd_sc_hd__a21bo_1 _23449_ (.A1(net88),
    .A2(_02883_),
    .B1_N(_02884_),
    .X(_00523_));
 sky130_fd_sc_hd__nor2_1 _23450_ (.A(_01230_),
    .B(_11519_),
    .Y(_02885_));
 sky130_fd_sc_hd__a21o_1 _23451_ (.A1(_02879_),
    .A2(_02878_),
    .B1(_02877_),
    .X(_02886_));
 sky130_fd_sc_hd__nor2_1 _23452_ (.A(net88),
    .B(_02878_),
    .Y(_02887_));
 sky130_fd_sc_hd__o21a_1 _23453_ (.A1(_02879_),
    .A2(_02877_),
    .B1(_02887_),
    .X(_02888_));
 sky130_fd_sc_hd__mux2_1 _23454_ (.A0(_11515_),
    .A1(_02878_),
    .S(net89),
    .X(_02889_));
 sky130_fd_sc_hd__nor2_1 _23455_ (.A(_02877_),
    .B(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__a211o_1 _23456_ (.A1(_02885_),
    .A2(_02886_),
    .B1(_02888_),
    .C1(_02890_),
    .X(_02891_));
 sky130_fd_sc_hd__xnor2_1 _23457_ (.A(_11789_),
    .B(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__nor3_1 _23458_ (.A(net85),
    .B(_11857_),
    .C(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__and3_1 _23459_ (.A(net85),
    .B(_11649_),
    .C(_02892_),
    .X(_02894_));
 sky130_fd_sc_hd__a211o_1 _23460_ (.A1(_11651_),
    .A2(net85),
    .B1(_02893_),
    .C1(_02894_),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _23461_ (.A0(\top0.cordic0.sin[0] ),
    .A1(\top0.matmul0.sin[0] ),
    .S(_05461_),
    .X(_02895_));
 sky130_fd_sc_hd__clkbuf_1 _23462_ (.A(_02895_),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _23463_ (.A0(net1003),
    .A1(\top0.matmul0.sin[1] ),
    .S(_05461_),
    .X(_02896_));
 sky130_fd_sc_hd__clkbuf_1 _23464_ (.A(_02896_),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _23465_ (.A0(\top0.cordic0.sin[2] ),
    .A1(\top0.matmul0.sin[2] ),
    .S(_05461_),
    .X(_02897_));
 sky130_fd_sc_hd__clkbuf_1 _23466_ (.A(_02897_),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _23467_ (.A0(net1010),
    .A1(\top0.matmul0.sin[3] ),
    .S(_05461_),
    .X(_02898_));
 sky130_fd_sc_hd__clkbuf_1 _23468_ (.A(_02898_),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _23469_ (.A0(net727),
    .A1(\top0.matmul0.sin[4] ),
    .S(_05461_),
    .X(_02899_));
 sky130_fd_sc_hd__clkbuf_1 _23470_ (.A(_02899_),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _23471_ (.A0(net920),
    .A1(\top0.matmul0.sin[5] ),
    .S(_05461_),
    .X(_02900_));
 sky130_fd_sc_hd__clkbuf_1 _23472_ (.A(_02900_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _23473_ (.A0(net1005),
    .A1(\top0.matmul0.sin[6] ),
    .S(_05461_),
    .X(_02901_));
 sky130_fd_sc_hd__clkbuf_1 _23474_ (.A(_02901_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _23475_ (.A0(net1000),
    .A1(\top0.matmul0.sin[7] ),
    .S(_05461_),
    .X(_02902_));
 sky130_fd_sc_hd__clkbuf_1 _23476_ (.A(_02902_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _23477_ (.A0(net1001),
    .A1(\top0.matmul0.sin[8] ),
    .S(_05461_),
    .X(_02903_));
 sky130_fd_sc_hd__clkbuf_1 _23478_ (.A(_02903_),
    .X(_00533_));
 sky130_fd_sc_hd__buf_4 _23479_ (.A(_05460_),
    .X(_02904_));
 sky130_fd_sc_hd__mux2_1 _23480_ (.A0(net999),
    .A1(\top0.matmul0.sin[9] ),
    .S(_02904_),
    .X(_02905_));
 sky130_fd_sc_hd__clkbuf_1 _23481_ (.A(_02905_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _23482_ (.A0(net928),
    .A1(\top0.matmul0.sin[10] ),
    .S(_02904_),
    .X(_02906_));
 sky130_fd_sc_hd__clkbuf_1 _23483_ (.A(_02906_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _23484_ (.A0(\top0.cordic0.sin[11] ),
    .A1(\top0.matmul0.sin[11] ),
    .S(_02904_),
    .X(_02907_));
 sky130_fd_sc_hd__clkbuf_1 _23485_ (.A(_02907_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _23486_ (.A0(net996),
    .A1(\top0.matmul0.sin[12] ),
    .S(_02904_),
    .X(_02908_));
 sky130_fd_sc_hd__clkbuf_1 _23487_ (.A(_02908_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _23488_ (.A0(net1007),
    .A1(\top0.matmul0.sin[13] ),
    .S(_02904_),
    .X(_02909_));
 sky130_fd_sc_hd__clkbuf_1 _23489_ (.A(_02909_),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _23490_ (.A0(net732),
    .A1(\top0.matmul0.cos[0] ),
    .S(_02904_),
    .X(_02910_));
 sky130_fd_sc_hd__clkbuf_1 _23491_ (.A(_02910_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _23492_ (.A0(\top0.cordic0.cos[1] ),
    .A1(\top0.matmul0.cos[1] ),
    .S(_02904_),
    .X(_02911_));
 sky130_fd_sc_hd__clkbuf_1 _23493_ (.A(_02911_),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_1 _23494_ (.A0(\top0.cordic0.cos[2] ),
    .A1(\top0.matmul0.cos[2] ),
    .S(_02904_),
    .X(_02912_));
 sky130_fd_sc_hd__clkbuf_1 _23495_ (.A(_02912_),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_1 _23496_ (.A0(net718),
    .A1(\top0.matmul0.cos[3] ),
    .S(_02904_),
    .X(_02913_));
 sky130_fd_sc_hd__clkbuf_1 _23497_ (.A(_02913_),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_1 _23498_ (.A0(net1002),
    .A1(\top0.matmul0.cos[4] ),
    .S(_02904_),
    .X(_02914_));
 sky130_fd_sc_hd__clkbuf_1 _23499_ (.A(_02914_),
    .X(_00543_));
 sky130_fd_sc_hd__clkbuf_4 _23500_ (.A(_05460_),
    .X(_02915_));
 sky130_fd_sc_hd__mux2_1 _23501_ (.A0(\top0.cordic0.cos[5] ),
    .A1(\top0.matmul0.cos[5] ),
    .S(_02915_),
    .X(_02916_));
 sky130_fd_sc_hd__clkbuf_1 _23502_ (.A(_02916_),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_1 _23503_ (.A0(net1008),
    .A1(\top0.matmul0.cos[6] ),
    .S(_02915_),
    .X(_02917_));
 sky130_fd_sc_hd__clkbuf_1 _23504_ (.A(_02917_),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _23505_ (.A0(\top0.cordic0.cos[7] ),
    .A1(\top0.matmul0.cos[7] ),
    .S(_02915_),
    .X(_02918_));
 sky130_fd_sc_hd__clkbuf_1 _23506_ (.A(_02918_),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _23507_ (.A0(net771),
    .A1(\top0.matmul0.cos[8] ),
    .S(_02915_),
    .X(_02919_));
 sky130_fd_sc_hd__clkbuf_1 _23508_ (.A(_02919_),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _23509_ (.A0(\top0.cordic0.cos[9] ),
    .A1(\top0.matmul0.cos[9] ),
    .S(_02915_),
    .X(_02920_));
 sky130_fd_sc_hd__clkbuf_1 _23510_ (.A(_02920_),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _23511_ (.A0(net794),
    .A1(\top0.matmul0.cos[10] ),
    .S(_02915_),
    .X(_02921_));
 sky130_fd_sc_hd__clkbuf_1 _23512_ (.A(_02921_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _23513_ (.A0(\top0.cordic0.cos[11] ),
    .A1(\top0.matmul0.cos[11] ),
    .S(_02915_),
    .X(_02922_));
 sky130_fd_sc_hd__clkbuf_1 _23514_ (.A(_02922_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _23515_ (.A0(\top0.cordic0.cos[12] ),
    .A1(\top0.matmul0.cos[12] ),
    .S(_02915_),
    .X(_02923_));
 sky130_fd_sc_hd__clkbuf_1 _23516_ (.A(_02923_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _23517_ (.A0(\top0.cordic0.cos[13] ),
    .A1(\top0.matmul0.cos[13] ),
    .S(_02915_),
    .X(_02924_));
 sky130_fd_sc_hd__clkbuf_1 _23518_ (.A(_02924_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _23519_ (.A0(\top0.a_in_matmul[0] ),
    .A1(\top0.matmul0.a[0] ),
    .S(_02915_),
    .X(_02925_));
 sky130_fd_sc_hd__clkbuf_1 _23520_ (.A(_02925_),
    .X(_00553_));
 sky130_fd_sc_hd__clkbuf_4 _23521_ (.A(_05460_),
    .X(_02926_));
 sky130_fd_sc_hd__mux2_1 _23522_ (.A0(\top0.a_in_matmul[1] ),
    .A1(\top0.matmul0.a[1] ),
    .S(_02926_),
    .X(_02927_));
 sky130_fd_sc_hd__clkbuf_1 _23523_ (.A(_02927_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _23524_ (.A0(net979),
    .A1(\top0.matmul0.a[2] ),
    .S(_02926_),
    .X(_02928_));
 sky130_fd_sc_hd__clkbuf_1 _23525_ (.A(_02928_),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _23526_ (.A0(\top0.a_in_matmul[3] ),
    .A1(\top0.matmul0.a[3] ),
    .S(_02926_),
    .X(_02929_));
 sky130_fd_sc_hd__clkbuf_1 _23527_ (.A(_02929_),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _23528_ (.A0(\top0.a_in_matmul[4] ),
    .A1(\top0.matmul0.a[4] ),
    .S(_02926_),
    .X(_02930_));
 sky130_fd_sc_hd__clkbuf_1 _23529_ (.A(_02930_),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _23530_ (.A0(\top0.a_in_matmul[5] ),
    .A1(\top0.matmul0.a[5] ),
    .S(_02926_),
    .X(_02931_));
 sky130_fd_sc_hd__clkbuf_1 _23531_ (.A(_02931_),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _23532_ (.A0(\top0.a_in_matmul[6] ),
    .A1(\top0.matmul0.a[6] ),
    .S(_02926_),
    .X(_02932_));
 sky130_fd_sc_hd__clkbuf_1 _23533_ (.A(_02932_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _23534_ (.A0(\top0.a_in_matmul[7] ),
    .A1(\top0.matmul0.a[7] ),
    .S(_02926_),
    .X(_02933_));
 sky130_fd_sc_hd__clkbuf_1 _23535_ (.A(_02933_),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _23536_ (.A0(net985),
    .A1(\top0.matmul0.a[8] ),
    .S(_02926_),
    .X(_02934_));
 sky130_fd_sc_hd__clkbuf_1 _23537_ (.A(_02934_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _23538_ (.A0(\top0.a_in_matmul[9] ),
    .A1(\top0.matmul0.a[9] ),
    .S(_02926_),
    .X(_02935_));
 sky130_fd_sc_hd__clkbuf_1 _23539_ (.A(_02935_),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _23540_ (.A0(\top0.a_in_matmul[10] ),
    .A1(\top0.matmul0.a[10] ),
    .S(_02926_),
    .X(_02936_));
 sky130_fd_sc_hd__clkbuf_1 _23541_ (.A(_02936_),
    .X(_00563_));
 sky130_fd_sc_hd__clkbuf_4 _23542_ (.A(_05460_),
    .X(_02937_));
 sky130_fd_sc_hd__mux2_1 _23543_ (.A0(\top0.a_in_matmul[11] ),
    .A1(\top0.matmul0.a[11] ),
    .S(_02937_),
    .X(_02938_));
 sky130_fd_sc_hd__clkbuf_1 _23544_ (.A(_02938_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _23545_ (.A0(\top0.a_in_matmul[12] ),
    .A1(\top0.matmul0.a[12] ),
    .S(_02937_),
    .X(_02939_));
 sky130_fd_sc_hd__clkbuf_1 _23546_ (.A(_02939_),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _23547_ (.A0(\top0.a_in_matmul[13] ),
    .A1(\top0.matmul0.a[13] ),
    .S(_02937_),
    .X(_02940_));
 sky130_fd_sc_hd__clkbuf_1 _23548_ (.A(_02940_),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _23549_ (.A0(\top0.a_in_matmul[14] ),
    .A1(\top0.matmul0.a[14] ),
    .S(_02937_),
    .X(_02941_));
 sky130_fd_sc_hd__clkbuf_1 _23550_ (.A(_02941_),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _23551_ (.A0(\top0.a_in_matmul[15] ),
    .A1(\top0.matmul0.a[15] ),
    .S(_02937_),
    .X(_02942_));
 sky130_fd_sc_hd__clkbuf_1 _23552_ (.A(_02942_),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _23553_ (.A0(\top0.b_in_matmul[0] ),
    .A1(\top0.matmul0.b[0] ),
    .S(_02937_),
    .X(_02943_));
 sky130_fd_sc_hd__clkbuf_1 _23554_ (.A(_02943_),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _23555_ (.A0(\top0.b_in_matmul[1] ),
    .A1(\top0.matmul0.b[1] ),
    .S(_02937_),
    .X(_02944_));
 sky130_fd_sc_hd__clkbuf_1 _23556_ (.A(_02944_),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _23557_ (.A0(\top0.b_in_matmul[2] ),
    .A1(\top0.matmul0.b[2] ),
    .S(_02937_),
    .X(_02945_));
 sky130_fd_sc_hd__clkbuf_1 _23558_ (.A(_02945_),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _23559_ (.A0(\top0.b_in_matmul[3] ),
    .A1(\top0.matmul0.b[3] ),
    .S(_02937_),
    .X(_02946_));
 sky130_fd_sc_hd__clkbuf_1 _23560_ (.A(_02946_),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_1 _23561_ (.A0(\top0.b_in_matmul[4] ),
    .A1(\top0.matmul0.b[4] ),
    .S(_02937_),
    .X(_02947_));
 sky130_fd_sc_hd__clkbuf_1 _23562_ (.A(_02947_),
    .X(_00573_));
 sky130_fd_sc_hd__clkbuf_4 _23563_ (.A(_05460_),
    .X(_02948_));
 sky130_fd_sc_hd__mux2_1 _23564_ (.A0(net965),
    .A1(\top0.matmul0.b[5] ),
    .S(_02948_),
    .X(_02949_));
 sky130_fd_sc_hd__clkbuf_1 _23565_ (.A(_02949_),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _23566_ (.A0(net966),
    .A1(\top0.matmul0.b[6] ),
    .S(_02948_),
    .X(_02950_));
 sky130_fd_sc_hd__clkbuf_1 _23567_ (.A(_02950_),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _23568_ (.A0(\top0.b_in_matmul[7] ),
    .A1(\top0.matmul0.b[7] ),
    .S(_02948_),
    .X(_02951_));
 sky130_fd_sc_hd__clkbuf_1 _23569_ (.A(_02951_),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _23570_ (.A0(\top0.b_in_matmul[8] ),
    .A1(\top0.matmul0.b[8] ),
    .S(_02948_),
    .X(_02952_));
 sky130_fd_sc_hd__clkbuf_1 _23571_ (.A(_02952_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _23572_ (.A0(\top0.b_in_matmul[9] ),
    .A1(\top0.matmul0.b[9] ),
    .S(_02948_),
    .X(_02953_));
 sky130_fd_sc_hd__clkbuf_1 _23573_ (.A(_02953_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _23574_ (.A0(\top0.b_in_matmul[10] ),
    .A1(\top0.matmul0.b[10] ),
    .S(_02948_),
    .X(_02954_));
 sky130_fd_sc_hd__clkbuf_1 _23575_ (.A(_02954_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _23576_ (.A0(net980),
    .A1(\top0.matmul0.b[11] ),
    .S(_02948_),
    .X(_02955_));
 sky130_fd_sc_hd__clkbuf_1 _23577_ (.A(_02955_),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _23578_ (.A0(\top0.b_in_matmul[12] ),
    .A1(\top0.matmul0.b[12] ),
    .S(_02948_),
    .X(_02956_));
 sky130_fd_sc_hd__clkbuf_1 _23579_ (.A(_02956_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _23580_ (.A0(\top0.b_in_matmul[13] ),
    .A1(\top0.matmul0.b[13] ),
    .S(_02948_),
    .X(_02957_));
 sky130_fd_sc_hd__clkbuf_1 _23581_ (.A(_02957_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _23582_ (.A0(net1009),
    .A1(\top0.matmul0.b[14] ),
    .S(_02948_),
    .X(_02958_));
 sky130_fd_sc_hd__clkbuf_1 _23583_ (.A(_02958_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _23584_ (.A0(\top0.b_in_matmul[15] ),
    .A1(net943),
    .S(_05460_),
    .X(_02959_));
 sky130_fd_sc_hd__clkbuf_1 _23585_ (.A(_02959_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _23586_ (.A0(\top0.matmul0.alpha_pass[0] ),
    .A1(_09251_),
    .S(net560),
    .X(_02960_));
 sky130_fd_sc_hd__clkbuf_1 _23587_ (.A(_02960_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _23588_ (.A0(\top0.matmul0.alpha_pass[1] ),
    .A1(_09255_),
    .S(net560),
    .X(_02961_));
 sky130_fd_sc_hd__clkbuf_1 _23589_ (.A(_02961_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _23590_ (.A0(\top0.matmul0.alpha_pass[2] ),
    .A1(_09261_),
    .S(net559),
    .X(_02962_));
 sky130_fd_sc_hd__clkbuf_1 _23591_ (.A(_02962_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _23592_ (.A0(\top0.matmul0.alpha_pass[3] ),
    .A1(_09267_),
    .S(net559),
    .X(_02963_));
 sky130_fd_sc_hd__clkbuf_1 _23593_ (.A(_02963_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _23594_ (.A0(\top0.matmul0.alpha_pass[4] ),
    .A1(_09272_),
    .S(net559),
    .X(_02964_));
 sky130_fd_sc_hd__clkbuf_1 _23595_ (.A(_02964_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _23596_ (.A0(net76),
    .A1(_09278_),
    .S(net559),
    .X(_02965_));
 sky130_fd_sc_hd__clkbuf_1 _23597_ (.A(_02965_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _23598_ (.A0(\top0.matmul0.alpha_pass[6] ),
    .A1(_09284_),
    .S(net559),
    .X(_02966_));
 sky130_fd_sc_hd__clkbuf_1 _23599_ (.A(_02966_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _23600_ (.A0(\top0.matmul0.alpha_pass[7] ),
    .A1(_09290_),
    .S(net561),
    .X(_02967_));
 sky130_fd_sc_hd__clkbuf_1 _23601_ (.A(_02967_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _23602_ (.A0(net1024),
    .A1(_09296_),
    .S(net559),
    .X(_02968_));
 sky130_fd_sc_hd__clkbuf_1 _23603_ (.A(_02968_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _23604_ (.A0(\top0.matmul0.alpha_pass[9] ),
    .A1(_09302_),
    .S(net559),
    .X(_02969_));
 sky130_fd_sc_hd__clkbuf_1 _23605_ (.A(_02969_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _23606_ (.A0(\top0.matmul0.alpha_pass[10] ),
    .A1(_09308_),
    .S(net559),
    .X(_02970_));
 sky130_fd_sc_hd__clkbuf_1 _23607_ (.A(_02970_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _23608_ (.A0(\top0.matmul0.alpha_pass[11] ),
    .A1(_09314_),
    .S(net559),
    .X(_02971_));
 sky130_fd_sc_hd__clkbuf_1 _23609_ (.A(_02971_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _23610_ (.A0(\top0.matmul0.alpha_pass[12] ),
    .A1(_09320_),
    .S(net559),
    .X(_02972_));
 sky130_fd_sc_hd__clkbuf_1 _23611_ (.A(_02972_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _23612_ (.A0(\top0.matmul0.alpha_pass[13] ),
    .A1(_09325_),
    .S(net560),
    .X(_02973_));
 sky130_fd_sc_hd__clkbuf_1 _23613_ (.A(_02973_),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _23614_ (.A0(\top0.matmul0.alpha_pass[14] ),
    .A1(_09331_),
    .S(net561),
    .X(_02974_));
 sky130_fd_sc_hd__clkbuf_1 _23615_ (.A(_02974_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _23616_ (.A0(\top0.matmul0.alpha_pass[15] ),
    .A1(_09337_),
    .S(net561),
    .X(_02975_));
 sky130_fd_sc_hd__clkbuf_1 _23617_ (.A(_02975_),
    .X(_00600_));
 sky130_fd_sc_hd__o21a_4 _23618_ (.A1(net569),
    .A2(net572),
    .B1(\top0.matmul0.matmul_stage_inst.f[4] ),
    .X(_02976_));
 sky130_fd_sc_hd__o21a_4 _23619_ (.A1(net564),
    .A2(net557),
    .B1(\top0.matmul0.matmul_stage_inst.e[4] ),
    .X(_02977_));
 sky130_fd_sc_hd__nor2_2 _23620_ (.A(_02976_),
    .B(_02977_),
    .Y(_02978_));
 sky130_fd_sc_hd__a22o_2 _23621_ (.A1(net574),
    .A2(\top0.matmul0.matmul_stage_inst.d[8] ),
    .B1(\top0.matmul0.matmul_stage_inst.c[8] ),
    .B2(net558),
    .X(_02979_));
 sky130_fd_sc_hd__a22o_4 _23622_ (.A1(net570),
    .A2(\top0.matmul0.matmul_stage_inst.b[8] ),
    .B1(\top0.matmul0.matmul_stage_inst.a[8] ),
    .B2(net567),
    .X(_02980_));
 sky130_fd_sc_hd__nor2_1 _23623_ (.A(_02979_),
    .B(_02980_),
    .Y(_02981_));
 sky130_fd_sc_hd__buf_4 _23624_ (.A(_02981_),
    .X(_02982_));
 sky130_fd_sc_hd__nor2_2 _23625_ (.A(_02978_),
    .B(_02982_),
    .Y(_02983_));
 sky130_fd_sc_hd__o21a_1 _23626_ (.A1(net569),
    .A2(net572),
    .B1(\top0.matmul0.matmul_stage_inst.f[5] ),
    .X(_02984_));
 sky130_fd_sc_hd__clkbuf_4 _23627_ (.A(_02984_),
    .X(_02985_));
 sky130_fd_sc_hd__o21a_1 _23628_ (.A1(net565),
    .A2(net557),
    .B1(\top0.matmul0.matmul_stage_inst.e[5] ),
    .X(_02986_));
 sky130_fd_sc_hd__clkbuf_4 _23629_ (.A(_02986_),
    .X(_02987_));
 sky130_fd_sc_hd__a22o_1 _23630_ (.A1(net574),
    .A2(\top0.matmul0.matmul_stage_inst.d[7] ),
    .B1(\top0.matmul0.matmul_stage_inst.c[7] ),
    .B2(net558),
    .X(_02988_));
 sky130_fd_sc_hd__clkbuf_4 _23631_ (.A(_02988_),
    .X(_02989_));
 sky130_fd_sc_hd__a22o_1 _23632_ (.A1(net570),
    .A2(\top0.matmul0.matmul_stage_inst.b[7] ),
    .B1(\top0.matmul0.matmul_stage_inst.a[7] ),
    .B2(net566),
    .X(_02990_));
 sky130_fd_sc_hd__clkbuf_4 _23633_ (.A(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__o22a_1 _23634_ (.A1(_02985_),
    .A2(_02987_),
    .B1(_02989_),
    .B2(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__o21a_1 _23635_ (.A1(net568),
    .A2(net573),
    .B1(\top0.matmul0.matmul_stage_inst.f[6] ),
    .X(_02993_));
 sky130_fd_sc_hd__buf_2 _23636_ (.A(_02993_),
    .X(_02994_));
 sky130_fd_sc_hd__o21a_1 _23637_ (.A1(net565),
    .A2(net557),
    .B1(\top0.matmul0.matmul_stage_inst.e[6] ),
    .X(_02995_));
 sky130_fd_sc_hd__clkbuf_4 _23638_ (.A(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__a22o_1 _23639_ (.A1(net569),
    .A2(\top0.matmul0.matmul_stage_inst.b[6] ),
    .B1(\top0.matmul0.matmul_stage_inst.a[6] ),
    .B2(net564),
    .X(_02997_));
 sky130_fd_sc_hd__clkbuf_4 _23640_ (.A(_02997_),
    .X(_02998_));
 sky130_fd_sc_hd__a22o_1 _23641_ (.A1(net572),
    .A2(\top0.matmul0.matmul_stage_inst.d[6] ),
    .B1(\top0.matmul0.matmul_stage_inst.c[6] ),
    .B2(net558),
    .X(_02999_));
 sky130_fd_sc_hd__clkbuf_4 _23642_ (.A(_02999_),
    .X(_03000_));
 sky130_fd_sc_hd__o22a_1 _23643_ (.A1(_02994_),
    .A2(_02996_),
    .B1(_02998_),
    .B2(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__xor2_2 _23644_ (.A(_02992_),
    .B(_03001_),
    .X(_03002_));
 sky130_fd_sc_hd__xnor2_4 _23645_ (.A(_02983_),
    .B(_03002_),
    .Y(_03003_));
 sky130_fd_sc_hd__a22o_4 _23646_ (.A1(net570),
    .A2(\top0.matmul0.matmul_stage_inst.b[5] ),
    .B1(\top0.matmul0.matmul_stage_inst.a[5] ),
    .B2(net566),
    .X(_03004_));
 sky130_fd_sc_hd__a22o_4 _23647_ (.A1(net574),
    .A2(\top0.matmul0.matmul_stage_inst.d[5] ),
    .B1(\top0.matmul0.matmul_stage_inst.c[5] ),
    .B2(net558),
    .X(_03005_));
 sky130_fd_sc_hd__nor2_4 _23648_ (.A(_03004_),
    .B(_03005_),
    .Y(_03006_));
 sky130_fd_sc_hd__nor2_2 _23649_ (.A(_02993_),
    .B(_02995_),
    .Y(_03007_));
 sky130_fd_sc_hd__nor2_2 _23650_ (.A(_03006_),
    .B(_03007_),
    .Y(_03008_));
 sky130_fd_sc_hd__o22a_2 _23651_ (.A1(_02976_),
    .A2(_02977_),
    .B1(_02988_),
    .B2(_02990_),
    .X(_03009_));
 sky130_fd_sc_hd__or2_2 _23652_ (.A(_03004_),
    .B(_03005_),
    .X(_03010_));
 sky130_fd_sc_hd__or2_1 _23653_ (.A(_02993_),
    .B(_02995_),
    .X(_03011_));
 sky130_fd_sc_hd__o22a_1 _23654_ (.A1(_02984_),
    .A2(_02986_),
    .B1(_02997_),
    .B2(_02999_),
    .X(_03012_));
 sky130_fd_sc_hd__a31o_1 _23655_ (.A1(_03010_),
    .A2(_03011_),
    .A3(_03009_),
    .B1(_03012_),
    .X(_03013_));
 sky130_fd_sc_hd__o21ai_2 _23656_ (.A1(_03008_),
    .A2(_03009_),
    .B1(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__o21a_4 _23657_ (.A1(net569),
    .A2(net573),
    .B1(\top0.matmul0.matmul_stage_inst.f[2] ),
    .X(_03015_));
 sky130_fd_sc_hd__o21a_4 _23658_ (.A1(net565),
    .A2(net557),
    .B1(\top0.matmul0.matmul_stage_inst.e[2] ),
    .X(_03016_));
 sky130_fd_sc_hd__nor2_4 _23659_ (.A(_03015_),
    .B(_03016_),
    .Y(_03017_));
 sky130_fd_sc_hd__a22o_2 _23660_ (.A1(net572),
    .A2(\top0.matmul0.matmul_stage_inst.d[10] ),
    .B1(\top0.matmul0.matmul_stage_inst.c[10] ),
    .B2(net557),
    .X(_03018_));
 sky130_fd_sc_hd__a22o_2 _23661_ (.A1(net569),
    .A2(\top0.matmul0.matmul_stage_inst.b[10] ),
    .B1(\top0.matmul0.matmul_stage_inst.a[10] ),
    .B2(net564),
    .X(_03019_));
 sky130_fd_sc_hd__nor2_1 _23662_ (.A(_03018_),
    .B(_03019_),
    .Y(_03020_));
 sky130_fd_sc_hd__nor2_1 _23663_ (.A(_03017_),
    .B(net1017),
    .Y(_03021_));
 sky130_fd_sc_hd__o21a_1 _23664_ (.A1(net569),
    .A2(net573),
    .B1(\top0.matmul0.matmul_stage_inst.f[3] ),
    .X(_03022_));
 sky130_fd_sc_hd__o21a_1 _23665_ (.A1(net565),
    .A2(net557),
    .B1(\top0.matmul0.matmul_stage_inst.e[3] ),
    .X(_03023_));
 sky130_fd_sc_hd__a22o_4 _23666_ (.A1(net574),
    .A2(\top0.matmul0.matmul_stage_inst.d[9] ),
    .B1(\top0.matmul0.matmul_stage_inst.c[9] ),
    .B2(net558),
    .X(_03024_));
 sky130_fd_sc_hd__a22o_4 _23667_ (.A1(net570),
    .A2(\top0.matmul0.matmul_stage_inst.b[9] ),
    .B1(\top0.matmul0.matmul_stage_inst.a[9] ),
    .B2(net566),
    .X(_03025_));
 sky130_fd_sc_hd__o22a_1 _23668_ (.A1(_03022_),
    .A2(_03023_),
    .B1(_03024_),
    .B2(_03025_),
    .X(_03026_));
 sky130_fd_sc_hd__o21a_4 _23669_ (.A1(net569),
    .A2(net573),
    .B1(\top0.matmul0.matmul_stage_inst.f[1] ),
    .X(_03027_));
 sky130_fd_sc_hd__o21a_4 _23670_ (.A1(net565),
    .A2(net557),
    .B1(\top0.matmul0.matmul_stage_inst.e[1] ),
    .X(_03028_));
 sky130_fd_sc_hd__a22o_4 _23671_ (.A1(net568),
    .A2(\top0.matmul0.matmul_stage_inst.b[11] ),
    .B1(\top0.matmul0.matmul_stage_inst.a[11] ),
    .B2(net564),
    .X(_03029_));
 sky130_fd_sc_hd__a22o_4 _23672_ (.A1(net572),
    .A2(\top0.matmul0.matmul_stage_inst.d[11] ),
    .B1(\top0.matmul0.matmul_stage_inst.c[11] ),
    .B2(net556),
    .X(_03030_));
 sky130_fd_sc_hd__o22a_1 _23673_ (.A1(_03027_),
    .A2(_03028_),
    .B1(_03029_),
    .B2(_03030_),
    .X(_03031_));
 sky130_fd_sc_hd__xor2_1 _23674_ (.A(_03026_),
    .B(_03031_),
    .X(_03032_));
 sky130_fd_sc_hd__xnor2_2 _23675_ (.A(_03021_),
    .B(_03032_),
    .Y(_03033_));
 sky130_fd_sc_hd__xnor2_2 _23676_ (.A(_03014_),
    .B(_03033_),
    .Y(_03034_));
 sky130_fd_sc_hd__xnor2_4 _23677_ (.A(_03003_),
    .B(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__a22o_2 _23678_ (.A1(net568),
    .A2(\top0.matmul0.matmul_stage_inst.b[4] ),
    .B1(\top0.matmul0.matmul_stage_inst.a[4] ),
    .B2(net564),
    .X(_03036_));
 sky130_fd_sc_hd__a22o_2 _23679_ (.A1(net572),
    .A2(\top0.matmul0.matmul_stage_inst.d[4] ),
    .B1(\top0.matmul0.matmul_stage_inst.c[4] ),
    .B2(net556),
    .X(_03037_));
 sky130_fd_sc_hd__o22a_1 _23680_ (.A1(_03036_),
    .A2(_03037_),
    .B1(_02993_),
    .B2(_02995_),
    .X(_03038_));
 sky130_fd_sc_hd__o22a_1 _23681_ (.A1(_02997_),
    .A2(_02999_),
    .B1(_02976_),
    .B2(_02977_),
    .X(_03039_));
 sky130_fd_sc_hd__or2_1 _23682_ (.A(_02984_),
    .B(_02986_),
    .X(_03040_));
 sky130_fd_sc_hd__a22o_1 _23683_ (.A1(_03010_),
    .A2(_03040_),
    .B1(_03038_),
    .B2(_03039_),
    .X(_03041_));
 sky130_fd_sc_hd__o21a_2 _23684_ (.A1(_03038_),
    .A2(_03039_),
    .B1(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__xnor2_2 _23685_ (.A(_03012_),
    .B(_03009_),
    .Y(_03043_));
 sky130_fd_sc_hd__xnor2_4 _23686_ (.A(_03008_),
    .B(_03043_),
    .Y(_03044_));
 sky130_fd_sc_hd__clkbuf_4 _23687_ (.A(_03022_),
    .X(_03045_));
 sky130_fd_sc_hd__clkbuf_4 _23688_ (.A(_03023_),
    .X(_03046_));
 sky130_fd_sc_hd__nor2_2 _23689_ (.A(_03045_),
    .B(_03046_),
    .Y(_03047_));
 sky130_fd_sc_hd__nor2_2 _23690_ (.A(_03047_),
    .B(_02982_),
    .Y(_03048_));
 sky130_fd_sc_hd__o22a_2 _23691_ (.A1(_03024_),
    .A2(_03025_),
    .B1(_03015_),
    .B2(_03016_),
    .X(_03049_));
 sky130_fd_sc_hd__o22a_2 _23692_ (.A1(_03018_),
    .A2(_03019_),
    .B1(_03027_),
    .B2(_03028_),
    .X(_03050_));
 sky130_fd_sc_hd__xnor2_2 _23693_ (.A(_03049_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__xnor2_4 _23694_ (.A(_03048_),
    .B(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__o21a_1 _23695_ (.A1(_03042_),
    .A2(_03044_),
    .B1(_03052_),
    .X(_03053_));
 sky130_fd_sc_hd__o21a_4 _23696_ (.A1(net571),
    .A2(net574),
    .B1(\top0.matmul0.matmul_stage_inst.f[7] ),
    .X(_03054_));
 sky130_fd_sc_hd__o21a_4 _23697_ (.A1(net566),
    .A2(net560),
    .B1(\top0.matmul0.matmul_stage_inst.e[7] ),
    .X(_03055_));
 sky130_fd_sc_hd__or2_2 _23698_ (.A(_03054_),
    .B(_03055_),
    .X(_03056_));
 sky130_fd_sc_hd__o21a_2 _23699_ (.A1(net574),
    .A2(net566),
    .B1(\top0.matmul0.matmul_stage_inst.a[3] ),
    .X(_03057_));
 sky130_fd_sc_hd__a22o_2 _23700_ (.A1(net556),
    .A2(\top0.matmul0.matmul_stage_inst.c[3] ),
    .B1(\top0.matmul0.matmul_stage_inst.b[3] ),
    .B2(net568),
    .X(_03058_));
 sky130_fd_sc_hd__or2_1 _23701_ (.A(_03057_),
    .B(_03058_),
    .X(_03059_));
 sky130_fd_sc_hd__clkbuf_4 _23702_ (.A(_03059_),
    .X(_03060_));
 sky130_fd_sc_hd__o21a_4 _23703_ (.A1(net570),
    .A2(net575),
    .B1(\top0.matmul0.matmul_stage_inst.f[9] ),
    .X(_03061_));
 sky130_fd_sc_hd__o21a_4 _23704_ (.A1(net567),
    .A2(net560),
    .B1(\top0.matmul0.matmul_stage_inst.e[9] ),
    .X(_03062_));
 sky130_fd_sc_hd__a22o_4 _23705_ (.A1(net568),
    .A2(\top0.matmul0.matmul_stage_inst.b[1] ),
    .B1(\top0.matmul0.matmul_stage_inst.a[1] ),
    .B2(net564),
    .X(_03063_));
 sky130_fd_sc_hd__a22o_4 _23706_ (.A1(net572),
    .A2(\top0.matmul0.matmul_stage_inst.d[1] ),
    .B1(\top0.matmul0.matmul_stage_inst.c[1] ),
    .B2(net556),
    .X(_03064_));
 sky130_fd_sc_hd__o22a_2 _23707_ (.A1(_03061_),
    .A2(_03062_),
    .B1(_03063_),
    .B2(_03064_),
    .X(_03065_));
 sky130_fd_sc_hd__a22o_2 _23708_ (.A1(net568),
    .A2(\top0.matmul0.matmul_stage_inst.b[2] ),
    .B1(\top0.matmul0.matmul_stage_inst.a[2] ),
    .B2(net564),
    .X(_03066_));
 sky130_fd_sc_hd__a22o_2 _23709_ (.A1(net572),
    .A2(\top0.matmul0.matmul_stage_inst.d[2] ),
    .B1(\top0.matmul0.matmul_stage_inst.c[2] ),
    .B2(net556),
    .X(_03067_));
 sky130_fd_sc_hd__o21a_1 _23710_ (.A1(net571),
    .A2(net574),
    .B1(\top0.matmul0.matmul_stage_inst.f[8] ),
    .X(_03068_));
 sky130_fd_sc_hd__clkbuf_4 _23711_ (.A(_03068_),
    .X(_03069_));
 sky130_fd_sc_hd__o21a_1 _23712_ (.A1(net567),
    .A2(net558),
    .B1(\top0.matmul0.matmul_stage_inst.e[8] ),
    .X(_03070_));
 sky130_fd_sc_hd__clkbuf_4 _23713_ (.A(_03070_),
    .X(_03071_));
 sky130_fd_sc_hd__o22a_1 _23714_ (.A1(_03066_),
    .A2(_03067_),
    .B1(_03069_),
    .B2(_03071_),
    .X(_03072_));
 sky130_fd_sc_hd__a22o_1 _23715_ (.A1(_03056_),
    .A2(_03060_),
    .B1(_03065_),
    .B2(_03072_),
    .X(_03073_));
 sky130_fd_sc_hd__or2_1 _23716_ (.A(_03065_),
    .B(_03072_),
    .X(_03074_));
 sky130_fd_sc_hd__and2_2 _23717_ (.A(_03073_),
    .B(_03074_),
    .X(_03075_));
 sky130_fd_sc_hd__clkbuf_4 _23718_ (.A(_03066_),
    .X(_03076_));
 sky130_fd_sc_hd__clkbuf_4 _23719_ (.A(_03067_),
    .X(_03077_));
 sky130_fd_sc_hd__o22a_4 _23720_ (.A1(_03061_),
    .A2(_03062_),
    .B1(_03076_),
    .B2(_03077_),
    .X(_03078_));
 sky130_fd_sc_hd__o22a_1 _23721_ (.A1(_03036_),
    .A2(_03037_),
    .B1(_03054_),
    .B2(_03055_),
    .X(_03079_));
 sky130_fd_sc_hd__o22a_1 _23722_ (.A1(_03069_),
    .A2(_03071_),
    .B1(_03057_),
    .B2(_03058_),
    .X(_03080_));
 sky130_fd_sc_hd__xnor2_2 _23723_ (.A(_03079_),
    .B(_03080_),
    .Y(_03081_));
 sky130_fd_sc_hd__xnor2_4 _23724_ (.A(_03078_),
    .B(_03081_),
    .Y(_03082_));
 sky130_fd_sc_hd__a22o_1 _23725_ (.A1(_03042_),
    .A2(_03044_),
    .B1(_03075_),
    .B2(_03082_),
    .X(_03083_));
 sky130_fd_sc_hd__o211ai_1 _23726_ (.A1(_03042_),
    .A2(_03052_),
    .B1(_03075_),
    .C1(_03082_),
    .Y(_03084_));
 sky130_fd_sc_hd__a21oi_1 _23727_ (.A1(_03042_),
    .A2(_03052_),
    .B1(_03044_),
    .Y(_03085_));
 sky130_fd_sc_hd__o22a_2 _23728_ (.A1(_03053_),
    .A2(_03083_),
    .B1(_03084_),
    .B2(_03085_),
    .X(_03086_));
 sky130_fd_sc_hd__xor2_4 _23729_ (.A(_03035_),
    .B(_03086_),
    .X(_03087_));
 sky130_fd_sc_hd__a22o_2 _23730_ (.A1(net574),
    .A2(\top0.matmul0.matmul_stage_inst.d[0] ),
    .B1(\top0.matmul0.matmul_stage_inst.a[0] ),
    .B2(net566),
    .X(_03088_));
 sky130_fd_sc_hd__o21a_2 _23731_ (.A1(net569),
    .A2(net556),
    .B1(\top0.matmul0.matmul_stage_inst.b[0] ),
    .X(_03089_));
 sky130_fd_sc_hd__o21a_4 _23732_ (.A1(net570),
    .A2(net574),
    .B1(\top0.matmul0.matmul_stage_inst.f[11] ),
    .X(_03090_));
 sky130_fd_sc_hd__o21a_4 _23733_ (.A1(net567),
    .A2(net558),
    .B1(\top0.matmul0.matmul_stage_inst.e[11] ),
    .X(_03091_));
 sky130_fd_sc_hd__o22a_2 _23734_ (.A1(_03088_),
    .A2(_03089_),
    .B1(_03090_),
    .B2(_03091_),
    .X(_03092_));
 sky130_fd_sc_hd__o21a_2 _23735_ (.A1(net570),
    .A2(net575),
    .B1(\top0.matmul0.matmul_stage_inst.f[10] ),
    .X(_03093_));
 sky130_fd_sc_hd__o21a_2 _23736_ (.A1(net567),
    .A2(net560),
    .B1(\top0.matmul0.matmul_stage_inst.e[10] ),
    .X(_03094_));
 sky130_fd_sc_hd__o22a_2 _23737_ (.A1(_03063_),
    .A2(_03064_),
    .B1(_03093_),
    .B2(_03094_),
    .X(_03095_));
 sky130_fd_sc_hd__xor2_1 _23738_ (.A(_03092_),
    .B(_03095_),
    .X(_03096_));
 sky130_fd_sc_hd__nand3_1 _23739_ (.A(_03073_),
    .B(_03074_),
    .C(_03096_),
    .Y(_03097_));
 sky130_fd_sc_hd__xnor2_4 _23740_ (.A(_03092_),
    .B(_03095_),
    .Y(_03098_));
 sky130_fd_sc_hd__a21o_1 _23741_ (.A1(_03073_),
    .A2(_03074_),
    .B1(_03098_),
    .X(_03099_));
 sky130_fd_sc_hd__mux2_2 _23742_ (.A0(_03097_),
    .A1(_03099_),
    .S(_03082_),
    .X(_03100_));
 sky130_fd_sc_hd__nand2_1 _23743_ (.A(_03087_),
    .B(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__o22a_2 _23744_ (.A1(_03063_),
    .A2(_03064_),
    .B1(_03090_),
    .B2(_03091_),
    .X(_03102_));
 sky130_fd_sc_hd__o21a_2 _23745_ (.A1(net571),
    .A2(net575),
    .B1(\top0.matmul0.matmul_stage_inst.f[12] ),
    .X(_03103_));
 sky130_fd_sc_hd__o21a_2 _23746_ (.A1(net566),
    .A2(net558),
    .B1(\top0.matmul0.matmul_stage_inst.e[12] ),
    .X(_03104_));
 sky130_fd_sc_hd__o22a_2 _23747_ (.A1(_03088_),
    .A2(_03089_),
    .B1(_03103_),
    .B2(_03104_),
    .X(_03105_));
 sky130_fd_sc_hd__nor2_4 _23748_ (.A(_03066_),
    .B(_03067_),
    .Y(_03106_));
 sky130_fd_sc_hd__nor2_1 _23749_ (.A(_03093_),
    .B(_03094_),
    .Y(_03107_));
 sky130_fd_sc_hd__nor2_1 _23750_ (.A(_03106_),
    .B(_03107_),
    .Y(_03108_));
 sky130_fd_sc_hd__xnor2_2 _23751_ (.A(_03105_),
    .B(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__xnor2_4 _23752_ (.A(_03102_),
    .B(_03109_),
    .Y(_03110_));
 sky130_fd_sc_hd__o21bai_1 _23753_ (.A1(_03087_),
    .A2(_03100_),
    .B1_N(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__nor2_4 _23754_ (.A(_03061_),
    .B(_03062_),
    .Y(_03112_));
 sky130_fd_sc_hd__nor2_1 _23755_ (.A(_03057_),
    .B(_03058_),
    .Y(_03113_));
 sky130_fd_sc_hd__buf_4 _23756_ (.A(_03113_),
    .X(_03114_));
 sky130_fd_sc_hd__nor2_2 _23757_ (.A(_03112_),
    .B(_03114_),
    .Y(_03115_));
 sky130_fd_sc_hd__o22a_1 _23758_ (.A1(_03036_),
    .A2(_03037_),
    .B1(_03069_),
    .B2(_03071_),
    .X(_03116_));
 sky130_fd_sc_hd__o22a_1 _23759_ (.A1(_03004_),
    .A2(_03005_),
    .B1(_03054_),
    .B2(_03055_),
    .X(_03117_));
 sky130_fd_sc_hd__xnor2_2 _23760_ (.A(_03116_),
    .B(_03117_),
    .Y(_03118_));
 sky130_fd_sc_hd__xnor2_4 _23761_ (.A(_03115_),
    .B(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__or2_4 _23762_ (.A(_03088_),
    .B(_03089_),
    .X(_03120_));
 sky130_fd_sc_hd__or2_1 _23763_ (.A(_03063_),
    .B(_03064_),
    .X(_03121_));
 sky130_fd_sc_hd__or2_1 _23764_ (.A(_03090_),
    .B(_03091_),
    .X(_03122_));
 sky130_fd_sc_hd__buf_6 _23765_ (.A(_03122_),
    .X(_03123_));
 sky130_fd_sc_hd__or2_2 _23766_ (.A(_03093_),
    .B(_03094_),
    .X(_03124_));
 sky130_fd_sc_hd__and4_2 _23767_ (.A(_03120_),
    .B(_03121_),
    .C(_03123_),
    .D(_03124_),
    .X(_03125_));
 sky130_fd_sc_hd__and2_1 _23768_ (.A(_03078_),
    .B(_03079_),
    .X(_03126_));
 sky130_fd_sc_hd__o21a_1 _23769_ (.A1(_03078_),
    .A2(_03079_),
    .B1(_03080_),
    .X(_03127_));
 sky130_fd_sc_hd__nor2_1 _23770_ (.A(_03126_),
    .B(_03127_),
    .Y(_03128_));
 sky130_fd_sc_hd__xnor2_2 _23771_ (.A(_03125_),
    .B(_03128_),
    .Y(_03129_));
 sky130_fd_sc_hd__xor2_4 _23772_ (.A(_03119_),
    .B(_03129_),
    .X(_03130_));
 sky130_fd_sc_hd__a21oi_2 _23773_ (.A1(_03101_),
    .A2(_03111_),
    .B1(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__nor2_1 _23774_ (.A(_03087_),
    .B(_03100_),
    .Y(_03132_));
 sky130_fd_sc_hd__and2_1 _23775_ (.A(_03110_),
    .B(_03130_),
    .X(_03133_));
 sky130_fd_sc_hd__xnor2_4 _23776_ (.A(_03075_),
    .B(_03082_),
    .Y(_03134_));
 sky130_fd_sc_hd__nor2_1 _23777_ (.A(_03098_),
    .B(_03134_),
    .Y(_03135_));
 sky130_fd_sc_hd__nor2_1 _23778_ (.A(_03110_),
    .B(_03135_),
    .Y(_03136_));
 sky130_fd_sc_hd__a22o_1 _23779_ (.A1(_03132_),
    .A2(_03133_),
    .B1(_03136_),
    .B2(_03087_),
    .X(_03137_));
 sky130_fd_sc_hd__nand2_1 _23780_ (.A(_03075_),
    .B(_03082_),
    .Y(_03138_));
 sky130_fd_sc_hd__or2_1 _23781_ (.A(_03035_),
    .B(_03138_),
    .X(_03139_));
 sky130_fd_sc_hd__nor2_1 _23782_ (.A(_03042_),
    .B(_03052_),
    .Y(_03140_));
 sky130_fd_sc_hd__a211o_1 _23783_ (.A1(_03035_),
    .A2(_03138_),
    .B1(_03140_),
    .C1(_03085_),
    .X(_03141_));
 sky130_fd_sc_hd__nor2_1 _23784_ (.A(_03049_),
    .B(_03050_),
    .Y(_03142_));
 sky130_fd_sc_hd__nand2_1 _23785_ (.A(_03049_),
    .B(_03050_),
    .Y(_03143_));
 sky130_fd_sc_hd__o31ai_2 _23786_ (.A1(_03047_),
    .A2(_02982_),
    .A3(_03142_),
    .B1(_03143_),
    .Y(_03144_));
 sky130_fd_sc_hd__or2_1 _23787_ (.A(net571),
    .B(net575),
    .X(_03145_));
 sky130_fd_sc_hd__buf_4 _23788_ (.A(_03145_),
    .X(_03146_));
 sky130_fd_sc_hd__or2_1 _23789_ (.A(net567),
    .B(net560),
    .X(_03147_));
 sky130_fd_sc_hd__buf_4 _23790_ (.A(_03147_),
    .X(_03148_));
 sky130_fd_sc_hd__a22oi_4 _23791_ (.A1(\top0.matmul0.matmul_stage_inst.f[0] ),
    .A2(_03146_),
    .B1(_03148_),
    .B2(\top0.matmul0.matmul_stage_inst.e[0] ),
    .Y(_03149_));
 sky130_fd_sc_hd__a22o_2 _23792_ (.A1(net568),
    .A2(\top0.matmul0.matmul_stage_inst.b[12] ),
    .B1(\top0.matmul0.matmul_stage_inst.a[12] ),
    .B2(net564),
    .X(_03150_));
 sky130_fd_sc_hd__a22o_2 _23793_ (.A1(net572),
    .A2(\top0.matmul0.matmul_stage_inst.d[12] ),
    .B1(\top0.matmul0.matmul_stage_inst.c[12] ),
    .B2(net556),
    .X(_03151_));
 sky130_fd_sc_hd__nor2_2 _23794_ (.A(_03150_),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__nor2_1 _23795_ (.A(_03149_),
    .B(_03152_),
    .Y(_03153_));
 sky130_fd_sc_hd__and2_1 _23796_ (.A(_03144_),
    .B(_03153_),
    .X(_03154_));
 sky130_fd_sc_hd__o21ai_2 _23797_ (.A1(net569),
    .A2(net573),
    .B1(\top0.matmul0.matmul_stage_inst.f[2] ),
    .Y(_03155_));
 sky130_fd_sc_hd__o21ai_2 _23798_ (.A1(net565),
    .A2(net557),
    .B1(\top0.matmul0.matmul_stage_inst.e[2] ),
    .Y(_03156_));
 sky130_fd_sc_hd__nand2_2 _23799_ (.A(_03155_),
    .B(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__or2_2 _23800_ (.A(_03018_),
    .B(_03019_),
    .X(_03158_));
 sky130_fd_sc_hd__a31o_1 _23801_ (.A1(_03157_),
    .A2(_03158_),
    .A3(_03031_),
    .B1(_03026_),
    .X(_03159_));
 sky130_fd_sc_hd__o21a_2 _23802_ (.A1(_03021_),
    .A2(_03031_),
    .B1(_03159_),
    .X(_03160_));
 sky130_fd_sc_hd__buf_4 _23803_ (.A(_03149_),
    .X(_03161_));
 sky130_fd_sc_hd__a22o_2 _23804_ (.A1(net572),
    .A2(\top0.matmul0.matmul_stage_inst.d[13] ),
    .B1(\top0.matmul0.matmul_stage_inst.c[13] ),
    .B2(net556),
    .X(_03162_));
 sky130_fd_sc_hd__a22o_2 _23805_ (.A1(net568),
    .A2(\top0.matmul0.matmul_stage_inst.b[13] ),
    .B1(\top0.matmul0.matmul_stage_inst.a[13] ),
    .B2(net564),
    .X(_03163_));
 sky130_fd_sc_hd__nor2_1 _23806_ (.A(_03162_),
    .B(_03163_),
    .Y(_03164_));
 sky130_fd_sc_hd__nor2_2 _23807_ (.A(_03161_),
    .B(_03164_),
    .Y(_03165_));
 sky130_fd_sc_hd__xnor2_4 _23808_ (.A(_03160_),
    .B(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__xor2_1 _23809_ (.A(_03154_),
    .B(_03166_),
    .X(_03167_));
 sky130_fd_sc_hd__and3_1 _23810_ (.A(_03139_),
    .B(_03141_),
    .C(_03167_),
    .X(_03168_));
 sky130_fd_sc_hd__a21oi_2 _23811_ (.A1(_03139_),
    .A2(_03141_),
    .B1(_03167_),
    .Y(_03169_));
 sky130_fd_sc_hd__or2_1 _23812_ (.A(_03014_),
    .B(_03033_),
    .X(_03170_));
 sky130_fd_sc_hd__a21o_1 _23813_ (.A1(_03014_),
    .A2(_03033_),
    .B1(_03003_),
    .X(_03171_));
 sky130_fd_sc_hd__or3_1 _23814_ (.A(_03125_),
    .B(_03126_),
    .C(_03127_),
    .X(_03172_));
 sky130_fd_sc_hd__o21a_1 _23815_ (.A1(_03126_),
    .A2(_03127_),
    .B1(_03125_),
    .X(_03173_));
 sky130_fd_sc_hd__a21o_1 _23816_ (.A1(_03119_),
    .A2(_03172_),
    .B1(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__a21o_1 _23817_ (.A1(_03170_),
    .A2(_03171_),
    .B1(_03174_),
    .X(_03175_));
 sky130_fd_sc_hd__nand3_1 _23818_ (.A(_03174_),
    .B(_03170_),
    .C(_03171_),
    .Y(_03176_));
 sky130_fd_sc_hd__o22a_2 _23819_ (.A1(_02976_),
    .A2(_02977_),
    .B1(_03024_),
    .B2(_03025_),
    .X(_03177_));
 sky130_fd_sc_hd__o22a_1 _23820_ (.A1(_02985_),
    .A2(_02987_),
    .B1(_02979_),
    .B2(_02980_),
    .X(_03178_));
 sky130_fd_sc_hd__o22a_1 _23821_ (.A1(_02994_),
    .A2(_02996_),
    .B1(_02989_),
    .B2(_02991_),
    .X(_03179_));
 sky130_fd_sc_hd__xnor2_1 _23822_ (.A(_03178_),
    .B(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__xnor2_2 _23823_ (.A(_03177_),
    .B(_03180_),
    .Y(_03181_));
 sky130_fd_sc_hd__and2_1 _23824_ (.A(_02992_),
    .B(_03001_),
    .X(_03182_));
 sky130_fd_sc_hd__nor2_1 _23825_ (.A(_02992_),
    .B(_03001_),
    .Y(_03183_));
 sky130_fd_sc_hd__o21ba_1 _23826_ (.A1(_02983_),
    .A2(_03182_),
    .B1_N(_03183_),
    .X(_03184_));
 sky130_fd_sc_hd__nor2_4 _23827_ (.A(_03027_),
    .B(_03028_),
    .Y(_03185_));
 sky130_fd_sc_hd__nor2_2 _23828_ (.A(_03185_),
    .B(_03152_),
    .Y(_03186_));
 sky130_fd_sc_hd__o22a_1 _23829_ (.A1(_03015_),
    .A2(_03016_),
    .B1(_03029_),
    .B2(_03030_),
    .X(_03187_));
 sky130_fd_sc_hd__o22a_1 _23830_ (.A1(_03045_),
    .A2(_03046_),
    .B1(_03018_),
    .B2(_03019_),
    .X(_03188_));
 sky130_fd_sc_hd__xnor2_1 _23831_ (.A(_03187_),
    .B(_03188_),
    .Y(_03189_));
 sky130_fd_sc_hd__xnor2_2 _23832_ (.A(_03186_),
    .B(_03189_),
    .Y(_03190_));
 sky130_fd_sc_hd__xnor2_1 _23833_ (.A(_03184_),
    .B(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__xnor2_2 _23834_ (.A(_03181_),
    .B(_03191_),
    .Y(_03192_));
 sky130_fd_sc_hd__a21o_1 _23835_ (.A1(_03175_),
    .A2(_03176_),
    .B1(_03192_),
    .X(_03193_));
 sky130_fd_sc_hd__nand3_2 _23836_ (.A(_03192_),
    .B(_03175_),
    .C(_03176_),
    .Y(_03194_));
 sky130_fd_sc_hd__nor2_4 _23837_ (.A(_03088_),
    .B(_03089_),
    .Y(_03195_));
 sky130_fd_sc_hd__o21a_2 _23838_ (.A1(net570),
    .A2(net575),
    .B1(\top0.matmul0.matmul_stage_inst.f[13] ),
    .X(_03196_));
 sky130_fd_sc_hd__o21a_2 _23839_ (.A1(net566),
    .A2(net560),
    .B1(\top0.matmul0.matmul_stage_inst.e[13] ),
    .X(_03197_));
 sky130_fd_sc_hd__nor2_2 _23840_ (.A(_03196_),
    .B(_03197_),
    .Y(_03198_));
 sky130_fd_sc_hd__nor2_2 _23841_ (.A(_03195_),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__buf_4 _23842_ (.A(_03107_),
    .X(_03200_));
 sky130_fd_sc_hd__nor2_1 _23843_ (.A(_03114_),
    .B(_03200_),
    .Y(_03201_));
 sky130_fd_sc_hd__o22a_1 _23844_ (.A1(_03063_),
    .A2(_03064_),
    .B1(_03103_),
    .B2(_03104_),
    .X(_03202_));
 sky130_fd_sc_hd__o22a_1 _23845_ (.A1(_03076_),
    .A2(_03077_),
    .B1(_03090_),
    .B2(_03091_),
    .X(_03203_));
 sky130_fd_sc_hd__xnor2_1 _23846_ (.A(_03202_),
    .B(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__xnor2_2 _23847_ (.A(_03201_),
    .B(_03204_),
    .Y(_03205_));
 sky130_fd_sc_hd__xor2_2 _23848_ (.A(_03199_),
    .B(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__clkbuf_4 _23849_ (.A(_03036_),
    .X(_03207_));
 sky130_fd_sc_hd__clkbuf_4 _23850_ (.A(_03037_),
    .X(_03208_));
 sky130_fd_sc_hd__o22a_1 _23851_ (.A1(_03207_),
    .A2(_03208_),
    .B1(_03061_),
    .B2(_03062_),
    .X(_03209_));
 sky130_fd_sc_hd__o22a_1 _23852_ (.A1(_02998_),
    .A2(_03000_),
    .B1(_03054_),
    .B2(_03055_),
    .X(_03210_));
 sky130_fd_sc_hd__o22a_1 _23853_ (.A1(_03004_),
    .A2(_03005_),
    .B1(_03069_),
    .B2(_03071_),
    .X(_03211_));
 sky130_fd_sc_hd__xor2_1 _23854_ (.A(_03210_),
    .B(_03211_),
    .X(_03212_));
 sky130_fd_sc_hd__xnor2_2 _23855_ (.A(_03209_),
    .B(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hd__o2bb2a_1 _23856_ (.A1_N(_03116_),
    .A2_N(_03117_),
    .B1(_03112_),
    .B2(_03113_),
    .X(_03214_));
 sky130_fd_sc_hd__nor2_1 _23857_ (.A(_03116_),
    .B(_03117_),
    .Y(_03215_));
 sky130_fd_sc_hd__or2_1 _23858_ (.A(_03076_),
    .B(_03077_),
    .X(_03216_));
 sky130_fd_sc_hd__clkbuf_4 _23859_ (.A(_03216_),
    .X(_03217_));
 sky130_fd_sc_hd__o211ai_1 _23860_ (.A1(_03102_),
    .A2(_03105_),
    .B1(_03124_),
    .C1(_03217_),
    .Y(_03218_));
 sky130_fd_sc_hd__nand2_1 _23861_ (.A(_03102_),
    .B(_03105_),
    .Y(_03219_));
 sky130_fd_sc_hd__o211a_1 _23862_ (.A1(_03214_),
    .A2(_03215_),
    .B1(_03218_),
    .C1(_03219_),
    .X(_03220_));
 sky130_fd_sc_hd__a211o_1 _23863_ (.A1(_03218_),
    .A2(_03219_),
    .B1(_03214_),
    .C1(_03215_),
    .X(_03221_));
 sky130_fd_sc_hd__and2b_1 _23864_ (.A_N(_03220_),
    .B(_03221_),
    .X(_03222_));
 sky130_fd_sc_hd__xnor2_2 _23865_ (.A(_03213_),
    .B(_03222_),
    .Y(_03223_));
 sky130_fd_sc_hd__xnor2_2 _23866_ (.A(_03206_),
    .B(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__a21o_2 _23867_ (.A1(_03193_),
    .A2(_03194_),
    .B1(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__nand3_4 _23868_ (.A(_03193_),
    .B(_03194_),
    .C(_03224_),
    .Y(_03226_));
 sky130_fd_sc_hd__o211ai_4 _23869_ (.A1(_03168_),
    .A2(_03169_),
    .B1(_03225_),
    .C1(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__a211o_1 _23870_ (.A1(_03225_),
    .A2(_03226_),
    .B1(_03168_),
    .C1(_03169_),
    .X(_03228_));
 sky130_fd_sc_hd__o211ai_4 _23871_ (.A1(_03131_),
    .A2(_03137_),
    .B1(_03227_),
    .C1(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__a211o_1 _23872_ (.A1(_03227_),
    .A2(_03228_),
    .B1(_03131_),
    .C1(_03137_),
    .X(_03230_));
 sky130_fd_sc_hd__xnor2_4 _23873_ (.A(_03098_),
    .B(_03134_),
    .Y(_03231_));
 sky130_fd_sc_hd__xor2_2 _23874_ (.A(_03042_),
    .B(_03052_),
    .X(_03232_));
 sky130_fd_sc_hd__xnor2_4 _23875_ (.A(_03044_),
    .B(_03232_),
    .Y(_03233_));
 sky130_fd_sc_hd__nor2_2 _23876_ (.A(_02984_),
    .B(_02986_),
    .Y(_03234_));
 sky130_fd_sc_hd__nor2_2 _23877_ (.A(_03006_),
    .B(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__xnor2_2 _23878_ (.A(_03038_),
    .B(_03039_),
    .Y(_03236_));
 sky130_fd_sc_hd__xnor2_4 _23879_ (.A(_03235_),
    .B(_03236_),
    .Y(_03237_));
 sky130_fd_sc_hd__nor2_2 _23880_ (.A(_02981_),
    .B(_03017_),
    .Y(_03238_));
 sky130_fd_sc_hd__o22a_1 _23881_ (.A1(_03024_),
    .A2(_03025_),
    .B1(_03027_),
    .B2(_03028_),
    .X(_03239_));
 sky130_fd_sc_hd__o22a_1 _23882_ (.A1(_03022_),
    .A2(_03023_),
    .B1(_02988_),
    .B2(_02990_),
    .X(_03240_));
 sky130_fd_sc_hd__xnor2_2 _23883_ (.A(_03239_),
    .B(_03240_),
    .Y(_03241_));
 sky130_fd_sc_hd__xnor2_4 _23884_ (.A(_03238_),
    .B(_03241_),
    .Y(_03242_));
 sky130_fd_sc_hd__o22a_1 _23885_ (.A1(_03004_),
    .A2(_03005_),
    .B1(_02976_),
    .B2(_02977_),
    .X(_03243_));
 sky130_fd_sc_hd__o22a_1 _23886_ (.A1(_02984_),
    .A2(_02986_),
    .B1(_03207_),
    .B2(_03208_),
    .X(_03244_));
 sky130_fd_sc_hd__a22o_1 _23887_ (.A1(_03011_),
    .A2(_03060_),
    .B1(_03243_),
    .B2(_03244_),
    .X(_03245_));
 sky130_fd_sc_hd__o21a_1 _23888_ (.A1(_03243_),
    .A2(_03244_),
    .B1(_03245_),
    .X(_03246_));
 sky130_fd_sc_hd__a21oi_1 _23889_ (.A1(_03237_),
    .A2(_03242_),
    .B1(_03246_),
    .Y(_03247_));
 sky130_fd_sc_hd__or2_2 _23890_ (.A(_03061_),
    .B(_03062_),
    .X(_03248_));
 sky130_fd_sc_hd__nand2_1 _23891_ (.A(_03248_),
    .B(_03120_),
    .Y(_03249_));
 sky130_fd_sc_hd__nor2_2 _23892_ (.A(_03054_),
    .B(_03055_),
    .Y(_03250_));
 sky130_fd_sc_hd__nor2_1 _23893_ (.A(_03068_),
    .B(_03070_),
    .Y(_03251_));
 sky130_fd_sc_hd__nor2_4 _23894_ (.A(_03063_),
    .B(_03064_),
    .Y(_03252_));
 sky130_fd_sc_hd__or4_2 _23895_ (.A(_03250_),
    .B(_03106_),
    .C(_03251_),
    .D(_03252_),
    .X(_03253_));
 sky130_fd_sc_hd__clkbuf_4 _23896_ (.A(_03251_),
    .X(_03254_));
 sky130_fd_sc_hd__o22a_1 _23897_ (.A1(_03250_),
    .A2(_03106_),
    .B1(_03254_),
    .B2(_03252_),
    .X(_03255_));
 sky130_fd_sc_hd__a21oi_2 _23898_ (.A1(_03249_),
    .A2(_03253_),
    .B1(_03255_),
    .Y(_03256_));
 sky130_fd_sc_hd__nor2_2 _23899_ (.A(_03250_),
    .B(_03113_),
    .Y(_03257_));
 sky130_fd_sc_hd__xnor2_2 _23900_ (.A(_03065_),
    .B(_03072_),
    .Y(_03258_));
 sky130_fd_sc_hd__xnor2_1 _23901_ (.A(_03257_),
    .B(_03258_),
    .Y(_03259_));
 sky130_fd_sc_hd__a2bb2o_1 _23902_ (.A1_N(_03237_),
    .A2_N(_03242_),
    .B1(_03256_),
    .B2(_03259_),
    .X(_03260_));
 sky130_fd_sc_hd__a21o_1 _23903_ (.A1(_03249_),
    .A2(_03253_),
    .B1(_03255_),
    .X(_03261_));
 sky130_fd_sc_hd__xor2_2 _23904_ (.A(_03257_),
    .B(_03258_),
    .X(_03262_));
 sky130_fd_sc_hd__a211o_1 _23905_ (.A1(_03237_),
    .A2(_03242_),
    .B1(_03261_),
    .C1(_03262_),
    .X(_03263_));
 sky130_fd_sc_hd__o21a_1 _23906_ (.A1(_03237_),
    .A2(_03242_),
    .B1(_03246_),
    .X(_03264_));
 sky130_fd_sc_hd__o22a_2 _23907_ (.A1(_03247_),
    .A2(_03260_),
    .B1(_03263_),
    .B2(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__xnor2_4 _23908_ (.A(_03233_),
    .B(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__xnor2_2 _23909_ (.A(_03256_),
    .B(_03262_),
    .Y(_03267_));
 sky130_fd_sc_hd__nor2_1 _23910_ (.A(_03195_),
    .B(_03200_),
    .Y(_03268_));
 sky130_fd_sc_hd__nand2_2 _23911_ (.A(_03267_),
    .B(_03268_),
    .Y(_03269_));
 sky130_fd_sc_hd__a21oi_1 _23912_ (.A1(_03231_),
    .A2(_03266_),
    .B1(_03269_),
    .Y(_03270_));
 sky130_fd_sc_hd__nor2_1 _23913_ (.A(_03231_),
    .B(_03266_),
    .Y(_03271_));
 sky130_fd_sc_hd__nand2_1 _23914_ (.A(_03256_),
    .B(_03259_),
    .Y(_03272_));
 sky130_fd_sc_hd__nand2_1 _23915_ (.A(_03237_),
    .B(_03242_),
    .Y(_03273_));
 sky130_fd_sc_hd__o21ai_1 _23916_ (.A1(_03237_),
    .A2(_03242_),
    .B1(_03246_),
    .Y(_03274_));
 sky130_fd_sc_hd__a21o_1 _23917_ (.A1(_03273_),
    .A2(_03274_),
    .B1(_03272_),
    .X(_03275_));
 sky130_fd_sc_hd__a32o_2 _23918_ (.A1(_03272_),
    .A2(_03273_),
    .A3(_03274_),
    .B1(_03275_),
    .B2(_03233_),
    .X(_03276_));
 sky130_fd_sc_hd__and2_1 _23919_ (.A(_03239_),
    .B(_03240_),
    .X(_03277_));
 sky130_fd_sc_hd__nor2_1 _23920_ (.A(_03239_),
    .B(_03240_),
    .Y(_03278_));
 sky130_fd_sc_hd__o21ba_1 _23921_ (.A1(_03238_),
    .A2(_03277_),
    .B1_N(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__nor2_4 _23922_ (.A(_03029_),
    .B(_03030_),
    .Y(_03280_));
 sky130_fd_sc_hd__nor2_1 _23923_ (.A(_03280_),
    .B(_03149_),
    .Y(_03281_));
 sky130_fd_sc_hd__nand2_1 _23924_ (.A(_03279_),
    .B(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__xnor2_1 _23925_ (.A(_03144_),
    .B(_03153_),
    .Y(_03283_));
 sky130_fd_sc_hd__and2_1 _23926_ (.A(_03282_),
    .B(_03283_),
    .X(_03284_));
 sky130_fd_sc_hd__or2_1 _23927_ (.A(_03282_),
    .B(_03283_),
    .X(_03285_));
 sky130_fd_sc_hd__and2b_1 _23928_ (.A_N(_03284_),
    .B(_03285_),
    .X(_03286_));
 sky130_fd_sc_hd__xnor2_4 _23929_ (.A(_03276_),
    .B(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__xnor2_1 _23930_ (.A(_03110_),
    .B(_03100_),
    .Y(_03288_));
 sky130_fd_sc_hd__xor2_2 _23931_ (.A(_03130_),
    .B(_03288_),
    .X(_03289_));
 sky130_fd_sc_hd__xnor2_4 _23932_ (.A(_03087_),
    .B(_03289_),
    .Y(_03290_));
 sky130_fd_sc_hd__o21a_1 _23933_ (.A1(_03276_),
    .A2(_03284_),
    .B1(_03285_),
    .X(_03291_));
 sky130_fd_sc_hd__o311a_1 _23934_ (.A1(_03270_),
    .A2(_03271_),
    .A3(_03287_),
    .B1(_03290_),
    .C1(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__o21ai_2 _23935_ (.A1(_03269_),
    .A2(_03266_),
    .B1(_03231_),
    .Y(_03293_));
 sky130_fd_sc_hd__nand2_1 _23936_ (.A(_03269_),
    .B(_03266_),
    .Y(_03294_));
 sky130_fd_sc_hd__and4_1 _23937_ (.A(_03291_),
    .B(_03293_),
    .C(_03294_),
    .D(_03287_),
    .X(_03295_));
 sky130_fd_sc_hd__or4_1 _23938_ (.A(_03291_),
    .B(_03270_),
    .C(_03271_),
    .D(_03287_),
    .X(_03296_));
 sky130_fd_sc_hd__a311o_1 _23939_ (.A1(_03293_),
    .A2(_03294_),
    .A3(_03287_),
    .B1(_03290_),
    .C1(_03291_),
    .X(_03297_));
 sky130_fd_sc_hd__and4bb_1 _23940_ (.A_N(_03292_),
    .B_N(_03295_),
    .C(_03296_),
    .D(_03297_),
    .X(_03298_));
 sky130_fd_sc_hd__a21oi_2 _23941_ (.A1(_03229_),
    .A2(_03230_),
    .B1(_03298_),
    .Y(_03299_));
 sky130_fd_sc_hd__and3_1 _23942_ (.A(_03229_),
    .B(_03230_),
    .C(_03298_),
    .X(_03300_));
 sky130_fd_sc_hd__nor2_2 _23943_ (.A(_03299_),
    .B(_03300_),
    .Y(_03301_));
 sky130_fd_sc_hd__nor2_2 _23944_ (.A(_03234_),
    .B(_03114_),
    .Y(_03302_));
 sky130_fd_sc_hd__o22a_1 _23945_ (.A1(_03207_),
    .A2(_03208_),
    .B1(_02976_),
    .B2(_02977_),
    .X(_03303_));
 sky130_fd_sc_hd__or2_1 _23946_ (.A(_03207_),
    .B(_03208_),
    .X(_03304_));
 sky130_fd_sc_hd__o22a_2 _23947_ (.A1(_02985_),
    .A2(_02987_),
    .B1(_02976_),
    .B2(_02977_),
    .X(_03305_));
 sky130_fd_sc_hd__o22a_1 _23948_ (.A1(_02994_),
    .A2(_02996_),
    .B1(_03076_),
    .B2(_03077_),
    .X(_03306_));
 sky130_fd_sc_hd__a31o_1 _23949_ (.A1(_03304_),
    .A2(_03305_),
    .A3(_03060_),
    .B1(_03306_),
    .X(_03307_));
 sky130_fd_sc_hd__o21a_2 _23950_ (.A1(_03302_),
    .A2(_03303_),
    .B1(_03307_),
    .X(_03308_));
 sky130_fd_sc_hd__nor2_2 _23951_ (.A(_03007_),
    .B(_03114_),
    .Y(_03309_));
 sky130_fd_sc_hd__xnor2_2 _23952_ (.A(_03243_),
    .B(_03244_),
    .Y(_03310_));
 sky130_fd_sc_hd__xnor2_4 _23953_ (.A(_03309_),
    .B(_03310_),
    .Y(_03311_));
 sky130_fd_sc_hd__nand2_1 _23954_ (.A(_03308_),
    .B(_03311_),
    .Y(_03312_));
 sky130_fd_sc_hd__or2_2 _23955_ (.A(_02998_),
    .B(_03000_),
    .X(_03313_));
 sky130_fd_sc_hd__or2_1 _23956_ (.A(_03045_),
    .B(_03046_),
    .X(_03314_));
 sky130_fd_sc_hd__clkbuf_4 _23957_ (.A(_03314_),
    .X(_03315_));
 sky130_fd_sc_hd__nand2_2 _23958_ (.A(_03313_),
    .B(_03315_),
    .Y(_03316_));
 sky130_fd_sc_hd__o22a_2 _23959_ (.A1(_03015_),
    .A2(_03016_),
    .B1(_02989_),
    .B2(_02991_),
    .X(_03317_));
 sky130_fd_sc_hd__o22a_1 _23960_ (.A1(_02979_),
    .A2(_02980_),
    .B1(_03027_),
    .B2(_03028_),
    .X(_03318_));
 sky130_fd_sc_hd__xnor2_2 _23961_ (.A(_03317_),
    .B(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__xnor2_4 _23962_ (.A(_03316_),
    .B(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__o21bai_2 _23963_ (.A1(_03308_),
    .A2(_03311_),
    .B1_N(_03320_),
    .Y(_03321_));
 sky130_fd_sc_hd__nor2_1 _23964_ (.A(_03248_),
    .B(_03217_),
    .Y(_03322_));
 sky130_fd_sc_hd__clkbuf_4 _23965_ (.A(_03120_),
    .X(_03323_));
 sky130_fd_sc_hd__clkbuf_4 _23966_ (.A(_03121_),
    .X(_03324_));
 sky130_fd_sc_hd__buf_4 _23967_ (.A(_03250_),
    .X(_03325_));
 sky130_fd_sc_hd__nor2_2 _23968_ (.A(_03325_),
    .B(_03254_),
    .Y(_03326_));
 sky130_fd_sc_hd__o2111ai_4 _23969_ (.A1(_03078_),
    .A2(_03322_),
    .B1(_03323_),
    .C1(_03324_),
    .D1(_03326_),
    .Y(_03327_));
 sky130_fd_sc_hd__a21o_1 _23970_ (.A1(_03312_),
    .A2(_03321_),
    .B1(_03327_),
    .X(_03328_));
 sky130_fd_sc_hd__nand3_2 _23971_ (.A(_03312_),
    .B(_03321_),
    .C(_03327_),
    .Y(_03329_));
 sky130_fd_sc_hd__nand2_1 _23972_ (.A(_03328_),
    .B(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__xnor2_1 _23973_ (.A(_03237_),
    .B(_03246_),
    .Y(_03331_));
 sky130_fd_sc_hd__xnor2_2 _23974_ (.A(_03242_),
    .B(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__xnor2_1 _23975_ (.A(_03267_),
    .B(_03268_),
    .Y(_03333_));
 sky130_fd_sc_hd__xor2_1 _23976_ (.A(_03332_),
    .B(_03333_),
    .X(_03334_));
 sky130_fd_sc_hd__xnor2_2 _23977_ (.A(_03330_),
    .B(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__o22a_1 _23978_ (.A1(_03004_),
    .A2(_03005_),
    .B1(_03022_),
    .B2(_03023_),
    .X(_03336_));
 sky130_fd_sc_hd__or2_2 _23979_ (.A(_03027_),
    .B(_03028_),
    .X(_03337_));
 sky130_fd_sc_hd__or2_1 _23980_ (.A(_02989_),
    .B(_02991_),
    .X(_03338_));
 sky130_fd_sc_hd__o22a_1 _23981_ (.A1(_02998_),
    .A2(_03000_),
    .B1(_03015_),
    .B2(_03016_),
    .X(_03339_));
 sky130_fd_sc_hd__a21o_1 _23982_ (.A1(_03337_),
    .A2(_03338_),
    .B1(_03339_),
    .X(_03340_));
 sky130_fd_sc_hd__and3_1 _23983_ (.A(_03337_),
    .B(_03338_),
    .C(_03339_),
    .X(_03341_));
 sky130_fd_sc_hd__a21o_2 _23984_ (.A1(_03336_),
    .A2(_03340_),
    .B1(_03341_),
    .X(_03342_));
 sky130_fd_sc_hd__nor2_4 _23985_ (.A(_03024_),
    .B(_03025_),
    .Y(_03343_));
 sky130_fd_sc_hd__nor2_2 _23986_ (.A(_03343_),
    .B(_03149_),
    .Y(_03344_));
 sky130_fd_sc_hd__and2_1 _23987_ (.A(_03342_),
    .B(_03344_),
    .X(_03345_));
 sky130_fd_sc_hd__nor2_1 _23988_ (.A(net1017),
    .B(_03161_),
    .Y(_03346_));
 sky130_fd_sc_hd__o211a_1 _23989_ (.A1(_03317_),
    .A2(_03318_),
    .B1(_03313_),
    .C1(_03315_),
    .X(_03347_));
 sky130_fd_sc_hd__a21o_1 _23990_ (.A1(_03317_),
    .A2(_03318_),
    .B1(_03347_),
    .X(_03348_));
 sky130_fd_sc_hd__xnor2_2 _23991_ (.A(_03346_),
    .B(_03348_),
    .Y(_03349_));
 sky130_fd_sc_hd__xnor2_2 _23992_ (.A(_03345_),
    .B(_03349_),
    .Y(_03350_));
 sky130_fd_sc_hd__nand2_1 _23993_ (.A(_03337_),
    .B(_03338_),
    .Y(_03351_));
 sky130_fd_sc_hd__xnor2_1 _23994_ (.A(_03336_),
    .B(_03339_),
    .Y(_03352_));
 sky130_fd_sc_hd__xnor2_2 _23995_ (.A(_03351_),
    .B(_03352_),
    .Y(_03353_));
 sky130_fd_sc_hd__o22a_2 _23996_ (.A1(_02993_),
    .A2(_02995_),
    .B1(_03063_),
    .B2(_03064_),
    .X(_03354_));
 sky130_fd_sc_hd__clkbuf_4 _23997_ (.A(_03040_),
    .X(_03355_));
 sky130_fd_sc_hd__o22a_1 _23998_ (.A1(_02976_),
    .A2(_02977_),
    .B1(_03057_),
    .B2(_03058_),
    .X(_03356_));
 sky130_fd_sc_hd__a21o_1 _23999_ (.A1(_03355_),
    .A2(_03216_),
    .B1(_03356_),
    .X(_03357_));
 sky130_fd_sc_hd__a32oi_4 _24000_ (.A1(_03305_),
    .A2(_03217_),
    .A3(_03060_),
    .B1(_03354_),
    .B2(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__or2_1 _24001_ (.A(_03353_),
    .B(_03358_),
    .X(_03359_));
 sky130_fd_sc_hd__xor2_2 _24002_ (.A(_03306_),
    .B(_03303_),
    .X(_03360_));
 sky130_fd_sc_hd__xnor2_4 _24003_ (.A(_03302_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__a21o_1 _24004_ (.A1(_03353_),
    .A2(_03358_),
    .B1(_03361_),
    .X(_03362_));
 sky130_fd_sc_hd__or2_2 _24005_ (.A(_03069_),
    .B(_03071_),
    .X(_03363_));
 sky130_fd_sc_hd__nor2_1 _24006_ (.A(_03325_),
    .B(_03106_),
    .Y(_03364_));
 sky130_fd_sc_hd__a31o_1 _24007_ (.A1(_03325_),
    .A2(_03363_),
    .A3(_03324_),
    .B1(_03364_),
    .X(_03365_));
 sky130_fd_sc_hd__a21o_1 _24008_ (.A1(_03363_),
    .A2(_03324_),
    .B1(_03056_),
    .X(_03366_));
 sky130_fd_sc_hd__or3_1 _24009_ (.A(_03195_),
    .B(_03250_),
    .C(_03217_),
    .X(_03367_));
 sky130_fd_sc_hd__a21oi_1 _24010_ (.A1(_03366_),
    .A2(_03367_),
    .B1(_03248_),
    .Y(_03368_));
 sky130_fd_sc_hd__a22o_1 _24011_ (.A1(_03056_),
    .A2(_03217_),
    .B1(_03363_),
    .B2(_03324_),
    .X(_03369_));
 sky130_fd_sc_hd__a21oi_1 _24012_ (.A1(_03253_),
    .A2(_03369_),
    .B1(_03323_),
    .Y(_03370_));
 sky130_fd_sc_hd__a311o_2 _24013_ (.A1(_03248_),
    .A2(_03323_),
    .A3(_03365_),
    .B1(_03368_),
    .C1(_03370_),
    .X(_03371_));
 sky130_fd_sc_hd__a21o_1 _24014_ (.A1(_03359_),
    .A2(_03362_),
    .B1(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__xnor2_2 _24015_ (.A(_03308_),
    .B(_03311_),
    .Y(_03373_));
 sky130_fd_sc_hd__xnor2_4 _24016_ (.A(_03320_),
    .B(_03373_),
    .Y(_03374_));
 sky130_fd_sc_hd__nand3_1 _24017_ (.A(_03359_),
    .B(_03362_),
    .C(_03371_),
    .Y(_03375_));
 sky130_fd_sc_hd__a21bo_1 _24018_ (.A1(_03372_),
    .A2(_03374_),
    .B1_N(_03375_),
    .X(_03376_));
 sky130_fd_sc_hd__xnor2_1 _24019_ (.A(_03350_),
    .B(_03376_),
    .Y(_03377_));
 sky130_fd_sc_hd__xnor2_2 _24020_ (.A(_03335_),
    .B(_03377_),
    .Y(_03378_));
 sky130_fd_sc_hd__nor2_2 _24021_ (.A(_02982_),
    .B(_03161_),
    .Y(_03379_));
 sky130_fd_sc_hd__o22a_1 _24022_ (.A1(_03036_),
    .A2(_03037_),
    .B1(_03045_),
    .B2(_03046_),
    .X(_03380_));
 sky130_fd_sc_hd__o22a_1 _24023_ (.A1(_02998_),
    .A2(_03000_),
    .B1(_03027_),
    .B2(_03028_),
    .X(_03381_));
 sky130_fd_sc_hd__o211a_1 _24024_ (.A1(_03380_),
    .A2(_03381_),
    .B1(_03010_),
    .C1(_03157_),
    .X(_03382_));
 sky130_fd_sc_hd__a21o_2 _24025_ (.A1(_03380_),
    .A2(_03381_),
    .B1(_03382_),
    .X(_03383_));
 sky130_fd_sc_hd__and2_2 _24026_ (.A(_03379_),
    .B(_03383_),
    .X(_03384_));
 sky130_fd_sc_hd__nand2_1 _24027_ (.A(_03010_),
    .B(_03157_),
    .Y(_03385_));
 sky130_fd_sc_hd__xnor2_1 _24028_ (.A(_03380_),
    .B(_03381_),
    .Y(_03386_));
 sky130_fd_sc_hd__xnor2_2 _24029_ (.A(_03385_),
    .B(_03386_),
    .Y(_03387_));
 sky130_fd_sc_hd__o22a_1 _24030_ (.A1(_02985_),
    .A2(_02987_),
    .B1(_03063_),
    .B2(_03064_),
    .X(_03388_));
 sky130_fd_sc_hd__o22a_2 _24031_ (.A1(_02976_),
    .A2(_02977_),
    .B1(_03076_),
    .B2(_03077_),
    .X(_03389_));
 sky130_fd_sc_hd__o22a_2 _24032_ (.A1(_02994_),
    .A2(_02996_),
    .B1(_03088_),
    .B2(_03089_),
    .X(_03390_));
 sky130_fd_sc_hd__a21o_1 _24033_ (.A1(_03388_),
    .A2(_03389_),
    .B1(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__o21ai_2 _24034_ (.A1(_03388_),
    .A2(_03389_),
    .B1(_03391_),
    .Y(_03392_));
 sky130_fd_sc_hd__or2_1 _24035_ (.A(_03387_),
    .B(_03392_),
    .X(_03393_));
 sky130_fd_sc_hd__nand2_2 _24036_ (.A(_03355_),
    .B(_03217_),
    .Y(_03394_));
 sky130_fd_sc_hd__xnor2_2 _24037_ (.A(_03354_),
    .B(_03356_),
    .Y(_03395_));
 sky130_fd_sc_hd__xnor2_4 _24038_ (.A(_03394_),
    .B(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__a21o_1 _24039_ (.A1(_03387_),
    .A2(_03392_),
    .B1(_03396_),
    .X(_03397_));
 sky130_fd_sc_hd__and2_1 _24040_ (.A(_03393_),
    .B(_03397_),
    .X(_03398_));
 sky130_fd_sc_hd__xnor2_2 _24041_ (.A(_03353_),
    .B(_03358_),
    .Y(_03399_));
 sky130_fd_sc_hd__xnor2_4 _24042_ (.A(_03361_),
    .B(_03399_),
    .Y(_03400_));
 sky130_fd_sc_hd__nor2_1 _24043_ (.A(_03398_),
    .B(_03400_),
    .Y(_03401_));
 sky130_fd_sc_hd__xnor2_4 _24044_ (.A(_03342_),
    .B(_03344_),
    .Y(_03402_));
 sky130_fd_sc_hd__o21ba_1 _24045_ (.A1(_03384_),
    .A2(_03401_),
    .B1_N(_03402_),
    .X(_03403_));
 sky130_fd_sc_hd__o211a_1 _24046_ (.A1(_03195_),
    .A2(_03254_),
    .B1(_03324_),
    .C1(_03056_),
    .X(_03404_));
 sky130_fd_sc_hd__o211a_1 _24047_ (.A1(_03250_),
    .A2(_03252_),
    .B1(_03363_),
    .C1(_03120_),
    .X(_03405_));
 sky130_fd_sc_hd__nor2_1 _24048_ (.A(_03404_),
    .B(_03405_),
    .Y(_03406_));
 sky130_fd_sc_hd__a21o_1 _24049_ (.A1(_03393_),
    .A2(_03397_),
    .B1(_03406_),
    .X(_03407_));
 sky130_fd_sc_hd__and3_1 _24050_ (.A(_03393_),
    .B(_03397_),
    .C(_03406_),
    .X(_03408_));
 sky130_fd_sc_hd__a21oi_2 _24051_ (.A1(_03400_),
    .A2(_03407_),
    .B1(_03408_),
    .Y(_03409_));
 sky130_fd_sc_hd__xnor2_4 _24052_ (.A(_03384_),
    .B(_03402_),
    .Y(_03410_));
 sky130_fd_sc_hd__nand2_1 _24053_ (.A(_03398_),
    .B(_03400_),
    .Y(_03411_));
 sky130_fd_sc_hd__o211a_1 _24054_ (.A1(_03404_),
    .A2(_03405_),
    .B1(_03410_),
    .C1(_03411_),
    .X(_03412_));
 sky130_fd_sc_hd__nand3_2 _24055_ (.A(_03372_),
    .B(_03374_),
    .C(_03375_),
    .Y(_03413_));
 sky130_fd_sc_hd__a21o_1 _24056_ (.A1(_03372_),
    .A2(_03375_),
    .B1(_03374_),
    .X(_03414_));
 sky130_fd_sc_hd__nand2_1 _24057_ (.A(_03413_),
    .B(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__nand2_1 _24058_ (.A(_03401_),
    .B(_03410_),
    .Y(_03416_));
 sky130_fd_sc_hd__o221a_1 _24059_ (.A1(_03409_),
    .A2(_03410_),
    .B1(_03412_),
    .B2(_03415_),
    .C1(_03416_),
    .X(_03417_));
 sky130_fd_sc_hd__a211o_1 _24060_ (.A1(_03384_),
    .A2(_03401_),
    .B1(_03403_),
    .C1(_03417_),
    .X(_03418_));
 sky130_fd_sc_hd__and2b_1 _24061_ (.A_N(_03402_),
    .B(_03384_),
    .X(_03419_));
 sky130_fd_sc_hd__inv_2 _24062_ (.A(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__a21o_1 _24063_ (.A1(_03400_),
    .A2(_03407_),
    .B1(_03408_),
    .X(_03421_));
 sky130_fd_sc_hd__a211o_1 _24064_ (.A1(_03413_),
    .A2(_03414_),
    .B1(_03420_),
    .C1(_03421_),
    .X(_03422_));
 sky130_fd_sc_hd__a21boi_1 _24065_ (.A1(_03378_),
    .A2(_03418_),
    .B1_N(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__inv_2 _24066_ (.A(_03350_),
    .Y(_03424_));
 sky130_fd_sc_hd__o21a_1 _24067_ (.A1(_03424_),
    .A2(_03371_),
    .B1(_03335_),
    .X(_03425_));
 sky130_fd_sc_hd__and2_1 _24068_ (.A(_03359_),
    .B(_03362_),
    .X(_03426_));
 sky130_fd_sc_hd__and3_1 _24069_ (.A(_03335_),
    .B(_03426_),
    .C(_03374_),
    .X(_03427_));
 sky130_fd_sc_hd__nor2_1 _24070_ (.A(_03426_),
    .B(_03374_),
    .Y(_03428_));
 sky130_fd_sc_hd__o211a_1 _24071_ (.A1(_03426_),
    .A2(_03374_),
    .B1(_03371_),
    .C1(_03424_),
    .X(_03429_));
 sky130_fd_sc_hd__and3_1 _24072_ (.A(_03424_),
    .B(_03426_),
    .C(_03374_),
    .X(_03430_));
 sky130_fd_sc_hd__a211o_1 _24073_ (.A1(_03350_),
    .A2(_03428_),
    .B1(_03429_),
    .C1(_03430_),
    .X(_03431_));
 sky130_fd_sc_hd__nor3_1 _24074_ (.A(_03425_),
    .B(_03427_),
    .C(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__a21bo_1 _24075_ (.A1(_03345_),
    .A2(_03428_),
    .B1_N(_03349_),
    .X(_03433_));
 sky130_fd_sc_hd__o21a_1 _24076_ (.A1(_03345_),
    .A2(_03428_),
    .B1(_03433_),
    .X(_03434_));
 sky130_fd_sc_hd__xnor2_2 _24077_ (.A(_03231_),
    .B(_03269_),
    .Y(_03435_));
 sky130_fd_sc_hd__xnor2_4 _24078_ (.A(_03266_),
    .B(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__a21oi_1 _24079_ (.A1(_03312_),
    .A2(_03321_),
    .B1(_03327_),
    .Y(_03437_));
 sky130_fd_sc_hd__o21ai_2 _24080_ (.A1(_03437_),
    .A2(_03332_),
    .B1(_03329_),
    .Y(_03438_));
 sky130_fd_sc_hd__nand2_1 _24081_ (.A(_03346_),
    .B(_03348_),
    .Y(_03439_));
 sky130_fd_sc_hd__xnor2_2 _24082_ (.A(_03279_),
    .B(_03281_),
    .Y(_03440_));
 sky130_fd_sc_hd__xnor2_1 _24083_ (.A(_03439_),
    .B(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__xnor2_2 _24084_ (.A(_03438_),
    .B(_03441_),
    .Y(_03442_));
 sky130_fd_sc_hd__and3_1 _24085_ (.A(_03328_),
    .B(_03329_),
    .C(_03332_),
    .X(_03443_));
 sky130_fd_sc_hd__a21oi_1 _24086_ (.A1(_03328_),
    .A2(_03329_),
    .B1(_03332_),
    .Y(_03444_));
 sky130_fd_sc_hd__or3_2 _24087_ (.A(_03333_),
    .B(_03443_),
    .C(_03444_),
    .X(_03445_));
 sky130_fd_sc_hd__xor2_2 _24088_ (.A(_03442_),
    .B(_03445_),
    .X(_03446_));
 sky130_fd_sc_hd__xnor2_4 _24089_ (.A(_03436_),
    .B(_03446_),
    .Y(_03447_));
 sky130_fd_sc_hd__xor2_1 _24090_ (.A(_03434_),
    .B(_03447_),
    .X(_03448_));
 sky130_fd_sc_hd__xnor2_1 _24091_ (.A(_03432_),
    .B(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__and2_1 _24092_ (.A(_03423_),
    .B(_03449_),
    .X(_03450_));
 sky130_fd_sc_hd__or2b_1 _24093_ (.A(_03384_),
    .B_N(_03402_),
    .X(_03451_));
 sky130_fd_sc_hd__o21a_1 _24094_ (.A1(_03419_),
    .A2(_03409_),
    .B1(_03451_),
    .X(_03452_));
 sky130_fd_sc_hd__o221a_1 _24095_ (.A1(_03451_),
    .A2(_03409_),
    .B1(_03452_),
    .B2(_03415_),
    .C1(_03422_),
    .X(_03453_));
 sky130_fd_sc_hd__xor2_2 _24096_ (.A(_03378_),
    .B(_03453_),
    .X(_03454_));
 sky130_fd_sc_hd__inv_2 _24097_ (.A(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__xnor2_4 _24098_ (.A(_03379_),
    .B(_03383_),
    .Y(_03456_));
 sky130_fd_sc_hd__nor2_2 _24099_ (.A(_03006_),
    .B(_03185_),
    .Y(_03457_));
 sky130_fd_sc_hd__o22a_1 _24100_ (.A1(_03045_),
    .A2(_03046_),
    .B1(_03057_),
    .B2(_03058_),
    .X(_03458_));
 sky130_fd_sc_hd__o22a_1 _24101_ (.A1(_03207_),
    .A2(_03208_),
    .B1(_03015_),
    .B2(_03016_),
    .X(_03459_));
 sky130_fd_sc_hd__xnor2_1 _24102_ (.A(_03458_),
    .B(_03459_),
    .Y(_03460_));
 sky130_fd_sc_hd__xnor2_2 _24103_ (.A(_03457_),
    .B(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__xor2_2 _24104_ (.A(_03389_),
    .B(_03390_),
    .X(_03462_));
 sky130_fd_sc_hd__nand2_1 _24105_ (.A(_03355_),
    .B(_03324_),
    .Y(_03463_));
 sky130_fd_sc_hd__nor2_2 _24106_ (.A(_02978_),
    .B(_03195_),
    .Y(_03464_));
 sky130_fd_sc_hd__or2_1 _24107_ (.A(_03463_),
    .B(_03464_),
    .X(_03465_));
 sky130_fd_sc_hd__nor2_1 _24108_ (.A(_03463_),
    .B(_03462_),
    .Y(_03466_));
 sky130_fd_sc_hd__a31o_1 _24109_ (.A1(_03305_),
    .A2(_03120_),
    .A3(_03324_),
    .B1(_03461_),
    .X(_03467_));
 sky130_fd_sc_hd__a32o_2 _24110_ (.A1(_03461_),
    .A2(_03462_),
    .A3(_03465_),
    .B1(_03466_),
    .B2(_03467_),
    .X(_03468_));
 sky130_fd_sc_hd__xor2_2 _24111_ (.A(_03387_),
    .B(_03392_),
    .X(_03469_));
 sky130_fd_sc_hd__xnor2_4 _24112_ (.A(_03396_),
    .B(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__nand2_2 _24113_ (.A(_03468_),
    .B(_03470_),
    .Y(_03471_));
 sky130_fd_sc_hd__o21a_1 _24114_ (.A1(_03458_),
    .A2(_03457_),
    .B1(_03459_),
    .X(_03472_));
 sky130_fd_sc_hd__a21o_1 _24115_ (.A1(_03458_),
    .A2(_03457_),
    .B1(_03472_),
    .X(_03473_));
 sky130_fd_sc_hd__nor2_4 _24116_ (.A(_02989_),
    .B(_02991_),
    .Y(_03474_));
 sky130_fd_sc_hd__nor2_1 _24117_ (.A(_03474_),
    .B(_03161_),
    .Y(_03475_));
 sky130_fd_sc_hd__nand2_1 _24118_ (.A(_03473_),
    .B(_03475_),
    .Y(_03476_));
 sky130_fd_sc_hd__o21a_1 _24119_ (.A1(_03456_),
    .A2(_03471_),
    .B1(_03476_),
    .X(_03477_));
 sky130_fd_sc_hd__a21oi_4 _24120_ (.A1(_03456_),
    .A2(_03471_),
    .B1(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__a21oi_1 _24121_ (.A1(_03393_),
    .A2(_03397_),
    .B1(_03406_),
    .Y(_03479_));
 sky130_fd_sc_hd__or3_1 _24122_ (.A(_03400_),
    .B(_03479_),
    .C(_03408_),
    .X(_03480_));
 sky130_fd_sc_hd__o21ai_1 _24123_ (.A1(_03479_),
    .A2(_03408_),
    .B1(_03400_),
    .Y(_03481_));
 sky130_fd_sc_hd__and2_1 _24124_ (.A(_03480_),
    .B(_03481_),
    .X(_03482_));
 sky130_fd_sc_hd__nand2_1 _24125_ (.A(_03323_),
    .B(_03056_),
    .Y(_03483_));
 sky130_fd_sc_hd__o21ba_1 _24126_ (.A1(_03468_),
    .A2(_03470_),
    .B1_N(_03483_),
    .X(_03484_));
 sky130_fd_sc_hd__and2_1 _24127_ (.A(_03468_),
    .B(_03470_),
    .X(_03485_));
 sky130_fd_sc_hd__o211a_1 _24128_ (.A1(_03485_),
    .A2(_03484_),
    .B1(_03481_),
    .C1(_03480_),
    .X(_03486_));
 sky130_fd_sc_hd__xor2_2 _24129_ (.A(_03476_),
    .B(_03456_),
    .X(_03487_));
 sky130_fd_sc_hd__nand2_1 _24130_ (.A(_03485_),
    .B(_03487_),
    .Y(_03488_));
 sky130_fd_sc_hd__o221a_2 _24131_ (.A1(_03482_),
    .A2(_03484_),
    .B1(_03486_),
    .B2(_03487_),
    .C1(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__xnor2_2 _24132_ (.A(_03473_),
    .B(_03475_),
    .Y(_03490_));
 sky130_fd_sc_hd__o22a_1 _24133_ (.A1(_03036_),
    .A2(_03037_),
    .B1(_03027_),
    .B2(_03028_),
    .X(_03491_));
 sky130_fd_sc_hd__o22a_1 _24134_ (.A1(_03045_),
    .A2(_03046_),
    .B1(_03076_),
    .B2(_03077_),
    .X(_03492_));
 sky130_fd_sc_hd__nor2_1 _24135_ (.A(_03491_),
    .B(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__nand2_1 _24136_ (.A(_03491_),
    .B(_03492_),
    .Y(_03494_));
 sky130_fd_sc_hd__o31ai_4 _24137_ (.A1(_03017_),
    .A2(_03114_),
    .A3(_03493_),
    .B1(_03494_),
    .Y(_03495_));
 sky130_fd_sc_hd__nor2_2 _24138_ (.A(_02998_),
    .B(_03000_),
    .Y(_03496_));
 sky130_fd_sc_hd__nor2_2 _24139_ (.A(_03496_),
    .B(_03161_),
    .Y(_03497_));
 sky130_fd_sc_hd__nand2_1 _24140_ (.A(_03495_),
    .B(_03497_),
    .Y(_03498_));
 sky130_fd_sc_hd__xnor2_1 _24141_ (.A(_03462_),
    .B(_03465_),
    .Y(_03499_));
 sky130_fd_sc_hd__xnor2_1 _24142_ (.A(_03461_),
    .B(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hd__or2_1 _24143_ (.A(_02976_),
    .B(_02977_),
    .X(_03501_));
 sky130_fd_sc_hd__clkbuf_4 _24144_ (.A(_03501_),
    .X(_03502_));
 sky130_fd_sc_hd__o211a_1 _24145_ (.A1(_03234_),
    .A2(_03195_),
    .B1(_03121_),
    .C1(_03502_),
    .X(_03503_));
 sky130_fd_sc_hd__o211a_1 _24146_ (.A1(_02978_),
    .A2(_03252_),
    .B1(_03120_),
    .C1(_03355_),
    .X(_03504_));
 sky130_fd_sc_hd__nor2_2 _24147_ (.A(_03503_),
    .B(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__nand2_1 _24148_ (.A(_03157_),
    .B(_03060_),
    .Y(_03506_));
 sky130_fd_sc_hd__xnor2_1 _24149_ (.A(_03491_),
    .B(_03492_),
    .Y(_03507_));
 sky130_fd_sc_hd__xnor2_2 _24150_ (.A(_03506_),
    .B(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__or3_2 _24151_ (.A(_03500_),
    .B(_03505_),
    .C(_03508_),
    .X(_03509_));
 sky130_fd_sc_hd__o21a_1 _24152_ (.A1(_03490_),
    .A2(_03498_),
    .B1(_03509_),
    .X(_03510_));
 sky130_fd_sc_hd__a21o_1 _24153_ (.A1(_03490_),
    .A2(_03498_),
    .B1(_03510_),
    .X(_03511_));
 sky130_fd_sc_hd__xnor2_1 _24154_ (.A(_03483_),
    .B(_03468_),
    .Y(_03512_));
 sky130_fd_sc_hd__xnor2_2 _24155_ (.A(_03470_),
    .B(_03512_),
    .Y(_03513_));
 sky130_fd_sc_hd__xnor2_1 _24156_ (.A(_03490_),
    .B(_03498_),
    .Y(_03514_));
 sky130_fd_sc_hd__xnor2_1 _24157_ (.A(_03509_),
    .B(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__or2_2 _24158_ (.A(_03513_),
    .B(_03515_),
    .X(_03516_));
 sky130_fd_sc_hd__o21bai_1 _24159_ (.A1(_03468_),
    .A2(_03470_),
    .B1_N(_03483_),
    .Y(_03517_));
 sky130_fd_sc_hd__and3_1 _24160_ (.A(_03471_),
    .B(_03517_),
    .C(_03487_),
    .X(_03518_));
 sky130_fd_sc_hd__a21oi_1 _24161_ (.A1(_03471_),
    .A2(_03517_),
    .B1(_03487_),
    .Y(_03519_));
 sky130_fd_sc_hd__nor2_1 _24162_ (.A(_03518_),
    .B(_03519_),
    .Y(_03520_));
 sky130_fd_sc_hd__or3_1 _24163_ (.A(_03509_),
    .B(_03490_),
    .C(_03498_),
    .X(_03521_));
 sky130_fd_sc_hd__o21ba_1 _24164_ (.A1(_03513_),
    .A2(_03521_),
    .B1_N(_03482_),
    .X(_03522_));
 sky130_fd_sc_hd__o221a_1 _24165_ (.A1(_03518_),
    .A2(_03519_),
    .B1(_03521_),
    .B2(_03513_),
    .C1(_03482_),
    .X(_03523_));
 sky130_fd_sc_hd__a221oi_4 _24166_ (.A1(_03511_),
    .A2(_03516_),
    .B1(_03520_),
    .B2(_03522_),
    .C1(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__a21o_1 _24167_ (.A1(_03478_),
    .A2(_03489_),
    .B1(_03524_),
    .X(_03525_));
 sky130_fd_sc_hd__a21oi_1 _24168_ (.A1(_03398_),
    .A2(_03400_),
    .B1(_03410_),
    .Y(_03526_));
 sky130_fd_sc_hd__o21ai_1 _24169_ (.A1(_03398_),
    .A2(_03400_),
    .B1(_03406_),
    .Y(_03527_));
 sky130_fd_sc_hd__mux2_1 _24170_ (.A0(_03410_),
    .A1(_03526_),
    .S(_03527_),
    .X(_03528_));
 sky130_fd_sc_hd__inv_2 _24171_ (.A(_03410_),
    .Y(_03529_));
 sky130_fd_sc_hd__o211ai_1 _24172_ (.A1(_03411_),
    .A2(_03529_),
    .B1(_03413_),
    .C1(_03414_),
    .Y(_03530_));
 sky130_fd_sc_hd__a32o_1 _24173_ (.A1(_03411_),
    .A2(_03527_),
    .A3(_03410_),
    .B1(_03414_),
    .B2(_03413_),
    .X(_03531_));
 sky130_fd_sc_hd__nor2_1 _24174_ (.A(_03409_),
    .B(_03410_),
    .Y(_03532_));
 sky130_fd_sc_hd__o22a_2 _24175_ (.A1(_03528_),
    .A2(_03530_),
    .B1(_03531_),
    .B2(_03532_),
    .X(_03533_));
 sky130_fd_sc_hd__o21a_1 _24176_ (.A1(_03478_),
    .A2(_03489_),
    .B1(_03533_),
    .X(_03534_));
 sky130_fd_sc_hd__or3_1 _24177_ (.A(_03478_),
    .B(_03489_),
    .C(_03533_),
    .X(_03535_));
 sky130_fd_sc_hd__nand2_1 _24178_ (.A(_03478_),
    .B(_03533_),
    .Y(_03536_));
 sky130_fd_sc_hd__o21ai_1 _24179_ (.A1(_03478_),
    .A2(_03533_),
    .B1(_03489_),
    .Y(_03537_));
 sky130_fd_sc_hd__o2111a_1 _24180_ (.A1(_03524_),
    .A2(_03535_),
    .B1(_03536_),
    .C1(_03537_),
    .D1(_03454_),
    .X(_03538_));
 sky130_fd_sc_hd__a31o_1 _24181_ (.A1(_03455_),
    .A2(_03525_),
    .A3(_03534_),
    .B1(_03538_),
    .X(_03539_));
 sky130_fd_sc_hd__xnor2_2 _24182_ (.A(_03505_),
    .B(_03508_),
    .Y(_03540_));
 sky130_fd_sc_hd__nor2_1 _24183_ (.A(_03185_),
    .B(_03114_),
    .Y(_03541_));
 sky130_fd_sc_hd__o22a_1 _24184_ (.A1(_03015_),
    .A2(_03016_),
    .B1(_03076_),
    .B2(_03077_),
    .X(_03542_));
 sky130_fd_sc_hd__o22a_1 _24185_ (.A1(_03045_),
    .A2(_03046_),
    .B1(_03063_),
    .B2(_03064_),
    .X(_03543_));
 sky130_fd_sc_hd__xnor2_1 _24186_ (.A(_03542_),
    .B(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__xnor2_2 _24187_ (.A(_03541_),
    .B(_03544_),
    .Y(_03545_));
 sky130_fd_sc_hd__nand2_2 _24188_ (.A(_03464_),
    .B(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__nor2_1 _24189_ (.A(_03540_),
    .B(_03546_),
    .Y(_03547_));
 sky130_fd_sc_hd__xnor2_2 _24190_ (.A(_03495_),
    .B(_03497_),
    .Y(_03548_));
 sky130_fd_sc_hd__a22o_4 _24191_ (.A1(\top0.matmul0.matmul_stage_inst.f[0] ),
    .A2(_03146_),
    .B1(_03148_),
    .B2(\top0.matmul0.matmul_stage_inst.e[0] ),
    .X(_03549_));
 sky130_fd_sc_hd__nor2_1 _24192_ (.A(_03542_),
    .B(_03543_),
    .Y(_03550_));
 sky130_fd_sc_hd__nand2_1 _24193_ (.A(_03542_),
    .B(_03543_),
    .Y(_03551_));
 sky130_fd_sc_hd__o31ai_2 _24194_ (.A1(_03185_),
    .A2(_03114_),
    .A3(_03550_),
    .B1(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__and3_1 _24195_ (.A(_03010_),
    .B(_03549_),
    .C(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__xor2_1 _24196_ (.A(_03548_),
    .B(_03553_),
    .X(_03554_));
 sky130_fd_sc_hd__xnor2_1 _24197_ (.A(_03547_),
    .B(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__nor2_1 _24198_ (.A(_03505_),
    .B(_03508_),
    .Y(_03556_));
 sky130_fd_sc_hd__xnor2_1 _24199_ (.A(_03500_),
    .B(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__xor2_1 _24200_ (.A(_03555_),
    .B(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__xor2_2 _24201_ (.A(_03540_),
    .B(_03546_),
    .X(_03559_));
 sky130_fd_sc_hd__a22o_1 _24202_ (.A1(_03315_),
    .A2(_03323_),
    .B1(_03217_),
    .B2(_03337_),
    .X(_03560_));
 sky130_fd_sc_hd__nor2_1 _24203_ (.A(_03017_),
    .B(_03252_),
    .Y(_03561_));
 sky130_fd_sc_hd__and4_1 _24204_ (.A(_03315_),
    .B(_03337_),
    .C(_03323_),
    .D(_03217_),
    .X(_03562_));
 sky130_fd_sc_hd__a21o_1 _24205_ (.A1(_03560_),
    .A2(_03561_),
    .B1(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__nor2_2 _24206_ (.A(_03207_),
    .B(_03208_),
    .Y(_03564_));
 sky130_fd_sc_hd__nor2_1 _24207_ (.A(_03564_),
    .B(_03161_),
    .Y(_03565_));
 sky130_fd_sc_hd__and2_1 _24208_ (.A(_03563_),
    .B(_03565_),
    .X(_03566_));
 sky130_fd_sc_hd__nand2_1 _24209_ (.A(_03010_),
    .B(_03549_),
    .Y(_03567_));
 sky130_fd_sc_hd__xnor2_2 _24210_ (.A(_03567_),
    .B(_03552_),
    .Y(_03568_));
 sky130_fd_sc_hd__a21o_1 _24211_ (.A1(_03559_),
    .A2(_03566_),
    .B1(_03568_),
    .X(_03569_));
 sky130_fd_sc_hd__o21a_1 _24212_ (.A1(_03559_),
    .A2(_03566_),
    .B1(_03569_),
    .X(_03570_));
 sky130_fd_sc_hd__o211a_1 _24213_ (.A1(_03185_),
    .A2(_03106_),
    .B1(_03323_),
    .C1(_03315_),
    .X(_03571_));
 sky130_fd_sc_hd__buf_2 _24214_ (.A(_03337_),
    .X(_03572_));
 sky130_fd_sc_hd__o211a_1 _24215_ (.A1(_03047_),
    .A2(_03195_),
    .B1(_03217_),
    .C1(_03572_),
    .X(_03573_));
 sky130_fd_sc_hd__nor2_1 _24216_ (.A(_03571_),
    .B(_03573_),
    .Y(_03574_));
 sky130_fd_sc_hd__xnor2_1 _24217_ (.A(_03561_),
    .B(_03574_),
    .Y(_03575_));
 sky130_fd_sc_hd__and3_1 _24218_ (.A(_03572_),
    .B(_03323_),
    .C(_03561_),
    .X(_03576_));
 sky130_fd_sc_hd__nor2_1 _24219_ (.A(_03114_),
    .B(_03161_),
    .Y(_03577_));
 sky130_fd_sc_hd__xor2_1 _24220_ (.A(_03576_),
    .B(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__a21o_1 _24221_ (.A1(_03017_),
    .A2(_03323_),
    .B1(_03217_),
    .X(_03579_));
 sky130_fd_sc_hd__a32o_1 _24222_ (.A1(_03572_),
    .A2(_03324_),
    .A3(_03579_),
    .B1(_03542_),
    .B2(_03323_),
    .X(_03580_));
 sky130_fd_sc_hd__a22o_1 _24223_ (.A1(_03549_),
    .A2(_03580_),
    .B1(_03578_),
    .B2(_03575_),
    .X(_03581_));
 sky130_fd_sc_hd__o21a_1 _24224_ (.A1(_03575_),
    .A2(_03578_),
    .B1(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__and2_1 _24225_ (.A(_03576_),
    .B(_03577_),
    .X(_03583_));
 sky130_fd_sc_hd__xor2_1 _24226_ (.A(_03565_),
    .B(_03583_),
    .X(_03584_));
 sky130_fd_sc_hd__xor2_2 _24227_ (.A(_03464_),
    .B(_03545_),
    .X(_03585_));
 sky130_fd_sc_hd__and2_1 _24228_ (.A(_03563_),
    .B(_03585_),
    .X(_03586_));
 sky130_fd_sc_hd__nor2_1 _24229_ (.A(_03563_),
    .B(_03585_),
    .Y(_03587_));
 sky130_fd_sc_hd__xor2_2 _24230_ (.A(_03559_),
    .B(_03568_),
    .X(_03588_));
 sky130_fd_sc_hd__mux2_1 _24231_ (.A0(_03586_),
    .A1(_03587_),
    .S(_03588_),
    .X(_03589_));
 sky130_fd_sc_hd__nor2_1 _24232_ (.A(_03586_),
    .B(_03587_),
    .Y(_03590_));
 sky130_fd_sc_hd__and3_1 _24233_ (.A(_03565_),
    .B(_03576_),
    .C(_03577_),
    .X(_03591_));
 sky130_fd_sc_hd__nor2_1 _24234_ (.A(_03565_),
    .B(_03583_),
    .Y(_03592_));
 sky130_fd_sc_hd__mux2_1 _24235_ (.A0(_03591_),
    .A1(_03592_),
    .S(_03588_),
    .X(_03593_));
 sky130_fd_sc_hd__a22o_1 _24236_ (.A1(_03584_),
    .A2(_03589_),
    .B1(_03590_),
    .B2(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__and3_1 _24237_ (.A(_03566_),
    .B(_03583_),
    .C(_03585_),
    .X(_03595_));
 sky130_fd_sc_hd__or2_1 _24238_ (.A(_03583_),
    .B(_03585_),
    .X(_03596_));
 sky130_fd_sc_hd__a211o_1 _24239_ (.A1(_03583_),
    .A2(_03585_),
    .B1(_03563_),
    .C1(_03565_),
    .X(_03597_));
 sky130_fd_sc_hd__and3b_1 _24240_ (.A_N(_03566_),
    .B(_03596_),
    .C(_03597_),
    .X(_03598_));
 sky130_fd_sc_hd__mux2_1 _24241_ (.A0(_03595_),
    .A1(_03598_),
    .S(_03588_),
    .X(_03599_));
 sky130_fd_sc_hd__a221o_1 _24242_ (.A1(_03558_),
    .A2(_03570_),
    .B1(_03582_),
    .B2(_03594_),
    .C1(_03599_),
    .X(_03600_));
 sky130_fd_sc_hd__or2_1 _24243_ (.A(_03558_),
    .B(_03570_),
    .X(_03601_));
 sky130_fd_sc_hd__xor2_1 _24244_ (.A(_03513_),
    .B(_03515_),
    .X(_03602_));
 sky130_fd_sc_hd__and2_1 _24245_ (.A(_03555_),
    .B(_03557_),
    .X(_03603_));
 sky130_fd_sc_hd__a211o_1 _24246_ (.A1(_03600_),
    .A2(_03601_),
    .B1(_03602_),
    .C1(_03603_),
    .X(_03604_));
 sky130_fd_sc_hd__a22o_1 _24247_ (.A1(_03603_),
    .A2(_03570_),
    .B1(_03601_),
    .B2(_03602_),
    .X(_03605_));
 sky130_fd_sc_hd__o21ai_1 _24248_ (.A1(_03540_),
    .A2(_03546_),
    .B1(_03548_),
    .Y(_03606_));
 sky130_fd_sc_hd__and2b_1 _24249_ (.A_N(_03548_),
    .B(_03547_),
    .X(_03607_));
 sky130_fd_sc_hd__a221o_1 _24250_ (.A1(_03603_),
    .A2(_03602_),
    .B1(_03606_),
    .B2(_03553_),
    .C1(_03607_),
    .X(_03608_));
 sky130_fd_sc_hd__a21o_1 _24251_ (.A1(_03600_),
    .A2(_03605_),
    .B1(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__xnor2_1 _24252_ (.A(_03482_),
    .B(_03520_),
    .Y(_03610_));
 sky130_fd_sc_hd__xor2_1 _24253_ (.A(_03511_),
    .B(_03516_),
    .X(_03611_));
 sky130_fd_sc_hd__xor2_1 _24254_ (.A(_03610_),
    .B(_03611_),
    .X(_03612_));
 sky130_fd_sc_hd__xnor2_1 _24255_ (.A(_03478_),
    .B(_03489_),
    .Y(_03613_));
 sky130_fd_sc_hd__xnor2_1 _24256_ (.A(_03533_),
    .B(_03613_),
    .Y(_03614_));
 sky130_fd_sc_hd__a32o_1 _24257_ (.A1(_03604_),
    .A2(_03609_),
    .A3(_03612_),
    .B1(_03614_),
    .B2(_03524_),
    .X(_03615_));
 sky130_fd_sc_hd__nand2_1 _24258_ (.A(_03536_),
    .B(_03537_),
    .Y(_03616_));
 sky130_fd_sc_hd__a21boi_1 _24259_ (.A1(_03454_),
    .A2(_03616_),
    .B1_N(_03423_),
    .Y(_03617_));
 sky130_fd_sc_hd__o2bb2a_1 _24260_ (.A1_N(_03539_),
    .A2_N(_03615_),
    .B1(_03617_),
    .B2(_03449_),
    .X(_03618_));
 sky130_fd_sc_hd__a21o_1 _24261_ (.A1(_03439_),
    .A2(_03440_),
    .B1(_03438_),
    .X(_03619_));
 sky130_fd_sc_hd__o21a_1 _24262_ (.A1(_03439_),
    .A2(_03440_),
    .B1(_03619_),
    .X(_03620_));
 sky130_fd_sc_hd__o21a_1 _24263_ (.A1(_03442_),
    .A2(_03436_),
    .B1(_03445_),
    .X(_03621_));
 sky130_fd_sc_hd__a21o_1 _24264_ (.A1(_03442_),
    .A2(_03436_),
    .B1(_03621_),
    .X(_03622_));
 sky130_fd_sc_hd__nand2_1 _24265_ (.A(_03620_),
    .B(_03622_),
    .Y(_03623_));
 sky130_fd_sc_hd__nand2_2 _24266_ (.A(net8),
    .B(_03447_),
    .Y(_03624_));
 sky130_fd_sc_hd__o21ai_4 _24267_ (.A1(net8),
    .A2(_03447_),
    .B1(_03434_),
    .Y(_03625_));
 sky130_fd_sc_hd__and2_1 _24268_ (.A(_03624_),
    .B(_03625_),
    .X(_03626_));
 sky130_fd_sc_hd__or2b_1 _24269_ (.A(_03623_),
    .B_N(_03626_),
    .X(_03627_));
 sky130_fd_sc_hd__nand2_2 _24270_ (.A(_03293_),
    .B(_03294_),
    .Y(_03628_));
 sky130_fd_sc_hd__xnor2_4 _24271_ (.A(_03628_),
    .B(_03287_),
    .Y(_03629_));
 sky130_fd_sc_hd__xnor2_4 _24272_ (.A(_03290_),
    .B(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__or2_1 _24273_ (.A(_03620_),
    .B(_03622_),
    .X(_03631_));
 sky130_fd_sc_hd__a21bo_1 _24274_ (.A1(_03626_),
    .A2(_03631_),
    .B1_N(_03623_),
    .X(_03632_));
 sky130_fd_sc_hd__nand2_1 _24275_ (.A(_03630_),
    .B(_03632_),
    .Y(_03633_));
 sky130_fd_sc_hd__a2bb2o_1 _24276_ (.A1_N(_03450_),
    .A2_N(_03618_),
    .B1(_03627_),
    .B2(_03633_),
    .X(_03634_));
 sky130_fd_sc_hd__xor2_1 _24277_ (.A(_03290_),
    .B(_03629_),
    .X(_03635_));
 sky130_fd_sc_hd__or2_1 _24278_ (.A(_03627_),
    .B(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__or3_1 _24279_ (.A(_03626_),
    .B(_03630_),
    .C(_03631_),
    .X(_03637_));
 sky130_fd_sc_hd__or2_1 _24280_ (.A(_03630_),
    .B(_03632_),
    .X(_03638_));
 sky130_fd_sc_hd__or3_1 _24281_ (.A(_03450_),
    .B(_03618_),
    .C(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__and4_2 _24282_ (.A(_03634_),
    .B(_03636_),
    .C(_03637_),
    .D(_03639_),
    .X(_03640_));
 sky130_fd_sc_hd__xnor2_4 _24283_ (.A(_03301_),
    .B(_03640_),
    .Y(_03641_));
 sky130_fd_sc_hd__clkbuf_4 _24284_ (.A(_03146_),
    .X(_03642_));
 sky130_fd_sc_hd__mux2_1 _24285_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[0] ),
    .A1(_03641_),
    .S(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__clkbuf_1 _24286_ (.A(_03643_),
    .X(_00601_));
 sky130_fd_sc_hd__a2111oi_1 _24287_ (.A1(_03624_),
    .A2(_03625_),
    .B1(_03630_),
    .C1(_03300_),
    .D1(_03299_),
    .Y(_03644_));
 sky130_fd_sc_hd__o2111a_1 _24288_ (.A1(_03299_),
    .A2(_03300_),
    .B1(_03624_),
    .C1(_03625_),
    .D1(_03630_),
    .X(_03645_));
 sky130_fd_sc_hd__o211ai_1 _24289_ (.A1(_03644_),
    .A2(_03645_),
    .B1(_03623_),
    .C1(_03631_),
    .Y(_03646_));
 sky130_fd_sc_hd__a21oi_1 _24290_ (.A1(_03624_),
    .A2(_03625_),
    .B1(_03635_),
    .Y(_03647_));
 sky130_fd_sc_hd__and3_1 _24291_ (.A(_03624_),
    .B(_03625_),
    .C(_03635_),
    .X(_03648_));
 sky130_fd_sc_hd__o21bai_1 _24292_ (.A1(_03299_),
    .A2(_03300_),
    .B1_N(_03623_),
    .Y(_03649_));
 sky130_fd_sc_hd__or3_1 _24293_ (.A(_03299_),
    .B(_03300_),
    .C(_03631_),
    .X(_03650_));
 sky130_fd_sc_hd__a2bb2o_1 _24294_ (.A1_N(_03647_),
    .A2_N(_03648_),
    .B1(_03649_),
    .B2(_03650_),
    .X(_03651_));
 sky130_fd_sc_hd__a211o_2 _24295_ (.A1(_03646_),
    .A2(_03651_),
    .B1(_03450_),
    .C1(_03618_),
    .X(_03652_));
 sky130_fd_sc_hd__a21o_1 _24296_ (.A1(_03624_),
    .A2(_03625_),
    .B1(_03622_),
    .X(_03653_));
 sky130_fd_sc_hd__a211o_2 _24297_ (.A1(_03301_),
    .A2(_03653_),
    .B1(_03630_),
    .C1(_03620_),
    .X(_03654_));
 sky130_fd_sc_hd__a31o_1 _24298_ (.A1(_03624_),
    .A2(_03625_),
    .A3(_03622_),
    .B1(_03630_),
    .X(_03655_));
 sky130_fd_sc_hd__a31o_1 _24299_ (.A1(_03624_),
    .A2(_03625_),
    .A3(_03622_),
    .B1(_03620_),
    .X(_03656_));
 sky130_fd_sc_hd__a31o_2 _24300_ (.A1(_03653_),
    .A2(_03655_),
    .A3(_03656_),
    .B1(_03301_),
    .X(_03657_));
 sky130_fd_sc_hd__and3_1 _24301_ (.A(_03652_),
    .B(_03654_),
    .C(_03657_),
    .X(_03658_));
 sky130_fd_sc_hd__o211a_1 _24302_ (.A1(_03290_),
    .A2(_03287_),
    .B1(_03294_),
    .C1(_03293_),
    .X(_03659_));
 sky130_fd_sc_hd__a21o_1 _24303_ (.A1(_03290_),
    .A2(_03287_),
    .B1(_03659_),
    .X(_03660_));
 sky130_fd_sc_hd__a21bo_1 _24304_ (.A1(_03229_),
    .A2(_03230_),
    .B1_N(_03291_),
    .X(_03661_));
 sky130_fd_sc_hd__and3b_1 _24305_ (.A_N(_03291_),
    .B(_03229_),
    .C(_03230_),
    .X(_03662_));
 sky130_fd_sc_hd__a21oi_4 _24306_ (.A1(_03660_),
    .A2(_03661_),
    .B1(_03662_),
    .Y(_03663_));
 sky130_fd_sc_hd__nor2_1 _24307_ (.A(_03168_),
    .B(_03169_),
    .Y(_03664_));
 sky130_fd_sc_hd__and2_1 _24308_ (.A(_03130_),
    .B(_03135_),
    .X(_03665_));
 sky130_fd_sc_hd__and2_1 _24309_ (.A(_03225_),
    .B(_03226_),
    .X(_03666_));
 sky130_fd_sc_hd__o21a_1 _24310_ (.A1(_03110_),
    .A2(_03130_),
    .B1(_03135_),
    .X(_03667_));
 sky130_fd_sc_hd__a21bo_1 _24311_ (.A1(_03666_),
    .A2(_03667_),
    .B1_N(_03087_),
    .X(_03668_));
 sky130_fd_sc_hd__or2_1 _24312_ (.A(_03130_),
    .B(_03135_),
    .X(_03669_));
 sky130_fd_sc_hd__a31o_1 _24313_ (.A1(_03225_),
    .A2(_03226_),
    .A3(_03669_),
    .B1(_03110_),
    .X(_03670_));
 sky130_fd_sc_hd__o211a_1 _24314_ (.A1(_03665_),
    .A2(_03666_),
    .B1(_03668_),
    .C1(_03670_),
    .X(_03671_));
 sky130_fd_sc_hd__o21ai_1 _24315_ (.A1(_03110_),
    .A2(_03665_),
    .B1(_03669_),
    .Y(_03672_));
 sky130_fd_sc_hd__o2bb2a_1 _24316_ (.A1_N(_03087_),
    .A2_N(_03672_),
    .B1(_03669_),
    .B2(_03110_),
    .X(_03673_));
 sky130_fd_sc_hd__a21bo_1 _24317_ (.A1(_03132_),
    .A2(_03664_),
    .B1_N(_03133_),
    .X(_03674_));
 sky130_fd_sc_hd__mux2_1 _24318_ (.A0(_03673_),
    .A1(_03674_),
    .S(_03666_),
    .X(_03675_));
 sky130_fd_sc_hd__o21ai_4 _24319_ (.A1(_03664_),
    .A2(_03671_),
    .B1(_03675_),
    .Y(_03676_));
 sky130_fd_sc_hd__and2_1 _24320_ (.A(_03139_),
    .B(_03141_),
    .X(_03677_));
 sky130_fd_sc_hd__a21bo_1 _24321_ (.A1(_03677_),
    .A2(_03166_),
    .B1_N(_03154_),
    .X(_03678_));
 sky130_fd_sc_hd__o21ai_4 _24322_ (.A1(_03677_),
    .A2(_03166_),
    .B1(_03678_),
    .Y(_03679_));
 sky130_fd_sc_hd__nand2_2 _24323_ (.A(_03502_),
    .B(_03158_),
    .Y(_03680_));
 sky130_fd_sc_hd__o22a_2 _24324_ (.A1(_02985_),
    .A2(_02987_),
    .B1(_03024_),
    .B2(_03025_),
    .X(_03681_));
 sky130_fd_sc_hd__o22a_1 _24325_ (.A1(_02994_),
    .A2(_02996_),
    .B1(_02979_),
    .B2(_02980_),
    .X(_03682_));
 sky130_fd_sc_hd__xnor2_2 _24326_ (.A(_03681_),
    .B(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hd__xnor2_4 _24327_ (.A(_03680_),
    .B(_03683_),
    .Y(_03684_));
 sky130_fd_sc_hd__a21o_1 _24328_ (.A1(_03177_),
    .A2(_03179_),
    .B1(_03178_),
    .X(_03685_));
 sky130_fd_sc_hd__o21ai_2 _24329_ (.A1(_03177_),
    .A2(_03179_),
    .B1(_03685_),
    .Y(_03686_));
 sky130_fd_sc_hd__or2_2 _24330_ (.A(_03162_),
    .B(_03163_),
    .X(_03687_));
 sky130_fd_sc_hd__nand2_2 _24331_ (.A(_03572_),
    .B(_03687_),
    .Y(_03688_));
 sky130_fd_sc_hd__o22a_1 _24332_ (.A1(_03015_),
    .A2(_03016_),
    .B1(_03150_),
    .B2(_03151_),
    .X(_03689_));
 sky130_fd_sc_hd__o22a_1 _24333_ (.A1(_03045_),
    .A2(_03046_),
    .B1(_03029_),
    .B2(_03030_),
    .X(_03690_));
 sky130_fd_sc_hd__xnor2_2 _24334_ (.A(_03689_),
    .B(_03690_),
    .Y(_03691_));
 sky130_fd_sc_hd__xnor2_4 _24335_ (.A(_03688_),
    .B(_03691_),
    .Y(_03692_));
 sky130_fd_sc_hd__xnor2_2 _24336_ (.A(_03686_),
    .B(_03692_),
    .Y(_03693_));
 sky130_fd_sc_hd__xor2_4 _24337_ (.A(_03684_),
    .B(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__a21o_1 _24338_ (.A1(_03184_),
    .A2(_03190_),
    .B1(_03181_),
    .X(_03695_));
 sky130_fd_sc_hd__or2_1 _24339_ (.A(_03184_),
    .B(_03190_),
    .X(_03696_));
 sky130_fd_sc_hd__a21oi_2 _24340_ (.A1(_03213_),
    .A2(_03221_),
    .B1(_03220_),
    .Y(_03697_));
 sky130_fd_sc_hd__a21boi_1 _24341_ (.A1(_03695_),
    .A2(_03696_),
    .B1_N(_03697_),
    .Y(_03698_));
 sky130_fd_sc_hd__and3b_1 _24342_ (.A_N(_03697_),
    .B(_03695_),
    .C(_03696_),
    .X(_03699_));
 sky130_fd_sc_hd__nor2_1 _24343_ (.A(_03698_),
    .B(_03699_),
    .Y(_03700_));
 sky130_fd_sc_hd__xnor2_2 _24344_ (.A(_03694_),
    .B(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__and2_1 _24345_ (.A(_03206_),
    .B(_03223_),
    .X(_03702_));
 sky130_fd_sc_hd__nand2_1 _24346_ (.A(_03202_),
    .B(_03203_),
    .Y(_03703_));
 sky130_fd_sc_hd__o211ai_2 _24347_ (.A1(_03202_),
    .A2(_03203_),
    .B1(_03060_),
    .C1(_03124_),
    .Y(_03704_));
 sky130_fd_sc_hd__a21oi_1 _24348_ (.A1(_03210_),
    .A2(_03211_),
    .B1(_03209_),
    .Y(_03705_));
 sky130_fd_sc_hd__nor2_1 _24349_ (.A(_03210_),
    .B(_03211_),
    .Y(_03706_));
 sky130_fd_sc_hd__a211oi_1 _24350_ (.A1(_03703_),
    .A2(_03704_),
    .B1(_03705_),
    .C1(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__o211a_1 _24351_ (.A1(_03705_),
    .A2(_03706_),
    .B1(_03703_),
    .C1(_03704_),
    .X(_03708_));
 sky130_fd_sc_hd__o22a_1 _24352_ (.A1(_02989_),
    .A2(_02991_),
    .B1(_03054_),
    .B2(_03055_),
    .X(_03709_));
 sky130_fd_sc_hd__o22a_1 _24353_ (.A1(_02998_),
    .A2(_03000_),
    .B1(_03069_),
    .B2(_03071_),
    .X(_03710_));
 sky130_fd_sc_hd__o22a_1 _24354_ (.A1(_03004_),
    .A2(_03005_),
    .B1(_03061_),
    .B2(_03062_),
    .X(_03711_));
 sky130_fd_sc_hd__xor2_1 _24355_ (.A(_03710_),
    .B(_03711_),
    .X(_03712_));
 sky130_fd_sc_hd__xnor2_2 _24356_ (.A(_03709_),
    .B(_03712_),
    .Y(_03713_));
 sky130_fd_sc_hd__o21ai_1 _24357_ (.A1(_03707_),
    .A2(_03708_),
    .B1(_03713_),
    .Y(_03714_));
 sky130_fd_sc_hd__or3_1 _24358_ (.A(_03713_),
    .B(_03707_),
    .C(_03708_),
    .X(_03715_));
 sky130_fd_sc_hd__and2_1 _24359_ (.A(_03714_),
    .B(_03715_),
    .X(_03716_));
 sky130_fd_sc_hd__o21a_2 _24360_ (.A1(net571),
    .A2(net575),
    .B1(\top0.matmul0.matmul_stage_inst.f[14] ),
    .X(_03717_));
 sky130_fd_sc_hd__o21a_2 _24361_ (.A1(net566),
    .A2(net560),
    .B1(\top0.matmul0.matmul_stage_inst.e[14] ),
    .X(_03718_));
 sky130_fd_sc_hd__nor2_2 _24362_ (.A(_03717_),
    .B(_03718_),
    .Y(_03719_));
 sky130_fd_sc_hd__or2_2 _24363_ (.A(_03196_),
    .B(_03197_),
    .X(_03720_));
 sky130_fd_sc_hd__o211a_1 _24364_ (.A1(_03195_),
    .A2(_03719_),
    .B1(_03720_),
    .C1(_03324_),
    .X(_03721_));
 sky130_fd_sc_hd__or2_2 _24365_ (.A(_03717_),
    .B(_03718_),
    .X(_03722_));
 sky130_fd_sc_hd__o211a_1 _24366_ (.A1(_03252_),
    .A2(_03198_),
    .B1(_03722_),
    .C1(_03120_),
    .X(_03723_));
 sky130_fd_sc_hd__nor2_1 _24367_ (.A(_03721_),
    .B(_03723_),
    .Y(_03724_));
 sky130_fd_sc_hd__nand2_1 _24368_ (.A(_03060_),
    .B(_03123_),
    .Y(_03725_));
 sky130_fd_sc_hd__o22a_1 _24369_ (.A1(_03076_),
    .A2(_03077_),
    .B1(_03103_),
    .B2(_03104_),
    .X(_03726_));
 sky130_fd_sc_hd__o22a_1 _24370_ (.A1(_03207_),
    .A2(_03208_),
    .B1(_03093_),
    .B2(_03094_),
    .X(_03727_));
 sky130_fd_sc_hd__xnor2_1 _24371_ (.A(_03726_),
    .B(_03727_),
    .Y(_03728_));
 sky130_fd_sc_hd__xnor2_2 _24372_ (.A(_03725_),
    .B(_03728_),
    .Y(_03729_));
 sky130_fd_sc_hd__xnor2_2 _24373_ (.A(_03724_),
    .B(_03729_),
    .Y(_03730_));
 sky130_fd_sc_hd__nand2_1 _24374_ (.A(_03199_),
    .B(_03205_),
    .Y(_03731_));
 sky130_fd_sc_hd__xor2_2 _24375_ (.A(_03730_),
    .B(_03731_),
    .X(_03732_));
 sky130_fd_sc_hd__xor2_2 _24376_ (.A(_03716_),
    .B(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__xnor2_1 _24377_ (.A(_03702_),
    .B(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__xnor2_2 _24378_ (.A(_03701_),
    .B(_03734_),
    .Y(_03735_));
 sky130_fd_sc_hd__a21boi_2 _24379_ (.A1(_03133_),
    .A2(_03226_),
    .B1_N(_03225_),
    .Y(_03736_));
 sky130_fd_sc_hd__o2bb2a_1 _24380_ (.A1_N(_03170_),
    .A2_N(_03171_),
    .B1(_03192_),
    .B2(_03174_),
    .X(_03737_));
 sky130_fd_sc_hd__a21o_2 _24381_ (.A1(_03192_),
    .A2(_03174_),
    .B1(_03737_),
    .X(_03738_));
 sky130_fd_sc_hd__a21oi_1 _24382_ (.A1(_03186_),
    .A2(_03187_),
    .B1(_03188_),
    .Y(_03739_));
 sky130_fd_sc_hd__o21ba_1 _24383_ (.A1(_03186_),
    .A2(_03187_),
    .B1_N(_03739_),
    .X(_03740_));
 sky130_fd_sc_hd__o21a_4 _24384_ (.A1(net573),
    .A2(net564),
    .B1(\top0.matmul0.matmul_stage_inst.a[14] ),
    .X(_03741_));
 sky130_fd_sc_hd__a22o_4 _24385_ (.A1(net556),
    .A2(\top0.matmul0.matmul_stage_inst.c[14] ),
    .B1(\top0.matmul0.matmul_stage_inst.b[14] ),
    .B2(net568),
    .X(_03742_));
 sky130_fd_sc_hd__nor2_2 _24386_ (.A(_03741_),
    .B(_03742_),
    .Y(_03743_));
 sky130_fd_sc_hd__nor2_1 _24387_ (.A(_03161_),
    .B(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__xor2_2 _24388_ (.A(_03740_),
    .B(_03744_),
    .X(_03745_));
 sky130_fd_sc_hd__and2_1 _24389_ (.A(_03160_),
    .B(_03165_),
    .X(_03746_));
 sky130_fd_sc_hd__xnor2_1 _24390_ (.A(_03745_),
    .B(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__xnor2_2 _24391_ (.A(_03738_),
    .B(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__xor2_1 _24392_ (.A(_03736_),
    .B(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__xnor2_1 _24393_ (.A(_03735_),
    .B(_03749_),
    .Y(_03750_));
 sky130_fd_sc_hd__nand2_2 _24394_ (.A(_03679_),
    .B(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__or2_1 _24395_ (.A(_03679_),
    .B(_03750_),
    .X(_03752_));
 sky130_fd_sc_hd__nand2_1 _24396_ (.A(_03751_),
    .B(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__xor2_1 _24397_ (.A(_03676_),
    .B(_03753_),
    .X(_03754_));
 sky130_fd_sc_hd__xnor2_1 _24398_ (.A(_03663_),
    .B(_03754_),
    .Y(_03755_));
 sky130_fd_sc_hd__xnor2_1 _24399_ (.A(_03658_),
    .B(_03755_),
    .Y(_03756_));
 sky130_fd_sc_hd__mux2_1 _24400_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[1] ),
    .A1(_03756_),
    .S(_03642_),
    .X(_03757_));
 sky130_fd_sc_hd__clkbuf_1 _24401_ (.A(_03757_),
    .X(_00602_));
 sky130_fd_sc_hd__or2_2 _24402_ (.A(_03029_),
    .B(_03030_),
    .X(_03758_));
 sky130_fd_sc_hd__nand2_1 _24403_ (.A(_03502_),
    .B(_03758_),
    .Y(_03759_));
 sky130_fd_sc_hd__o22a_1 _24404_ (.A1(_02985_),
    .A2(_02987_),
    .B1(_03018_),
    .B2(_03019_),
    .X(_03760_));
 sky130_fd_sc_hd__o22a_1 _24405_ (.A1(_02994_),
    .A2(_02996_),
    .B1(_03024_),
    .B2(_03025_),
    .X(_03761_));
 sky130_fd_sc_hd__xnor2_1 _24406_ (.A(_03760_),
    .B(_03761_),
    .Y(_03762_));
 sky130_fd_sc_hd__xnor2_2 _24407_ (.A(_03759_),
    .B(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__a21oi_1 _24408_ (.A1(_03502_),
    .A2(_03158_),
    .B1(_03681_),
    .Y(_03764_));
 sky130_fd_sc_hd__clkbuf_4 _24409_ (.A(_02978_),
    .X(_03765_));
 sky130_fd_sc_hd__or3b_1 _24410_ (.A(_03765_),
    .B(net1017),
    .C_N(_03681_),
    .X(_03766_));
 sky130_fd_sc_hd__o31a_1 _24411_ (.A1(_03007_),
    .A2(_02982_),
    .A3(_03764_),
    .B1(_03766_),
    .X(_03767_));
 sky130_fd_sc_hd__nor2_2 _24412_ (.A(_03185_),
    .B(_03743_),
    .Y(_03768_));
 sky130_fd_sc_hd__o22a_1 _24413_ (.A1(_03015_),
    .A2(_03016_),
    .B1(_03162_),
    .B2(_03163_),
    .X(_03769_));
 sky130_fd_sc_hd__o22a_1 _24414_ (.A1(_03045_),
    .A2(_03046_),
    .B1(_03150_),
    .B2(_03151_),
    .X(_03770_));
 sky130_fd_sc_hd__xor2_1 _24415_ (.A(_03769_),
    .B(_03770_),
    .X(_03771_));
 sky130_fd_sc_hd__xnor2_2 _24416_ (.A(_03768_),
    .B(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__xnor2_1 _24417_ (.A(_03767_),
    .B(_03772_),
    .Y(_03773_));
 sky130_fd_sc_hd__xnor2_2 _24418_ (.A(_03763_),
    .B(_03773_),
    .Y(_03774_));
 sky130_fd_sc_hd__or2_1 _24419_ (.A(_03686_),
    .B(_03692_),
    .X(_03775_));
 sky130_fd_sc_hd__a21o_1 _24420_ (.A1(_03686_),
    .A2(_03692_),
    .B1(_03684_),
    .X(_03776_));
 sky130_fd_sc_hd__nand2_1 _24421_ (.A(_03775_),
    .B(_03776_),
    .Y(_03777_));
 sky130_fd_sc_hd__a211o_1 _24422_ (.A1(_03703_),
    .A2(_03704_),
    .B1(_03705_),
    .C1(_03706_),
    .X(_03778_));
 sky130_fd_sc_hd__o21ai_1 _24423_ (.A1(_03713_),
    .A2(_03708_),
    .B1(_03778_),
    .Y(_03779_));
 sky130_fd_sc_hd__xor2_1 _24424_ (.A(_03777_),
    .B(_03779_),
    .X(_03780_));
 sky130_fd_sc_hd__xnor2_2 _24425_ (.A(_03774_),
    .B(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__nor2_1 _24426_ (.A(_03730_),
    .B(_03731_),
    .Y(_03782_));
 sky130_fd_sc_hd__a21o_1 _24427_ (.A1(_03716_),
    .A2(_03732_),
    .B1(_03782_),
    .X(_03783_));
 sky130_fd_sc_hd__and2_1 _24428_ (.A(_03726_),
    .B(_03727_),
    .X(_03784_));
 sky130_fd_sc_hd__o211a_1 _24429_ (.A1(_03726_),
    .A2(_03727_),
    .B1(_03060_),
    .C1(_03123_),
    .X(_03785_));
 sky130_fd_sc_hd__a21o_1 _24430_ (.A1(_03709_),
    .A2(_03710_),
    .B1(_03711_),
    .X(_03786_));
 sky130_fd_sc_hd__or2_1 _24431_ (.A(_03709_),
    .B(_03710_),
    .X(_03787_));
 sky130_fd_sc_hd__o211a_1 _24432_ (.A1(_03784_),
    .A2(_03785_),
    .B1(_03786_),
    .C1(_03787_),
    .X(_03788_));
 sky130_fd_sc_hd__a211oi_2 _24433_ (.A1(_03786_),
    .A2(_03787_),
    .B1(_03784_),
    .C1(_03785_),
    .Y(_03789_));
 sky130_fd_sc_hd__o22a_1 _24434_ (.A1(_02989_),
    .A2(_02991_),
    .B1(_03069_),
    .B2(_03071_),
    .X(_03790_));
 sky130_fd_sc_hd__o22a_1 _24435_ (.A1(_02998_),
    .A2(_03000_),
    .B1(_03061_),
    .B2(_03062_),
    .X(_03791_));
 sky130_fd_sc_hd__o22a_1 _24436_ (.A1(_02979_),
    .A2(_02980_),
    .B1(_03054_),
    .B2(_03055_),
    .X(_03792_));
 sky130_fd_sc_hd__xor2_1 _24437_ (.A(_03791_),
    .B(_03792_),
    .X(_03793_));
 sky130_fd_sc_hd__xnor2_1 _24438_ (.A(_03790_),
    .B(_03793_),
    .Y(_03794_));
 sky130_fd_sc_hd__o21ai_1 _24439_ (.A1(_03788_),
    .A2(_03789_),
    .B1(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__or3_1 _24440_ (.A(_03794_),
    .B(_03788_),
    .C(_03789_),
    .X(_03796_));
 sky130_fd_sc_hd__and2_1 _24441_ (.A(_03795_),
    .B(_03796_),
    .X(_03797_));
 sky130_fd_sc_hd__nor2_1 _24442_ (.A(_03724_),
    .B(_03729_),
    .Y(_03798_));
 sky130_fd_sc_hd__nor2_1 _24443_ (.A(_03103_),
    .B(_03104_),
    .Y(_03799_));
 sky130_fd_sc_hd__nor2_1 _24444_ (.A(_03114_),
    .B(_03799_),
    .Y(_03800_));
 sky130_fd_sc_hd__o22a_1 _24445_ (.A1(_03207_),
    .A2(_03208_),
    .B1(_03090_),
    .B2(_03091_),
    .X(_03801_));
 sky130_fd_sc_hd__o22a_1 _24446_ (.A1(_03004_),
    .A2(_03005_),
    .B1(_03093_),
    .B2(_03094_),
    .X(_03802_));
 sky130_fd_sc_hd__xnor2_1 _24447_ (.A(_03801_),
    .B(_03802_),
    .Y(_03803_));
 sky130_fd_sc_hd__xnor2_2 _24448_ (.A(_03800_),
    .B(_03803_),
    .Y(_03804_));
 sky130_fd_sc_hd__o21ai_2 _24449_ (.A1(net570),
    .A2(net574),
    .B1(\top0.matmul0.matmul_stage_inst.f[15] ),
    .Y(_03805_));
 sky130_fd_sc_hd__o21ai_2 _24450_ (.A1(net566),
    .A2(net558),
    .B1(\top0.matmul0.matmul_stage_inst.e[15] ),
    .Y(_03806_));
 sky130_fd_sc_hd__a211o_2 _24451_ (.A1(_03805_),
    .A2(_03806_),
    .B1(_03088_),
    .C1(_03089_),
    .X(_03807_));
 sky130_fd_sc_hd__o22a_1 _24452_ (.A1(_03076_),
    .A2(_03077_),
    .B1(_03196_),
    .B2(_03197_),
    .X(_03808_));
 sky130_fd_sc_hd__xnor2_2 _24453_ (.A(_03807_),
    .B(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__o211a_1 _24454_ (.A1(_03195_),
    .A2(_03198_),
    .B1(_03722_),
    .C1(_03324_),
    .X(_03810_));
 sky130_fd_sc_hd__xnor2_1 _24455_ (.A(_03809_),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__xnor2_2 _24456_ (.A(_03804_),
    .B(_03811_),
    .Y(_03812_));
 sky130_fd_sc_hd__xnor2_1 _24457_ (.A(_03798_),
    .B(_03812_),
    .Y(_03813_));
 sky130_fd_sc_hd__xnor2_2 _24458_ (.A(_03797_),
    .B(_03813_),
    .Y(_03814_));
 sky130_fd_sc_hd__xor2_1 _24459_ (.A(_03783_),
    .B(_03814_),
    .X(_03815_));
 sky130_fd_sc_hd__xnor2_2 _24460_ (.A(_03781_),
    .B(_03815_),
    .Y(_03816_));
 sky130_fd_sc_hd__a21bo_1 _24461_ (.A1(_03206_),
    .A2(_03223_),
    .B1_N(_03694_),
    .X(_03817_));
 sky130_fd_sc_hd__a2111o_1 _24462_ (.A1(_03206_),
    .A2(_03223_),
    .B1(_03694_),
    .C1(_03698_),
    .D1(_03699_),
    .X(_03818_));
 sky130_fd_sc_hd__o221a_1 _24463_ (.A1(_03702_),
    .A2(_03733_),
    .B1(_03817_),
    .B2(_03700_),
    .C1(_03818_),
    .X(_03819_));
 sky130_fd_sc_hd__o21ai_2 _24464_ (.A1(_03701_),
    .A2(_03733_),
    .B1(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hd__nand2_1 _24465_ (.A(_03740_),
    .B(_03744_),
    .Y(_03821_));
 sky130_fd_sc_hd__a21o_1 _24466_ (.A1(_03572_),
    .A2(_03687_),
    .B1(_03689_),
    .X(_03822_));
 sky130_fd_sc_hd__and3_1 _24467_ (.A(_03572_),
    .B(_03687_),
    .C(_03689_),
    .X(_03823_));
 sky130_fd_sc_hd__a21o_1 _24468_ (.A1(_03690_),
    .A2(_03822_),
    .B1(_03823_),
    .X(_03824_));
 sky130_fd_sc_hd__nand2_2 _24469_ (.A(_03805_),
    .B(_03806_),
    .Y(_03825_));
 sky130_fd_sc_hd__clkbuf_4 _24470_ (.A(_03825_),
    .X(_03826_));
 sky130_fd_sc_hd__a22o_2 _24471_ (.A1(net556),
    .A2(\top0.matmul0.matmul_stage_inst.c[15] ),
    .B1(\top0.matmul0.matmul_stage_inst.b[15] ),
    .B2(net568),
    .X(_03827_));
 sky130_fd_sc_hd__or2_1 _24472_ (.A(_03741_),
    .B(_03827_),
    .X(_03828_));
 sky130_fd_sc_hd__clkbuf_4 _24473_ (.A(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__nand2_2 _24474_ (.A(_03549_),
    .B(_03829_),
    .Y(_03830_));
 sky130_fd_sc_hd__xnor2_1 _24475_ (.A(_03826_),
    .B(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__xnor2_1 _24476_ (.A(_03824_),
    .B(_03831_),
    .Y(_03832_));
 sky130_fd_sc_hd__or2_1 _24477_ (.A(_03821_),
    .B(_03832_),
    .X(_03833_));
 sky130_fd_sc_hd__nand2_1 _24478_ (.A(_03821_),
    .B(_03832_),
    .Y(_03834_));
 sky130_fd_sc_hd__nand2_1 _24479_ (.A(_03833_),
    .B(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__a22o_1 _24480_ (.A1(_03694_),
    .A2(_03697_),
    .B1(_03695_),
    .B2(_03696_),
    .X(_03836_));
 sky130_fd_sc_hd__o21ai_4 _24481_ (.A1(_03694_),
    .A2(_03697_),
    .B1(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__xnor2_2 _24482_ (.A(_03835_),
    .B(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__xnor2_1 _24483_ (.A(_03820_),
    .B(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__xnor2_2 _24484_ (.A(_03816_),
    .B(_03839_),
    .Y(_03840_));
 sky130_fd_sc_hd__o21bai_1 _24485_ (.A1(_03735_),
    .A2(_03748_),
    .B1_N(_03736_),
    .Y(_03841_));
 sky130_fd_sc_hd__a21bo_1 _24486_ (.A1(_03735_),
    .A2(_03748_),
    .B1_N(_03841_),
    .X(_03842_));
 sky130_fd_sc_hd__a21o_1 _24487_ (.A1(_03738_),
    .A2(_03745_),
    .B1(_03746_),
    .X(_03843_));
 sky130_fd_sc_hd__o21a_1 _24488_ (.A1(_03738_),
    .A2(_03745_),
    .B1(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__xnor2_1 _24489_ (.A(_03842_),
    .B(_03844_),
    .Y(_03845_));
 sky130_fd_sc_hd__xnor2_2 _24490_ (.A(_03840_),
    .B(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__or2_1 _24491_ (.A(_03663_),
    .B(_03676_),
    .X(_03847_));
 sky130_fd_sc_hd__nand2_1 _24492_ (.A(_03663_),
    .B(_03676_),
    .Y(_03848_));
 sky130_fd_sc_hd__inv_2 _24493_ (.A(_03752_),
    .Y(_03849_));
 sky130_fd_sc_hd__o21a_1 _24494_ (.A1(_03663_),
    .A2(_03849_),
    .B1(_03751_),
    .X(_03850_));
 sky130_fd_sc_hd__o22a_1 _24495_ (.A1(_03663_),
    .A2(_03751_),
    .B1(_03850_),
    .B2(_03676_),
    .X(_03851_));
 sky130_fd_sc_hd__a22oi_1 _24496_ (.A1(_03663_),
    .A2(_03849_),
    .B1(_03850_),
    .B2(_03676_),
    .Y(_03852_));
 sky130_fd_sc_hd__mux2_1 _24497_ (.A0(_03851_),
    .A1(_03852_),
    .S(_03658_),
    .X(_03853_));
 sky130_fd_sc_hd__o221a_1 _24498_ (.A1(_03751_),
    .A2(_03847_),
    .B1(_03848_),
    .B2(_03752_),
    .C1(_03853_),
    .X(_03854_));
 sky130_fd_sc_hd__xnor2_1 _24499_ (.A(_03846_),
    .B(_03854_),
    .Y(_03855_));
 sky130_fd_sc_hd__mux2_1 _24500_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[2] ),
    .A1(_03855_),
    .S(_03642_),
    .X(_03856_));
 sky130_fd_sc_hd__clkbuf_1 _24501_ (.A(_03856_),
    .X(_00603_));
 sky130_fd_sc_hd__and3_1 _24502_ (.A(_03654_),
    .B(_03657_),
    .C(_03847_),
    .X(_03857_));
 sky130_fd_sc_hd__and2_1 _24503_ (.A(_03663_),
    .B(_03676_),
    .X(_03858_));
 sky130_fd_sc_hd__a221oi_1 _24504_ (.A1(_03751_),
    .A2(_03846_),
    .B1(_03857_),
    .B2(_03652_),
    .C1(_03858_),
    .Y(_03859_));
 sky130_fd_sc_hd__nor2_1 _24505_ (.A(_03751_),
    .B(_03846_),
    .Y(_03860_));
 sky130_fd_sc_hd__o211a_1 _24506_ (.A1(_03846_),
    .A2(_03858_),
    .B1(_03654_),
    .C1(_03657_),
    .X(_03861_));
 sky130_fd_sc_hd__a221oi_1 _24507_ (.A1(_03846_),
    .A2(_03847_),
    .B1(_03861_),
    .B2(_03652_),
    .C1(_03849_),
    .Y(_03862_));
 sky130_fd_sc_hd__or3_2 _24508_ (.A(_03859_),
    .B(_03860_),
    .C(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__o22a_2 _24509_ (.A1(_03207_),
    .A2(_03208_),
    .B1(_03103_),
    .B2(_03104_),
    .X(_03864_));
 sky130_fd_sc_hd__o22a_2 _24510_ (.A1(_02998_),
    .A2(_03000_),
    .B1(_03093_),
    .B2(_03094_),
    .X(_03865_));
 sky130_fd_sc_hd__o22a_1 _24511_ (.A1(_03004_),
    .A2(_03005_),
    .B1(_03090_),
    .B2(_03091_),
    .X(_03866_));
 sky130_fd_sc_hd__xor2_2 _24512_ (.A(_03865_),
    .B(_03866_),
    .X(_03867_));
 sky130_fd_sc_hd__xnor2_4 _24513_ (.A(_03864_),
    .B(_03867_),
    .Y(_03868_));
 sky130_fd_sc_hd__nor2_1 _24514_ (.A(_03252_),
    .B(_03719_),
    .Y(_03869_));
 sky130_fd_sc_hd__and3_1 _24515_ (.A(_03195_),
    .B(_03825_),
    .C(_03808_),
    .X(_03870_));
 sky130_fd_sc_hd__o21ai_1 _24516_ (.A1(_03106_),
    .A2(_03198_),
    .B1(_03807_),
    .Y(_03871_));
 sky130_fd_sc_hd__o21a_1 _24517_ (.A1(_03869_),
    .A2(_03870_),
    .B1(_03871_),
    .X(_03872_));
 sky130_fd_sc_hd__nand2_1 _24518_ (.A(_03252_),
    .B(_03825_),
    .Y(_03873_));
 sky130_fd_sc_hd__o22a_1 _24519_ (.A1(_03057_),
    .A2(_03058_),
    .B1(_03196_),
    .B2(_03197_),
    .X(_03874_));
 sky130_fd_sc_hd__o22a_1 _24520_ (.A1(_03076_),
    .A2(_03077_),
    .B1(_03717_),
    .B2(_03718_),
    .X(_03875_));
 sky130_fd_sc_hd__xnor2_1 _24521_ (.A(_03874_),
    .B(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hd__xnor2_2 _24522_ (.A(_03873_),
    .B(_03876_),
    .Y(_03877_));
 sky130_fd_sc_hd__xnor2_2 _24523_ (.A(_03872_),
    .B(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__xnor2_4 _24524_ (.A(_03868_),
    .B(_03878_),
    .Y(_03879_));
 sky130_fd_sc_hd__a21boi_1 _24525_ (.A1(_03809_),
    .A2(_03869_),
    .B1_N(_03804_),
    .Y(_03880_));
 sky130_fd_sc_hd__mux2_1 _24526_ (.A0(_03869_),
    .A1(_03804_),
    .S(_03809_),
    .X(_03881_));
 sky130_fd_sc_hd__o21ai_4 _24527_ (.A1(_03199_),
    .A2(_03880_),
    .B1(_03881_),
    .Y(_03882_));
 sky130_fd_sc_hd__o22a_2 _24528_ (.A1(_03024_),
    .A2(_03025_),
    .B1(_03054_),
    .B2(_03055_),
    .X(_03883_));
 sky130_fd_sc_hd__o22a_2 _24529_ (.A1(_02979_),
    .A2(_02980_),
    .B1(_03069_),
    .B2(_03071_),
    .X(_03884_));
 sky130_fd_sc_hd__o22a_1 _24530_ (.A1(_02989_),
    .A2(_02991_),
    .B1(_03061_),
    .B2(_03062_),
    .X(_03885_));
 sky130_fd_sc_hd__xnor2_1 _24531_ (.A(_03884_),
    .B(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__xnor2_2 _24532_ (.A(_03883_),
    .B(_03886_),
    .Y(_03887_));
 sky130_fd_sc_hd__or2_1 _24533_ (.A(_03103_),
    .B(_03104_),
    .X(_03888_));
 sky130_fd_sc_hd__clkbuf_4 _24534_ (.A(_03888_),
    .X(_03889_));
 sky130_fd_sc_hd__a22o_1 _24535_ (.A1(_03060_),
    .A2(_03889_),
    .B1(_03801_),
    .B2(_03802_),
    .X(_03890_));
 sky130_fd_sc_hd__or2_1 _24536_ (.A(_03801_),
    .B(_03802_),
    .X(_03891_));
 sky130_fd_sc_hd__and2_1 _24537_ (.A(_03790_),
    .B(_03792_),
    .X(_03892_));
 sky130_fd_sc_hd__o21a_1 _24538_ (.A1(_03790_),
    .A2(_03792_),
    .B1(_03791_),
    .X(_03893_));
 sky130_fd_sc_hd__a211oi_1 _24539_ (.A1(_03890_),
    .A2(_03891_),
    .B1(_03892_),
    .C1(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__o211a_1 _24540_ (.A1(_03892_),
    .A2(_03893_),
    .B1(_03890_),
    .C1(_03891_),
    .X(_03895_));
 sky130_fd_sc_hd__nor2_1 _24541_ (.A(_03894_),
    .B(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__xnor2_2 _24542_ (.A(_03887_),
    .B(_03896_),
    .Y(_03897_));
 sky130_fd_sc_hd__xor2_2 _24543_ (.A(_03882_),
    .B(_03897_),
    .X(_03898_));
 sky130_fd_sc_hd__xnor2_4 _24544_ (.A(_03879_),
    .B(_03898_),
    .Y(_03899_));
 sky130_fd_sc_hd__buf_4 _24545_ (.A(_03152_),
    .X(_03900_));
 sky130_fd_sc_hd__nor2_1 _24546_ (.A(_03765_),
    .B(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__o22a_1 _24547_ (.A1(_02985_),
    .A2(_02987_),
    .B1(_03029_),
    .B2(_03030_),
    .X(_03902_));
 sky130_fd_sc_hd__o22a_1 _24548_ (.A1(_02994_),
    .A2(_02996_),
    .B1(_03018_),
    .B2(_03019_),
    .X(_03903_));
 sky130_fd_sc_hd__xnor2_1 _24549_ (.A(_03902_),
    .B(_03903_),
    .Y(_03904_));
 sky130_fd_sc_hd__xnor2_2 _24550_ (.A(_03901_),
    .B(_03904_),
    .Y(_03905_));
 sky130_fd_sc_hd__a22o_1 _24551_ (.A1(_03502_),
    .A2(_03758_),
    .B1(_03760_),
    .B2(_03761_),
    .X(_03906_));
 sky130_fd_sc_hd__o21a_1 _24552_ (.A1(_03760_),
    .A2(_03761_),
    .B1(_03906_),
    .X(_03907_));
 sky130_fd_sc_hd__nor2_2 _24553_ (.A(_03741_),
    .B(_03827_),
    .Y(_03908_));
 sky130_fd_sc_hd__nor2_1 _24554_ (.A(_03185_),
    .B(_03908_),
    .Y(_03909_));
 sky130_fd_sc_hd__o22a_1 _24555_ (.A1(_03015_),
    .A2(_03016_),
    .B1(_03741_),
    .B2(_03742_),
    .X(_03910_));
 sky130_fd_sc_hd__o22a_1 _24556_ (.A1(_03045_),
    .A2(_03046_),
    .B1(_03162_),
    .B2(_03163_),
    .X(_03911_));
 sky130_fd_sc_hd__xnor2_1 _24557_ (.A(_03910_),
    .B(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__xnor2_2 _24558_ (.A(_03909_),
    .B(_03912_),
    .Y(_03913_));
 sky130_fd_sc_hd__xnor2_1 _24559_ (.A(_03907_),
    .B(_03913_),
    .Y(_03914_));
 sky130_fd_sc_hd__xnor2_2 _24560_ (.A(_03905_),
    .B(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__or2_1 _24561_ (.A(_03767_),
    .B(_03772_),
    .X(_03916_));
 sky130_fd_sc_hd__a21o_1 _24562_ (.A1(_03767_),
    .A2(_03772_),
    .B1(_03763_),
    .X(_03917_));
 sky130_fd_sc_hd__o21bai_2 _24563_ (.A1(_03794_),
    .A2(_03789_),
    .B1_N(_03788_),
    .Y(_03918_));
 sky130_fd_sc_hd__a21oi_1 _24564_ (.A1(_03916_),
    .A2(_03917_),
    .B1(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__and3_1 _24565_ (.A(_03916_),
    .B(_03917_),
    .C(_03918_),
    .X(_03920_));
 sky130_fd_sc_hd__or3_2 _24566_ (.A(_03915_),
    .B(_03919_),
    .C(_03920_),
    .X(_03921_));
 sky130_fd_sc_hd__o21ai_2 _24567_ (.A1(_03919_),
    .A2(_03920_),
    .B1(_03915_),
    .Y(_03922_));
 sky130_fd_sc_hd__a31o_1 _24568_ (.A1(_03795_),
    .A2(_03796_),
    .A3(_03812_),
    .B1(_03798_),
    .X(_03923_));
 sky130_fd_sc_hd__o21ai_2 _24569_ (.A1(_03797_),
    .A2(_03812_),
    .B1(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__a21oi_1 _24570_ (.A1(_03921_),
    .A2(_03922_),
    .B1(_03924_),
    .Y(_03925_));
 sky130_fd_sc_hd__and3_1 _24571_ (.A(_03924_),
    .B(_03921_),
    .C(_03922_),
    .X(_03926_));
 sky130_fd_sc_hd__or2_1 _24572_ (.A(_03925_),
    .B(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__xnor2_2 _24573_ (.A(_03899_),
    .B(_03927_),
    .Y(_03928_));
 sky130_fd_sc_hd__and2_1 _24574_ (.A(_03783_),
    .B(_03814_),
    .X(_03929_));
 sky130_fd_sc_hd__nor2_1 _24575_ (.A(_03783_),
    .B(_03814_),
    .Y(_03930_));
 sky130_fd_sc_hd__o21bai_2 _24576_ (.A1(_03781_),
    .A2(_03929_),
    .B1_N(_03930_),
    .Y(_03931_));
 sky130_fd_sc_hd__a21bo_1 _24577_ (.A1(_03775_),
    .A2(_03776_),
    .B1_N(_03779_),
    .X(_03932_));
 sky130_fd_sc_hd__o2111a_1 _24578_ (.A1(_03713_),
    .A2(_03708_),
    .B1(_03775_),
    .C1(_03776_),
    .D1(_03778_),
    .X(_03933_));
 sky130_fd_sc_hd__a21o_1 _24579_ (.A1(_03774_),
    .A2(_03932_),
    .B1(_03933_),
    .X(_03934_));
 sky130_fd_sc_hd__nor2_1 _24580_ (.A(_03161_),
    .B(_03908_),
    .Y(_03935_));
 sky130_fd_sc_hd__clkbuf_4 _24581_ (.A(_03826_),
    .X(_03936_));
 sky130_fd_sc_hd__o21ai_1 _24582_ (.A1(_03824_),
    .A2(_03935_),
    .B1(_03936_),
    .Y(_03937_));
 sky130_fd_sc_hd__nand2_1 _24583_ (.A(_03824_),
    .B(_03935_),
    .Y(_03938_));
 sky130_fd_sc_hd__nand2_1 _24584_ (.A(_03937_),
    .B(_03938_),
    .Y(_03939_));
 sky130_fd_sc_hd__o21ai_2 _24585_ (.A1(_03768_),
    .A2(_03769_),
    .B1(_03770_),
    .Y(_03940_));
 sky130_fd_sc_hd__nand2_1 _24586_ (.A(_03768_),
    .B(_03769_),
    .Y(_03941_));
 sky130_fd_sc_hd__a21oi_2 _24587_ (.A1(_03940_),
    .A2(_03941_),
    .B1(_03830_),
    .Y(_03942_));
 sky130_fd_sc_hd__and3_1 _24588_ (.A(_03830_),
    .B(_03940_),
    .C(_03941_),
    .X(_03943_));
 sky130_fd_sc_hd__or2_1 _24589_ (.A(_03942_),
    .B(_03943_),
    .X(_03944_));
 sky130_fd_sc_hd__xnor2_1 _24590_ (.A(_03939_),
    .B(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__xnor2_2 _24591_ (.A(_03934_),
    .B(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__xnor2_1 _24592_ (.A(_03931_),
    .B(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__xnor2_2 _24593_ (.A(_03928_),
    .B(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__a21o_1 _24594_ (.A1(_03820_),
    .A2(_03838_),
    .B1(_03816_),
    .X(_03949_));
 sky130_fd_sc_hd__o21ai_2 _24595_ (.A1(_03820_),
    .A2(_03838_),
    .B1(_03949_),
    .Y(_03950_));
 sky130_fd_sc_hd__nand2_1 _24596_ (.A(_03833_),
    .B(_03837_),
    .Y(_03951_));
 sky130_fd_sc_hd__nand2_1 _24597_ (.A(_03834_),
    .B(_03951_),
    .Y(_03952_));
 sky130_fd_sc_hd__xor2_1 _24598_ (.A(_03950_),
    .B(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__xnor2_1 _24599_ (.A(_03948_),
    .B(_03953_),
    .Y(_03954_));
 sky130_fd_sc_hd__a21bo_1 _24600_ (.A1(_03842_),
    .A2(_03844_),
    .B1_N(_03840_),
    .X(_03955_));
 sky130_fd_sc_hd__o21ai_2 _24601_ (.A1(_03842_),
    .A2(_03844_),
    .B1(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__nand2_1 _24602_ (.A(_03954_),
    .B(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hd__or2_1 _24603_ (.A(_03954_),
    .B(_03956_),
    .X(_03958_));
 sky130_fd_sc_hd__nand2_1 _24604_ (.A(_03957_),
    .B(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__xnor2_1 _24605_ (.A(_03863_),
    .B(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__mux2_1 _24606_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[3] ),
    .A1(_03960_),
    .S(_03642_),
    .X(_03961_));
 sky130_fd_sc_hd__clkbuf_1 _24607_ (.A(_03961_),
    .X(_00604_));
 sky130_fd_sc_hd__nor2_1 _24608_ (.A(_03954_),
    .B(_03956_),
    .Y(_03962_));
 sky130_fd_sc_hd__a21o_1 _24609_ (.A1(_03863_),
    .A2(_03957_),
    .B1(_03962_),
    .X(_03963_));
 sky130_fd_sc_hd__a21boi_1 _24610_ (.A1(_03948_),
    .A2(_03952_),
    .B1_N(_03950_),
    .Y(_03964_));
 sky130_fd_sc_hd__o21ba_1 _24611_ (.A1(_03948_),
    .A2(_03952_),
    .B1_N(_03964_),
    .X(_03965_));
 sky130_fd_sc_hd__a211o_1 _24612_ (.A1(_03890_),
    .A2(_03891_),
    .B1(_03892_),
    .C1(_03893_),
    .X(_03966_));
 sky130_fd_sc_hd__o21a_1 _24613_ (.A1(_03887_),
    .A2(_03895_),
    .B1(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__or2_1 _24614_ (.A(_03907_),
    .B(_03913_),
    .X(_03968_));
 sky130_fd_sc_hd__a21o_1 _24615_ (.A1(_03907_),
    .A2(_03913_),
    .B1(_03905_),
    .X(_03969_));
 sky130_fd_sc_hd__nand3_1 _24616_ (.A(_03967_),
    .B(_03968_),
    .C(_03969_),
    .Y(_03970_));
 sky130_fd_sc_hd__a21o_1 _24617_ (.A1(_03968_),
    .A2(_03969_),
    .B1(_03967_),
    .X(_03971_));
 sky130_fd_sc_hd__a211o_1 _24618_ (.A1(_03155_),
    .A2(_03156_),
    .B1(_03027_),
    .C1(_03028_),
    .X(_03972_));
 sky130_fd_sc_hd__o211ai_2 _24619_ (.A1(_03027_),
    .A2(_03028_),
    .B1(_03155_),
    .C1(_03156_),
    .Y(_03973_));
 sky130_fd_sc_hd__nand2_2 _24620_ (.A(_03972_),
    .B(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__nand2_1 _24621_ (.A(_03315_),
    .B(_03974_),
    .Y(_03975_));
 sky130_fd_sc_hd__a21oi_2 _24622_ (.A1(_03742_),
    .A2(_03827_),
    .B1(_03741_),
    .Y(_03976_));
 sky130_fd_sc_hd__a211o_1 _24623_ (.A1(_03972_),
    .A2(_03973_),
    .B1(_03047_),
    .C1(_03827_),
    .X(_03977_));
 sky130_fd_sc_hd__o21a_1 _24624_ (.A1(_03741_),
    .A2(_03974_),
    .B1(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__a21o_1 _24625_ (.A1(_03829_),
    .A2(_03974_),
    .B1(_03315_),
    .X(_03979_));
 sky130_fd_sc_hd__o221ai_4 _24626_ (.A1(_03975_),
    .A2(_03976_),
    .B1(_03978_),
    .B2(_03742_),
    .C1(_03979_),
    .Y(_03980_));
 sky130_fd_sc_hd__or2_2 _24627_ (.A(_03150_),
    .B(_03151_),
    .X(_03981_));
 sky130_fd_sc_hd__o211a_1 _24628_ (.A1(_03902_),
    .A2(_03903_),
    .B1(_03502_),
    .C1(_03981_),
    .X(_03982_));
 sky130_fd_sc_hd__a21o_1 _24629_ (.A1(_03902_),
    .A2(_03903_),
    .B1(_03982_),
    .X(_03983_));
 sky130_fd_sc_hd__nor2_1 _24630_ (.A(_03765_),
    .B(_03164_),
    .Y(_03984_));
 sky130_fd_sc_hd__o22a_1 _24631_ (.A1(_02994_),
    .A2(_02996_),
    .B1(_03029_),
    .B2(_03030_),
    .X(_03985_));
 sky130_fd_sc_hd__o22a_1 _24632_ (.A1(_02985_),
    .A2(_02987_),
    .B1(_03150_),
    .B2(_03151_),
    .X(_03986_));
 sky130_fd_sc_hd__xnor2_1 _24633_ (.A(_03985_),
    .B(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__xnor2_2 _24634_ (.A(_03984_),
    .B(_03987_),
    .Y(_03988_));
 sky130_fd_sc_hd__xnor2_1 _24635_ (.A(_03983_),
    .B(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__xnor2_2 _24636_ (.A(_03980_),
    .B(_03989_),
    .Y(_03990_));
 sky130_fd_sc_hd__a21o_1 _24637_ (.A1(_03970_),
    .A2(_03971_),
    .B1(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__nand3_2 _24638_ (.A(_03990_),
    .B(_03970_),
    .C(_03971_),
    .Y(_03992_));
 sky130_fd_sc_hd__nand2_2 _24639_ (.A(_03991_),
    .B(_03992_),
    .Y(_03993_));
 sky130_fd_sc_hd__o21ba_1 _24640_ (.A1(_03882_),
    .A2(_03897_),
    .B1_N(_03879_),
    .X(_03994_));
 sky130_fd_sc_hd__a21o_1 _24641_ (.A1(_03882_),
    .A2(_03897_),
    .B1(_03994_),
    .X(_03995_));
 sky130_fd_sc_hd__o22a_1 _24642_ (.A1(_03018_),
    .A2(_03019_),
    .B1(_03054_),
    .B2(_03055_),
    .X(_03996_));
 sky130_fd_sc_hd__o22a_1 _24643_ (.A1(_02979_),
    .A2(_02980_),
    .B1(_03061_),
    .B2(_03062_),
    .X(_03997_));
 sky130_fd_sc_hd__o22a_1 _24644_ (.A1(_03024_),
    .A2(_03025_),
    .B1(_03069_),
    .B2(_03071_),
    .X(_03998_));
 sky130_fd_sc_hd__xor2_1 _24645_ (.A(_03997_),
    .B(_03998_),
    .X(_03999_));
 sky130_fd_sc_hd__xnor2_1 _24646_ (.A(_03996_),
    .B(_03999_),
    .Y(_04000_));
 sky130_fd_sc_hd__a21o_1 _24647_ (.A1(_03883_),
    .A2(_03884_),
    .B1(_03885_),
    .X(_04001_));
 sky130_fd_sc_hd__or2_1 _24648_ (.A(_03883_),
    .B(_03884_),
    .X(_04002_));
 sky130_fd_sc_hd__a21oi_2 _24649_ (.A1(_03864_),
    .A2(_03865_),
    .B1(_03866_),
    .Y(_04003_));
 sky130_fd_sc_hd__nor2_1 _24650_ (.A(_03864_),
    .B(_03865_),
    .Y(_04004_));
 sky130_fd_sc_hd__a211o_1 _24651_ (.A1(_04001_),
    .A2(_04002_),
    .B1(_04003_),
    .C1(_04004_),
    .X(_04005_));
 sky130_fd_sc_hd__o211ai_1 _24652_ (.A1(_04003_),
    .A2(_04004_),
    .B1(_04001_),
    .C1(_04002_),
    .Y(_04006_));
 sky130_fd_sc_hd__and3_1 _24653_ (.A(_04000_),
    .B(_04005_),
    .C(_04006_),
    .X(_04007_));
 sky130_fd_sc_hd__a21oi_1 _24654_ (.A1(_04005_),
    .A2(_04006_),
    .B1(_04000_),
    .Y(_04008_));
 sky130_fd_sc_hd__a21bo_1 _24655_ (.A1(_03868_),
    .A2(_03877_),
    .B1_N(_03872_),
    .X(_04009_));
 sky130_fd_sc_hd__or2_1 _24656_ (.A(_03868_),
    .B(_03877_),
    .X(_04010_));
 sky130_fd_sc_hd__o211ai_2 _24657_ (.A1(_04007_),
    .A2(_04008_),
    .B1(_04009_),
    .C1(_04010_),
    .Y(_04011_));
 sky130_fd_sc_hd__a211o_1 _24658_ (.A1(_04009_),
    .A2(_04010_),
    .B1(_04007_),
    .C1(_04008_),
    .X(_04012_));
 sky130_fd_sc_hd__and2_1 _24659_ (.A(_03106_),
    .B(_03826_),
    .X(_04013_));
 sky130_fd_sc_hd__o22a_1 _24660_ (.A1(_03207_),
    .A2(_03208_),
    .B1(_03196_),
    .B2(_03197_),
    .X(_04014_));
 sky130_fd_sc_hd__o22a_1 _24661_ (.A1(_03057_),
    .A2(_03058_),
    .B1(_03717_),
    .B2(_03718_),
    .X(_04015_));
 sky130_fd_sc_hd__xor2_1 _24662_ (.A(_04014_),
    .B(_04015_),
    .X(_04016_));
 sky130_fd_sc_hd__xnor2_1 _24663_ (.A(_04013_),
    .B(_04016_),
    .Y(_04017_));
 sky130_fd_sc_hd__a21o_1 _24664_ (.A1(_03252_),
    .A2(_03825_),
    .B1(_03875_),
    .X(_04018_));
 sky130_fd_sc_hd__and3_1 _24665_ (.A(_03252_),
    .B(_03826_),
    .C(_03875_),
    .X(_04019_));
 sky130_fd_sc_hd__a21oi_2 _24666_ (.A1(_03874_),
    .A2(_04018_),
    .B1(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__o22a_2 _24667_ (.A1(_03004_),
    .A2(_03005_),
    .B1(_03103_),
    .B2(_03104_),
    .X(_04021_));
 sky130_fd_sc_hd__o22a_2 _24668_ (.A1(_02998_),
    .A2(_03000_),
    .B1(_03090_),
    .B2(_03091_),
    .X(_04022_));
 sky130_fd_sc_hd__o22a_1 _24669_ (.A1(_02989_),
    .A2(_02991_),
    .B1(_03093_),
    .B2(_03094_),
    .X(_04023_));
 sky130_fd_sc_hd__xor2_1 _24670_ (.A(_04022_),
    .B(_04023_),
    .X(_04024_));
 sky130_fd_sc_hd__xnor2_1 _24671_ (.A(_04021_),
    .B(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__xnor2_1 _24672_ (.A(_04020_),
    .B(_04025_),
    .Y(_04026_));
 sky130_fd_sc_hd__xnor2_1 _24673_ (.A(_04017_),
    .B(_04026_),
    .Y(_04027_));
 sky130_fd_sc_hd__a21boi_1 _24674_ (.A1(_04011_),
    .A2(_04012_),
    .B1_N(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__and3b_1 _24675_ (.A_N(_04027_),
    .B(_04011_),
    .C(_04012_),
    .X(_04029_));
 sky130_fd_sc_hd__or2_1 _24676_ (.A(_04028_),
    .B(_04029_),
    .X(_04030_));
 sky130_fd_sc_hd__xnor2_2 _24677_ (.A(_03995_),
    .B(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__xnor2_4 _24678_ (.A(_03993_),
    .B(_04031_),
    .Y(_04032_));
 sky130_fd_sc_hd__nand3b_2 _24679_ (.A_N(_03924_),
    .B(_03921_),
    .C(_03922_),
    .Y(_04033_));
 sky130_fd_sc_hd__a21boi_2 _24680_ (.A1(_03921_),
    .A2(_03922_),
    .B1_N(_03924_),
    .Y(_04034_));
 sky130_fd_sc_hd__a21oi_4 _24681_ (.A1(_03899_),
    .A2(_04033_),
    .B1(_04034_),
    .Y(_04035_));
 sky130_fd_sc_hd__nand2_1 _24682_ (.A(_03916_),
    .B(_03917_),
    .Y(_04036_));
 sky130_fd_sc_hd__o21a_1 _24683_ (.A1(_04036_),
    .A2(_03918_),
    .B1(_03915_),
    .X(_04037_));
 sky130_fd_sc_hd__a21oi_2 _24684_ (.A1(_04036_),
    .A2(_03918_),
    .B1(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__clkbuf_4 _24685_ (.A(_03908_),
    .X(_04039_));
 sky130_fd_sc_hd__or2_1 _24686_ (.A(_03910_),
    .B(_03911_),
    .X(_04040_));
 sky130_fd_sc_hd__a21oi_1 _24687_ (.A1(_03572_),
    .A2(_04040_),
    .B1(_03549_),
    .Y(_04041_));
 sky130_fd_sc_hd__and2_1 _24688_ (.A(_03910_),
    .B(_03911_),
    .X(_04042_));
 sky130_fd_sc_hd__o211a_1 _24689_ (.A1(_03572_),
    .A2(_04042_),
    .B1(_04040_),
    .C1(_03549_),
    .X(_04043_));
 sky130_fd_sc_hd__inv_2 _24690_ (.A(_04042_),
    .Y(_04044_));
 sky130_fd_sc_hd__o32a_2 _24691_ (.A1(_04039_),
    .A2(_04041_),
    .A3(_04043_),
    .B1(_03935_),
    .B2(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__xnor2_1 _24692_ (.A(_03942_),
    .B(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__xnor2_1 _24693_ (.A(_04038_),
    .B(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__xnor2_1 _24694_ (.A(_04035_),
    .B(_04047_),
    .Y(_04048_));
 sky130_fd_sc_hd__xnor2_2 _24695_ (.A(_04032_),
    .B(_04048_),
    .Y(_04049_));
 sky130_fd_sc_hd__inv_2 _24696_ (.A(_03946_),
    .Y(_04050_));
 sky130_fd_sc_hd__nor2_1 _24697_ (.A(_03931_),
    .B(_04050_),
    .Y(_04051_));
 sky130_fd_sc_hd__nand2_1 _24698_ (.A(_03931_),
    .B(_04050_),
    .Y(_04052_));
 sky130_fd_sc_hd__o21ai_1 _24699_ (.A1(_03928_),
    .A2(_04051_),
    .B1(_04052_),
    .Y(_04053_));
 sky130_fd_sc_hd__or2b_1 _24700_ (.A(_03944_),
    .B_N(_03939_),
    .X(_04054_));
 sky130_fd_sc_hd__and3_1 _24701_ (.A(_03937_),
    .B(_03938_),
    .C(_03944_),
    .X(_04055_));
 sky130_fd_sc_hd__a21oi_2 _24702_ (.A1(_03934_),
    .A2(_04054_),
    .B1(_04055_),
    .Y(_04056_));
 sky130_fd_sc_hd__xor2_1 _24703_ (.A(_04053_),
    .B(_04056_),
    .X(_04057_));
 sky130_fd_sc_hd__xnor2_1 _24704_ (.A(_04049_),
    .B(_04057_),
    .Y(_04058_));
 sky130_fd_sc_hd__and2b_1 _24705_ (.A_N(_03965_),
    .B(_04058_),
    .X(_04059_));
 sky130_fd_sc_hd__or2b_1 _24706_ (.A(_04058_),
    .B_N(_03965_),
    .X(_04060_));
 sky130_fd_sc_hd__or2b_1 _24707_ (.A(_04059_),
    .B_N(_04060_),
    .X(_04061_));
 sky130_fd_sc_hd__xnor2_1 _24708_ (.A(_03963_),
    .B(_04061_),
    .Y(_04062_));
 sky130_fd_sc_hd__mux2_1 _24709_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[4] ),
    .A1(_04062_),
    .S(_03642_),
    .X(_04063_));
 sky130_fd_sc_hd__clkbuf_1 _24710_ (.A(_04063_),
    .X(_00605_));
 sky130_fd_sc_hd__o21ai_1 _24711_ (.A1(_03963_),
    .A2(_04059_),
    .B1(_04060_),
    .Y(_04064_));
 sky130_fd_sc_hd__a21bo_1 _24712_ (.A1(_04049_),
    .A2(_04056_),
    .B1_N(_04053_),
    .X(_04065_));
 sky130_fd_sc_hd__o21a_1 _24713_ (.A1(_04049_),
    .A2(_04056_),
    .B1(_04065_),
    .X(_04066_));
 sky130_fd_sc_hd__xnor2_2 _24714_ (.A(_03315_),
    .B(_03974_),
    .Y(_04067_));
 sky130_fd_sc_hd__or2_1 _24715_ (.A(_03908_),
    .B(_04067_),
    .X(_04068_));
 sky130_fd_sc_hd__clkbuf_8 _24716_ (.A(_04068_),
    .X(_04069_));
 sky130_fd_sc_hd__a22o_1 _24717_ (.A1(_03502_),
    .A2(_03687_),
    .B1(_03985_),
    .B2(_03986_),
    .X(_04070_));
 sky130_fd_sc_hd__o21a_2 _24718_ (.A1(_03985_),
    .A2(_03986_),
    .B1(_04070_),
    .X(_04071_));
 sky130_fd_sc_hd__nor2_1 _24719_ (.A(_03765_),
    .B(_03743_),
    .Y(_04072_));
 sky130_fd_sc_hd__o22a_1 _24720_ (.A1(_02994_),
    .A2(_02996_),
    .B1(_03150_),
    .B2(_03151_),
    .X(_04073_));
 sky130_fd_sc_hd__o22a_1 _24721_ (.A1(_02985_),
    .A2(_02987_),
    .B1(_03162_),
    .B2(_03163_),
    .X(_04074_));
 sky130_fd_sc_hd__xnor2_1 _24722_ (.A(_04073_),
    .B(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__xnor2_2 _24723_ (.A(_04072_),
    .B(_04075_),
    .Y(_04076_));
 sky130_fd_sc_hd__xnor2_2 _24724_ (.A(_04071_),
    .B(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hd__xnor2_4 _24725_ (.A(_04069_),
    .B(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hd__nor2_1 _24726_ (.A(_03983_),
    .B(_03988_),
    .Y(_04079_));
 sky130_fd_sc_hd__nand2_1 _24727_ (.A(_03983_),
    .B(_03988_),
    .Y(_04080_));
 sky130_fd_sc_hd__o21ai_2 _24728_ (.A1(_03980_),
    .A2(_04079_),
    .B1(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__a21oi_1 _24729_ (.A1(_03883_),
    .A2(_03884_),
    .B1(_03885_),
    .Y(_04082_));
 sky130_fd_sc_hd__nor2_1 _24730_ (.A(_03883_),
    .B(_03884_),
    .Y(_04083_));
 sky130_fd_sc_hd__or4_1 _24731_ (.A(_04003_),
    .B(_04004_),
    .C(_04082_),
    .D(_04083_),
    .X(_04084_));
 sky130_fd_sc_hd__o22a_1 _24732_ (.A1(_04003_),
    .A2(_04004_),
    .B1(_04082_),
    .B2(_04083_),
    .X(_04085_));
 sky130_fd_sc_hd__a21o_2 _24733_ (.A1(_04000_),
    .A2(_04084_),
    .B1(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__xnor2_2 _24734_ (.A(_04081_),
    .B(_04086_),
    .Y(_04087_));
 sky130_fd_sc_hd__xor2_4 _24735_ (.A(_04078_),
    .B(_04087_),
    .X(_04088_));
 sky130_fd_sc_hd__a21boi_1 _24736_ (.A1(_04027_),
    .A2(_04012_),
    .B1_N(_04011_),
    .Y(_04089_));
 sky130_fd_sc_hd__nand2_1 _24737_ (.A(_03114_),
    .B(_03826_),
    .Y(_04090_));
 sky130_fd_sc_hd__nor2_1 _24738_ (.A(_03006_),
    .B(_03198_),
    .Y(_04091_));
 sky130_fd_sc_hd__nor2_1 _24739_ (.A(_03564_),
    .B(_03719_),
    .Y(_04092_));
 sky130_fd_sc_hd__xnor2_1 _24740_ (.A(_04091_),
    .B(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__xnor2_2 _24741_ (.A(_04090_),
    .B(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__a31o_1 _24742_ (.A1(_03106_),
    .A2(_03826_),
    .A3(_04014_),
    .B1(_04015_),
    .X(_04095_));
 sky130_fd_sc_hd__o21a_1 _24743_ (.A1(_04013_),
    .A2(_04014_),
    .B1(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__clkbuf_4 _24744_ (.A(_03799_),
    .X(_04097_));
 sky130_fd_sc_hd__nor2_1 _24745_ (.A(_03496_),
    .B(_04097_),
    .Y(_04098_));
 sky130_fd_sc_hd__o22a_1 _24746_ (.A1(_02989_),
    .A2(_02991_),
    .B1(_03090_),
    .B2(_03091_),
    .X(_04099_));
 sky130_fd_sc_hd__o22a_1 _24747_ (.A1(_02979_),
    .A2(_02980_),
    .B1(_03093_),
    .B2(_03094_),
    .X(_04100_));
 sky130_fd_sc_hd__xnor2_1 _24748_ (.A(_04099_),
    .B(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__xnor2_2 _24749_ (.A(_04098_),
    .B(_04101_),
    .Y(_04102_));
 sky130_fd_sc_hd__xnor2_1 _24750_ (.A(_04096_),
    .B(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__xnor2_2 _24751_ (.A(_04094_),
    .B(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hd__or2_1 _24752_ (.A(_04020_),
    .B(_04025_),
    .X(_04105_));
 sky130_fd_sc_hd__a21o_1 _24753_ (.A1(_04020_),
    .A2(_04025_),
    .B1(_04017_),
    .X(_04106_));
 sky130_fd_sc_hd__o22a_1 _24754_ (.A1(_03018_),
    .A2(_03019_),
    .B1(_03069_),
    .B2(_03071_),
    .X(_04107_));
 sky130_fd_sc_hd__o22a_1 _24755_ (.A1(_03054_),
    .A2(_03055_),
    .B1(_03029_),
    .B2(_03030_),
    .X(_04108_));
 sky130_fd_sc_hd__o22a_1 _24756_ (.A1(_03024_),
    .A2(_03025_),
    .B1(_03061_),
    .B2(_03062_),
    .X(_04109_));
 sky130_fd_sc_hd__xor2_1 _24757_ (.A(_04108_),
    .B(_04109_),
    .X(_04110_));
 sky130_fd_sc_hd__xnor2_2 _24758_ (.A(_04107_),
    .B(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__a21o_1 _24759_ (.A1(_04021_),
    .A2(_04022_),
    .B1(_04023_),
    .X(_04112_));
 sky130_fd_sc_hd__or2_1 _24760_ (.A(_04021_),
    .B(_04022_),
    .X(_04113_));
 sky130_fd_sc_hd__a21oi_2 _24761_ (.A1(_03996_),
    .A2(_03998_),
    .B1(_03997_),
    .Y(_04114_));
 sky130_fd_sc_hd__nor2_1 _24762_ (.A(_03996_),
    .B(_03998_),
    .Y(_04115_));
 sky130_fd_sc_hd__a211o_1 _24763_ (.A1(_04112_),
    .A2(_04113_),
    .B1(_04114_),
    .C1(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__o211ai_1 _24764_ (.A1(_04114_),
    .A2(_04115_),
    .B1(_04112_),
    .C1(_04113_),
    .Y(_04117_));
 sky130_fd_sc_hd__and3_1 _24765_ (.A(_04111_),
    .B(_04116_),
    .C(_04117_),
    .X(_04118_));
 sky130_fd_sc_hd__a21oi_1 _24766_ (.A1(_04116_),
    .A2(_04117_),
    .B1(_04111_),
    .Y(_04119_));
 sky130_fd_sc_hd__a211o_1 _24767_ (.A1(_04105_),
    .A2(_04106_),
    .B1(_04118_),
    .C1(_04119_),
    .X(_04120_));
 sky130_fd_sc_hd__o211ai_1 _24768_ (.A1(_04118_),
    .A2(_04119_),
    .B1(_04105_),
    .C1(_04106_),
    .Y(_04121_));
 sky130_fd_sc_hd__nand2_1 _24769_ (.A(_04120_),
    .B(_04121_),
    .Y(_04122_));
 sky130_fd_sc_hd__xnor2_2 _24770_ (.A(_04104_),
    .B(_04122_),
    .Y(_04123_));
 sky130_fd_sc_hd__xnor2_1 _24771_ (.A(_04089_),
    .B(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__xnor2_2 _24772_ (.A(_04088_),
    .B(_04124_),
    .Y(_04125_));
 sky130_fd_sc_hd__a211o_1 _24773_ (.A1(_03991_),
    .A2(_03992_),
    .B1(_04028_),
    .C1(_04029_),
    .X(_04126_));
 sky130_fd_sc_hd__o211a_1 _24774_ (.A1(_04028_),
    .A2(_04029_),
    .B1(_03991_),
    .C1(_03992_),
    .X(_04127_));
 sky130_fd_sc_hd__a21oi_1 _24775_ (.A1(_03995_),
    .A2(_04126_),
    .B1(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__a21oi_1 _24776_ (.A1(_03572_),
    .A2(_04040_),
    .B1(_04042_),
    .Y(_04129_));
 sky130_fd_sc_hd__nor2_1 _24777_ (.A(_03830_),
    .B(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__clkbuf_4 _24778_ (.A(_03743_),
    .X(_04131_));
 sky130_fd_sc_hd__o22a_1 _24779_ (.A1(_03017_),
    .A2(_03185_),
    .B1(_04131_),
    .B2(_03047_),
    .X(_04132_));
 sky130_fd_sc_hd__a21oi_1 _24780_ (.A1(_03017_),
    .A2(_03185_),
    .B1(_04132_),
    .Y(_04133_));
 sky130_fd_sc_hd__xnor2_1 _24781_ (.A(_03549_),
    .B(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hd__nor2_2 _24782_ (.A(_04039_),
    .B(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__xnor2_1 _24783_ (.A(_04130_),
    .B(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__inv_2 _24784_ (.A(_03990_),
    .Y(_04137_));
 sky130_fd_sc_hd__a21bo_1 _24785_ (.A1(_04137_),
    .A2(_03971_),
    .B1_N(_03970_),
    .X(_04138_));
 sky130_fd_sc_hd__xnor2_2 _24786_ (.A(_04136_),
    .B(_04138_),
    .Y(_04139_));
 sky130_fd_sc_hd__xnor2_1 _24787_ (.A(_04128_),
    .B(_04139_),
    .Y(_04140_));
 sky130_fd_sc_hd__xnor2_2 _24788_ (.A(_04125_),
    .B(_04140_),
    .Y(_04141_));
 sky130_fd_sc_hd__nand2_2 _24789_ (.A(_04038_),
    .B(_04045_),
    .Y(_04142_));
 sky130_fd_sc_hd__nor2_1 _24790_ (.A(_04038_),
    .B(_04045_),
    .Y(_04143_));
 sky130_fd_sc_hd__a21o_1 _24791_ (.A1(_04035_),
    .A2(_04142_),
    .B1(_04143_),
    .X(_04144_));
 sky130_fd_sc_hd__a21o_1 _24792_ (.A1(_03940_),
    .A2(_03941_),
    .B1(_03830_),
    .X(_04145_));
 sky130_fd_sc_hd__o221ai_2 _24793_ (.A1(_04035_),
    .A2(_04142_),
    .B1(_04144_),
    .B2(_04032_),
    .C1(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__and2_1 _24794_ (.A(_04035_),
    .B(_04143_),
    .X(_04147_));
 sky130_fd_sc_hd__a211o_1 _24795_ (.A1(_04032_),
    .A2(_04144_),
    .B1(_04147_),
    .C1(_04145_),
    .X(_04148_));
 sky130_fd_sc_hd__nor2_1 _24796_ (.A(_04035_),
    .B(_04142_),
    .Y(_04149_));
 sky130_fd_sc_hd__mux2_1 _24797_ (.A0(_04149_),
    .A1(_04147_),
    .S(_04032_),
    .X(_04150_));
 sky130_fd_sc_hd__a21o_1 _24798_ (.A1(_04146_),
    .A2(_04148_),
    .B1(_04150_),
    .X(_04151_));
 sky130_fd_sc_hd__xnor2_2 _24799_ (.A(_04141_),
    .B(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__xor2_1 _24800_ (.A(_04066_),
    .B(_04152_),
    .X(_04153_));
 sky130_fd_sc_hd__xnor2_1 _24801_ (.A(_04064_),
    .B(_04153_),
    .Y(_04154_));
 sky130_fd_sc_hd__mux2_1 _24802_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[5] ),
    .A1(_04154_),
    .S(_03642_),
    .X(_04155_));
 sky130_fd_sc_hd__clkbuf_1 _24803_ (.A(_04155_),
    .X(_00606_));
 sky130_fd_sc_hd__nor2_1 _24804_ (.A(_04066_),
    .B(_04152_),
    .Y(_04156_));
 sky130_fd_sc_hd__nand2_1 _24805_ (.A(_04066_),
    .B(_04152_),
    .Y(_04157_));
 sky130_fd_sc_hd__o21ai_1 _24806_ (.A1(_04064_),
    .A2(_04156_),
    .B1(_04157_),
    .Y(_04158_));
 sky130_fd_sc_hd__and2_1 _24807_ (.A(_04035_),
    .B(_04032_),
    .X(_04159_));
 sky130_fd_sc_hd__o21ai_1 _24808_ (.A1(_04035_),
    .A2(_04032_),
    .B1(_03942_),
    .Y(_04160_));
 sky130_fd_sc_hd__or2b_1 _24809_ (.A(_04159_),
    .B_N(_04160_),
    .X(_04161_));
 sky130_fd_sc_hd__or2_1 _24810_ (.A(_04141_),
    .B(_04143_),
    .X(_04162_));
 sky130_fd_sc_hd__o21a_1 _24811_ (.A1(_04035_),
    .A2(_04032_),
    .B1(_04142_),
    .X(_04163_));
 sky130_fd_sc_hd__o21a_1 _24812_ (.A1(_04143_),
    .A2(_04163_),
    .B1(_04141_),
    .X(_04164_));
 sky130_fd_sc_hd__o211a_1 _24813_ (.A1(_04141_),
    .A2(_04159_),
    .B1(_04142_),
    .C1(_03942_),
    .X(_04165_));
 sky130_fd_sc_hd__a211o_1 _24814_ (.A1(_04161_),
    .A2(_04162_),
    .B1(_04164_),
    .C1(_04165_),
    .X(_04166_));
 sky130_fd_sc_hd__a21o_1 _24815_ (.A1(_04125_),
    .A2(_04139_),
    .B1(_04128_),
    .X(_04167_));
 sky130_fd_sc_hd__o21a_1 _24816_ (.A1(_04125_),
    .A2(_04139_),
    .B1(_04167_),
    .X(_04168_));
 sky130_fd_sc_hd__a21bo_1 _24817_ (.A1(_04088_),
    .A2(_04123_),
    .B1_N(_04089_),
    .X(_04169_));
 sky130_fd_sc_hd__o21ai_4 _24818_ (.A1(_04088_),
    .A2(_04123_),
    .B1(_04169_),
    .Y(_04170_));
 sky130_fd_sc_hd__o21ba_1 _24819_ (.A1(_04078_),
    .A2(_04086_),
    .B1_N(_04081_),
    .X(_04171_));
 sky130_fd_sc_hd__a21oi_2 _24820_ (.A1(_04078_),
    .A2(_04086_),
    .B1(_04171_),
    .Y(_04172_));
 sky130_fd_sc_hd__or2_1 _24821_ (.A(_03741_),
    .B(_03742_),
    .X(_04173_));
 sky130_fd_sc_hd__buf_2 _24822_ (.A(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__a21oi_1 _24823_ (.A1(_03157_),
    .A2(_03572_),
    .B1(_03315_),
    .Y(_04175_));
 sky130_fd_sc_hd__a21oi_2 _24824_ (.A1(_03017_),
    .A2(_03185_),
    .B1(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hd__o21a_2 _24825_ (.A1(_03549_),
    .A2(_04176_),
    .B1(_03829_),
    .X(_04177_));
 sky130_fd_sc_hd__o31a_2 _24826_ (.A1(_03161_),
    .A2(_04174_),
    .A3(_03975_),
    .B1(_04177_),
    .X(_04178_));
 sky130_fd_sc_hd__xor2_1 _24827_ (.A(_04172_),
    .B(_04178_),
    .X(_04179_));
 sky130_fd_sc_hd__nand2_2 _24828_ (.A(_03564_),
    .B(_03826_),
    .Y(_04180_));
 sky130_fd_sc_hd__nand2_2 _24829_ (.A(_03313_),
    .B(_03720_),
    .Y(_04181_));
 sky130_fd_sc_hd__clkbuf_4 _24830_ (.A(_03719_),
    .X(_04182_));
 sky130_fd_sc_hd__nor2_1 _24831_ (.A(_03006_),
    .B(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__xor2_1 _24832_ (.A(_04181_),
    .B(_04183_),
    .X(_04184_));
 sky130_fd_sc_hd__xnor2_2 _24833_ (.A(_04180_),
    .B(_04184_),
    .Y(_04185_));
 sky130_fd_sc_hd__a21bo_1 _24834_ (.A1(_04091_),
    .A2(_04092_),
    .B1_N(_04090_),
    .X(_04186_));
 sky130_fd_sc_hd__o21a_1 _24835_ (.A1(_04091_),
    .A2(_04092_),
    .B1(_04186_),
    .X(_04187_));
 sky130_fd_sc_hd__nor2_1 _24836_ (.A(_03474_),
    .B(_04097_),
    .Y(_04188_));
 sky130_fd_sc_hd__nor2_1 _24837_ (.A(_03343_),
    .B(_03200_),
    .Y(_04189_));
 sky130_fd_sc_hd__nor2_4 _24838_ (.A(_03090_),
    .B(_03091_),
    .Y(_04190_));
 sky130_fd_sc_hd__nor2_1 _24839_ (.A(_02982_),
    .B(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__xnor2_1 _24840_ (.A(_04189_),
    .B(_04191_),
    .Y(_04192_));
 sky130_fd_sc_hd__xnor2_1 _24841_ (.A(_04188_),
    .B(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__xnor2_1 _24842_ (.A(_04187_),
    .B(_04193_),
    .Y(_04194_));
 sky130_fd_sc_hd__xnor2_2 _24843_ (.A(_04185_),
    .B(_04194_),
    .Y(_04195_));
 sky130_fd_sc_hd__nor2_1 _24844_ (.A(_04096_),
    .B(_04102_),
    .Y(_04196_));
 sky130_fd_sc_hd__nand2_1 _24845_ (.A(_04096_),
    .B(_04102_),
    .Y(_04197_));
 sky130_fd_sc_hd__o21ai_2 _24846_ (.A1(_04094_),
    .A2(_04196_),
    .B1(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__nor2_2 _24847_ (.A(_03325_),
    .B(_03900_),
    .Y(_04199_));
 sky130_fd_sc_hd__nor2_1 _24848_ (.A(_03254_),
    .B(_03280_),
    .Y(_04200_));
 sky130_fd_sc_hd__nor2_1 _24849_ (.A(net1017),
    .B(_03112_),
    .Y(_04201_));
 sky130_fd_sc_hd__xnor2_1 _24850_ (.A(_04200_),
    .B(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__xnor2_2 _24851_ (.A(_04199_),
    .B(_04202_),
    .Y(_04203_));
 sky130_fd_sc_hd__a21o_1 _24852_ (.A1(_03313_),
    .A2(_03889_),
    .B1(_04099_),
    .X(_04204_));
 sky130_fd_sc_hd__and3_1 _24853_ (.A(_03313_),
    .B(_03889_),
    .C(_04099_),
    .X(_04205_));
 sky130_fd_sc_hd__a21o_1 _24854_ (.A1(_04100_),
    .A2(_04204_),
    .B1(_04205_),
    .X(_04206_));
 sky130_fd_sc_hd__a21o_1 _24855_ (.A1(_04107_),
    .A2(_04108_),
    .B1(_04109_),
    .X(_04207_));
 sky130_fd_sc_hd__o21a_1 _24856_ (.A1(_04107_),
    .A2(_04108_),
    .B1(_04207_),
    .X(_04208_));
 sky130_fd_sc_hd__xnor2_1 _24857_ (.A(_04206_),
    .B(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__xnor2_2 _24858_ (.A(_04203_),
    .B(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__xnor2_1 _24859_ (.A(_04198_),
    .B(_04210_),
    .Y(_04211_));
 sky130_fd_sc_hd__xnor2_2 _24860_ (.A(_04195_),
    .B(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__o211a_1 _24861_ (.A1(_04118_),
    .A2(_04119_),
    .B1(_04105_),
    .C1(_04106_),
    .X(_04213_));
 sky130_fd_sc_hd__a21oi_1 _24862_ (.A1(_04104_),
    .A2(_04120_),
    .B1(_04213_),
    .Y(_04214_));
 sky130_fd_sc_hd__or2_1 _24863_ (.A(_04071_),
    .B(_04076_),
    .X(_04215_));
 sky130_fd_sc_hd__nand2_1 _24864_ (.A(_04071_),
    .B(_04076_),
    .Y(_04216_));
 sky130_fd_sc_hd__mux2_1 _24865_ (.A0(_04215_),
    .A1(_04216_),
    .S(_04069_),
    .X(_04217_));
 sky130_fd_sc_hd__nor2_1 _24866_ (.A(_03765_),
    .B(_03908_),
    .Y(_04218_));
 sky130_fd_sc_hd__o22a_1 _24867_ (.A1(_02994_),
    .A2(_02996_),
    .B1(_03162_),
    .B2(_03163_),
    .X(_04219_));
 sky130_fd_sc_hd__o22a_1 _24868_ (.A1(_02985_),
    .A2(_02987_),
    .B1(_03741_),
    .B2(_03742_),
    .X(_04220_));
 sky130_fd_sc_hd__xnor2_1 _24869_ (.A(_04219_),
    .B(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__xnor2_2 _24870_ (.A(_04218_),
    .B(_04221_),
    .Y(_04222_));
 sky130_fd_sc_hd__and2_1 _24871_ (.A(_04073_),
    .B(_04074_),
    .X(_04223_));
 sky130_fd_sc_hd__nor2_1 _24872_ (.A(_04073_),
    .B(_04074_),
    .Y(_04224_));
 sky130_fd_sc_hd__o21ba_1 _24873_ (.A1(_04072_),
    .A2(_04223_),
    .B1_N(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__xnor2_2 _24874_ (.A(_04222_),
    .B(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__a21oi_1 _24875_ (.A1(_04021_),
    .A2(_04022_),
    .B1(_04023_),
    .Y(_04227_));
 sky130_fd_sc_hd__nor2_1 _24876_ (.A(_04021_),
    .B(_04022_),
    .Y(_04228_));
 sky130_fd_sc_hd__or4_1 _24877_ (.A(_04114_),
    .B(_04115_),
    .C(_04227_),
    .D(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__o22a_1 _24878_ (.A1(_04114_),
    .A2(_04115_),
    .B1(_04227_),
    .B2(_04228_),
    .X(_04230_));
 sky130_fd_sc_hd__a21o_2 _24879_ (.A1(_04111_),
    .A2(_04229_),
    .B1(_04230_),
    .X(_04231_));
 sky130_fd_sc_hd__xnor2_1 _24880_ (.A(_04226_),
    .B(_04231_),
    .Y(_04232_));
 sky130_fd_sc_hd__xnor2_2 _24881_ (.A(_04217_),
    .B(_04232_),
    .Y(_04233_));
 sky130_fd_sc_hd__xnor2_1 _24882_ (.A(_04214_),
    .B(_04233_),
    .Y(_04234_));
 sky130_fd_sc_hd__xnor2_2 _24883_ (.A(_04212_),
    .B(_04234_),
    .Y(_04235_));
 sky130_fd_sc_hd__xnor2_1 _24884_ (.A(_04179_),
    .B(_04235_),
    .Y(_04236_));
 sky130_fd_sc_hd__xnor2_2 _24885_ (.A(_04170_),
    .B(_04236_),
    .Y(_04237_));
 sky130_fd_sc_hd__a21o_1 _24886_ (.A1(_04130_),
    .A2(_04135_),
    .B1(_04138_),
    .X(_04238_));
 sky130_fd_sc_hd__o21a_1 _24887_ (.A1(_04130_),
    .A2(_04135_),
    .B1(_04238_),
    .X(_04239_));
 sky130_fd_sc_hd__xnor2_1 _24888_ (.A(_04237_),
    .B(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__xnor2_2 _24889_ (.A(_04168_),
    .B(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__xnor2_1 _24890_ (.A(_04166_),
    .B(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__xnor2_1 _24891_ (.A(_04158_),
    .B(_04242_),
    .Y(_04243_));
 sky130_fd_sc_hd__mux2_1 _24892_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[6] ),
    .A1(_04243_),
    .S(_03642_),
    .X(_04244_));
 sky130_fd_sc_hd__clkbuf_1 _24893_ (.A(_04244_),
    .X(_00607_));
 sky130_fd_sc_hd__nor2_1 _24894_ (.A(_04166_),
    .B(_04241_),
    .Y(_04245_));
 sky130_fd_sc_hd__nor3_1 _24895_ (.A(_03959_),
    .B(_04061_),
    .C(_04245_),
    .Y(_04246_));
 sky130_fd_sc_hd__nand2_1 _24896_ (.A(_04166_),
    .B(_04241_),
    .Y(_04247_));
 sky130_fd_sc_hd__o21ai_1 _24897_ (.A1(_03962_),
    .A2(_04059_),
    .B1(_04060_),
    .Y(_04248_));
 sky130_fd_sc_hd__a21o_1 _24898_ (.A1(_04156_),
    .A2(_04247_),
    .B1(_04245_),
    .X(_04249_));
 sky130_fd_sc_hd__a31oi_1 _24899_ (.A1(_04157_),
    .A2(_04247_),
    .A3(_04248_),
    .B1(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__a31o_1 _24900_ (.A1(_03863_),
    .A2(_04153_),
    .A3(_04246_),
    .B1(_04250_),
    .X(_04251_));
 sky130_fd_sc_hd__buf_2 _24901_ (.A(_03011_),
    .X(_04252_));
 sky130_fd_sc_hd__xnor2_1 _24902_ (.A(_03355_),
    .B(_03765_),
    .Y(_04253_));
 sky130_fd_sc_hd__nand2_1 _24903_ (.A(_04252_),
    .B(_04253_),
    .Y(_04254_));
 sky130_fd_sc_hd__o22a_1 _24904_ (.A1(_04252_),
    .A2(_03741_),
    .B1(_03742_),
    .B2(_04254_),
    .X(_04255_));
 sky130_fd_sc_hd__a21o_1 _24905_ (.A1(_04252_),
    .A2(_04174_),
    .B1(_04253_),
    .X(_04256_));
 sky130_fd_sc_hd__o221a_4 _24906_ (.A1(_03976_),
    .A2(_04254_),
    .B1(_04255_),
    .B2(_03827_),
    .C1(_04256_),
    .X(_04257_));
 sky130_fd_sc_hd__nor2_4 _24907_ (.A(_04039_),
    .B(_04067_),
    .Y(_04258_));
 sky130_fd_sc_hd__a21o_1 _24908_ (.A1(_04219_),
    .A2(_04220_),
    .B1(_04218_),
    .X(_04259_));
 sky130_fd_sc_hd__o21a_2 _24909_ (.A1(_04219_),
    .A2(_04220_),
    .B1(_04259_),
    .X(_04260_));
 sky130_fd_sc_hd__xnor2_2 _24910_ (.A(_04258_),
    .B(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__xnor2_4 _24911_ (.A(_04257_),
    .B(_04261_),
    .Y(_04262_));
 sky130_fd_sc_hd__a21o_1 _24912_ (.A1(_04222_),
    .A2(_04225_),
    .B1(_04258_),
    .X(_04263_));
 sky130_fd_sc_hd__o21a_1 _24913_ (.A1(_04222_),
    .A2(_04225_),
    .B1(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__a21o_1 _24914_ (.A1(_04206_),
    .A2(_04208_),
    .B1(_04203_),
    .X(_04265_));
 sky130_fd_sc_hd__o21a_1 _24915_ (.A1(_04206_),
    .A2(_04208_),
    .B1(_04265_),
    .X(_04266_));
 sky130_fd_sc_hd__xnor2_2 _24916_ (.A(_04264_),
    .B(_04266_),
    .Y(_04267_));
 sky130_fd_sc_hd__xnor2_4 _24917_ (.A(_04262_),
    .B(_04267_),
    .Y(_04268_));
 sky130_fd_sc_hd__o21ba_1 _24918_ (.A1(_04198_),
    .A2(_04210_),
    .B1_N(_04195_),
    .X(_04269_));
 sky130_fd_sc_hd__a21oi_2 _24919_ (.A1(_04198_),
    .A2(_04210_),
    .B1(_04269_),
    .Y(_04270_));
 sky130_fd_sc_hd__nand2_1 _24920_ (.A(_03006_),
    .B(_03826_),
    .Y(_04271_));
 sky130_fd_sc_hd__buf_4 _24921_ (.A(_03198_),
    .X(_04272_));
 sky130_fd_sc_hd__nor2_1 _24922_ (.A(_03474_),
    .B(_04272_),
    .Y(_04273_));
 sky130_fd_sc_hd__nor2_1 _24923_ (.A(_03496_),
    .B(_04182_),
    .Y(_04274_));
 sky130_fd_sc_hd__xnor2_1 _24924_ (.A(_04273_),
    .B(_04274_),
    .Y(_04275_));
 sky130_fd_sc_hd__xnor2_2 _24925_ (.A(_04271_),
    .B(_04275_),
    .Y(_04276_));
 sky130_fd_sc_hd__o21ba_1 _24926_ (.A1(_04180_),
    .A2(_04181_),
    .B1_N(_04183_),
    .X(_04277_));
 sky130_fd_sc_hd__a21oi_2 _24927_ (.A1(_04180_),
    .A2(_04181_),
    .B1(_04277_),
    .Y(_04278_));
 sky130_fd_sc_hd__nor2_1 _24928_ (.A(_02982_),
    .B(_04097_),
    .Y(_04279_));
 sky130_fd_sc_hd__nor2_1 _24929_ (.A(net1017),
    .B(_03200_),
    .Y(_04280_));
 sky130_fd_sc_hd__nor2_1 _24930_ (.A(_03343_),
    .B(_04190_),
    .Y(_04281_));
 sky130_fd_sc_hd__xnor2_1 _24931_ (.A(_04280_),
    .B(_04281_),
    .Y(_04282_));
 sky130_fd_sc_hd__xnor2_2 _24932_ (.A(_04279_),
    .B(_04282_),
    .Y(_04283_));
 sky130_fd_sc_hd__xnor2_1 _24933_ (.A(_04278_),
    .B(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__xnor2_2 _24934_ (.A(_04276_),
    .B(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__a21bo_1 _24935_ (.A1(_04187_),
    .A2(_04193_),
    .B1_N(_04185_),
    .X(_04286_));
 sky130_fd_sc_hd__o21a_1 _24936_ (.A1(_04187_),
    .A2(_04193_),
    .B1(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__clkbuf_4 _24937_ (.A(_03164_),
    .X(_04288_));
 sky130_fd_sc_hd__nor2_1 _24938_ (.A(_03325_),
    .B(_04288_),
    .Y(_04289_));
 sky130_fd_sc_hd__nor2_1 _24939_ (.A(_03112_),
    .B(_03280_),
    .Y(_04290_));
 sky130_fd_sc_hd__nor2_1 _24940_ (.A(_03254_),
    .B(_03900_),
    .Y(_04291_));
 sky130_fd_sc_hd__xnor2_1 _24941_ (.A(_04290_),
    .B(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hd__xnor2_2 _24942_ (.A(_04289_),
    .B(_04292_),
    .Y(_04293_));
 sky130_fd_sc_hd__a21o_1 _24943_ (.A1(_04188_),
    .A2(_04191_),
    .B1(_04189_),
    .X(_04294_));
 sky130_fd_sc_hd__o21a_1 _24944_ (.A1(_04188_),
    .A2(_04191_),
    .B1(_04294_),
    .X(_04295_));
 sky130_fd_sc_hd__a21o_1 _24945_ (.A1(_04199_),
    .A2(_04200_),
    .B1(_04201_),
    .X(_04296_));
 sky130_fd_sc_hd__o21a_1 _24946_ (.A1(_04199_),
    .A2(_04200_),
    .B1(_04296_),
    .X(_04297_));
 sky130_fd_sc_hd__xnor2_1 _24947_ (.A(_04295_),
    .B(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hd__xnor2_2 _24948_ (.A(_04293_),
    .B(_04298_),
    .Y(_04299_));
 sky130_fd_sc_hd__xor2_1 _24949_ (.A(_04287_),
    .B(_04299_),
    .X(_04300_));
 sky130_fd_sc_hd__xnor2_2 _24950_ (.A(_04285_),
    .B(_04300_),
    .Y(_04301_));
 sky130_fd_sc_hd__xor2_2 _24951_ (.A(_04270_),
    .B(_04301_),
    .X(_04302_));
 sky130_fd_sc_hd__xnor2_4 _24952_ (.A(_04268_),
    .B(_04302_),
    .Y(_04303_));
 sky130_fd_sc_hd__o21ba_1 _24953_ (.A1(_04212_),
    .A2(_04233_),
    .B1_N(_04214_),
    .X(_04304_));
 sky130_fd_sc_hd__a21o_1 _24954_ (.A1(_04212_),
    .A2(_04233_),
    .B1(_04304_),
    .X(_04305_));
 sky130_fd_sc_hd__o21ai_4 _24955_ (.A1(_03549_),
    .A2(_04176_),
    .B1(_03829_),
    .Y(_04306_));
 sky130_fd_sc_hd__nor2_1 _24956_ (.A(_04071_),
    .B(_04076_),
    .Y(_04307_));
 sky130_fd_sc_hd__o21a_1 _24957_ (.A1(_04226_),
    .A2(_04231_),
    .B1(_04216_),
    .X(_04308_));
 sky130_fd_sc_hd__a21o_1 _24958_ (.A1(_04226_),
    .A2(_04231_),
    .B1(_04308_),
    .X(_04309_));
 sky130_fd_sc_hd__inv_2 _24959_ (.A(_04226_),
    .Y(_04310_));
 sky130_fd_sc_hd__o211a_1 _24960_ (.A1(_04307_),
    .A2(_04231_),
    .B1(_04258_),
    .C1(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__a221o_1 _24961_ (.A1(_04307_),
    .A2(_04231_),
    .B1(_04309_),
    .B2(_04069_),
    .C1(_04311_),
    .X(_04312_));
 sky130_fd_sc_hd__xnor2_1 _24962_ (.A(_04306_),
    .B(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__xnor2_1 _24963_ (.A(_04305_),
    .B(_04313_),
    .Y(_04314_));
 sky130_fd_sc_hd__xnor2_2 _24964_ (.A(_04303_),
    .B(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hd__or2_1 _24965_ (.A(_04172_),
    .B(_04178_),
    .X(_04316_));
 sky130_fd_sc_hd__and2_1 _24966_ (.A(_04172_),
    .B(_04178_),
    .X(_04317_));
 sky130_fd_sc_hd__a21o_1 _24967_ (.A1(_04170_),
    .A2(_04316_),
    .B1(_04317_),
    .X(_04318_));
 sky130_fd_sc_hd__nand2_1 _24968_ (.A(_04235_),
    .B(_04317_),
    .Y(_04319_));
 sky130_fd_sc_hd__mux2_1 _24969_ (.A0(_04316_),
    .A1(_04319_),
    .S(_04170_),
    .X(_04320_));
 sky130_fd_sc_hd__o21a_1 _24970_ (.A1(_04235_),
    .A2(_04318_),
    .B1(_04320_),
    .X(_04321_));
 sky130_fd_sc_hd__xnor2_1 _24971_ (.A(_04315_),
    .B(_04321_),
    .Y(_04322_));
 sky130_fd_sc_hd__o21a_1 _24972_ (.A1(_04237_),
    .A2(_04239_),
    .B1(_04168_),
    .X(_04323_));
 sky130_fd_sc_hd__a21oi_1 _24973_ (.A1(_04237_),
    .A2(_04239_),
    .B1(_04323_),
    .Y(_04324_));
 sky130_fd_sc_hd__nand2_1 _24974_ (.A(_04322_),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__or2_1 _24975_ (.A(_04322_),
    .B(_04324_),
    .X(_04326_));
 sky130_fd_sc_hd__nand2_1 _24976_ (.A(_04325_),
    .B(_04326_),
    .Y(_04327_));
 sky130_fd_sc_hd__xnor2_1 _24977_ (.A(_04251_),
    .B(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__mux2_1 _24978_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[7] ),
    .A1(_04328_),
    .S(_03642_),
    .X(_04329_));
 sky130_fd_sc_hd__clkbuf_1 _24979_ (.A(_04329_),
    .X(_00608_));
 sky130_fd_sc_hd__nor2_1 _24980_ (.A(_04322_),
    .B(_04324_),
    .Y(_04330_));
 sky130_fd_sc_hd__a21oi_1 _24981_ (.A1(_04251_),
    .A2(_04325_),
    .B1(_04330_),
    .Y(_04331_));
 sky130_fd_sc_hd__or2_1 _24982_ (.A(_04315_),
    .B(_04317_),
    .X(_04332_));
 sky130_fd_sc_hd__a22o_1 _24983_ (.A1(_04315_),
    .A2(_04316_),
    .B1(_04332_),
    .B2(_04170_),
    .X(_04333_));
 sky130_fd_sc_hd__a22o_1 _24984_ (.A1(_04315_),
    .A2(_04318_),
    .B1(_04333_),
    .B2(_04235_),
    .X(_04334_));
 sky130_fd_sc_hd__a21o_1 _24985_ (.A1(_04257_),
    .A2(_04260_),
    .B1(_04258_),
    .X(_04335_));
 sky130_fd_sc_hd__o21ai_4 _24986_ (.A1(_04257_),
    .A2(_04260_),
    .B1(_04335_),
    .Y(_04336_));
 sky130_fd_sc_hd__a21oi_1 _24987_ (.A1(_03234_),
    .A2(_04174_),
    .B1(_03765_),
    .Y(_04337_));
 sky130_fd_sc_hd__a21o_1 _24988_ (.A1(_03355_),
    .A2(_04131_),
    .B1(_04337_),
    .X(_04338_));
 sky130_fd_sc_hd__a31o_1 _24989_ (.A1(_03234_),
    .A2(_03007_),
    .A3(_03765_),
    .B1(_04039_),
    .X(_04339_));
 sky130_fd_sc_hd__a21oi_1 _24990_ (.A1(_04252_),
    .A2(_04338_),
    .B1(_04339_),
    .Y(_04340_));
 sky130_fd_sc_hd__xnor2_1 _24991_ (.A(_04069_),
    .B(_04340_),
    .Y(_04341_));
 sky130_fd_sc_hd__a21o_1 _24992_ (.A1(_04295_),
    .A2(_04297_),
    .B1(_04293_),
    .X(_04342_));
 sky130_fd_sc_hd__o21a_1 _24993_ (.A1(_04295_),
    .A2(_04297_),
    .B1(_04342_),
    .X(_04343_));
 sky130_fd_sc_hd__nor2_1 _24994_ (.A(_04341_),
    .B(_04343_),
    .Y(_04344_));
 sky130_fd_sc_hd__and2_1 _24995_ (.A(_04341_),
    .B(_04343_),
    .X(_04345_));
 sky130_fd_sc_hd__or2_2 _24996_ (.A(_04344_),
    .B(_04345_),
    .X(_04346_));
 sky130_fd_sc_hd__xor2_4 _24997_ (.A(_04336_),
    .B(_04346_),
    .X(_04347_));
 sky130_fd_sc_hd__nand2_1 _24998_ (.A(_03496_),
    .B(_03826_),
    .Y(_04348_));
 sky130_fd_sc_hd__nor2_1 _24999_ (.A(_02982_),
    .B(_04272_),
    .Y(_04349_));
 sky130_fd_sc_hd__nor2_1 _25000_ (.A(_03474_),
    .B(_03719_),
    .Y(_04350_));
 sky130_fd_sc_hd__xnor2_1 _25001_ (.A(_04349_),
    .B(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__xnor2_1 _25002_ (.A(_04348_),
    .B(_04351_),
    .Y(_04352_));
 sky130_fd_sc_hd__a21bo_1 _25003_ (.A1(_04273_),
    .A2(_04274_),
    .B1_N(_04271_),
    .X(_04353_));
 sky130_fd_sc_hd__o21a_1 _25004_ (.A1(_04273_),
    .A2(_04274_),
    .B1(_04353_),
    .X(_04354_));
 sky130_fd_sc_hd__nor2_2 _25005_ (.A(_03343_),
    .B(_04097_),
    .Y(_04355_));
 sky130_fd_sc_hd__nor2_1 _25006_ (.A(_03280_),
    .B(_03200_),
    .Y(_04356_));
 sky130_fd_sc_hd__nor2_1 _25007_ (.A(net1017),
    .B(_04190_),
    .Y(_04357_));
 sky130_fd_sc_hd__xnor2_1 _25008_ (.A(_04356_),
    .B(_04357_),
    .Y(_04358_));
 sky130_fd_sc_hd__xnor2_2 _25009_ (.A(_04355_),
    .B(_04358_),
    .Y(_04359_));
 sky130_fd_sc_hd__xnor2_1 _25010_ (.A(_04354_),
    .B(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__xnor2_1 _25011_ (.A(_04352_),
    .B(_04360_),
    .Y(_04361_));
 sky130_fd_sc_hd__a21bo_1 _25012_ (.A1(_04278_),
    .A2(_04283_),
    .B1_N(_04276_),
    .X(_04362_));
 sky130_fd_sc_hd__o21a_1 _25013_ (.A1(_04278_),
    .A2(_04283_),
    .B1(_04362_),
    .X(_04363_));
 sky130_fd_sc_hd__nor2_1 _25014_ (.A(_03325_),
    .B(_03743_),
    .Y(_04364_));
 sky130_fd_sc_hd__nor2_1 _25015_ (.A(_03112_),
    .B(_03900_),
    .Y(_04365_));
 sky130_fd_sc_hd__nor2_1 _25016_ (.A(_03254_),
    .B(_04288_),
    .Y(_04366_));
 sky130_fd_sc_hd__xnor2_1 _25017_ (.A(_04365_),
    .B(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__xnor2_2 _25018_ (.A(_04364_),
    .B(_04367_),
    .Y(_04368_));
 sky130_fd_sc_hd__a21o_1 _25019_ (.A1(_04279_),
    .A2(_04281_),
    .B1(_04280_),
    .X(_04369_));
 sky130_fd_sc_hd__o21a_1 _25020_ (.A1(_04279_),
    .A2(_04281_),
    .B1(_04369_),
    .X(_04370_));
 sky130_fd_sc_hd__clkbuf_4 _25021_ (.A(_03248_),
    .X(_04371_));
 sky130_fd_sc_hd__o211a_1 _25022_ (.A1(_04289_),
    .A2(_04291_),
    .B1(_04371_),
    .C1(_03758_),
    .X(_04372_));
 sky130_fd_sc_hd__a21o_1 _25023_ (.A1(_04289_),
    .A2(_04291_),
    .B1(_04372_),
    .X(_04373_));
 sky130_fd_sc_hd__xnor2_1 _25024_ (.A(_04370_),
    .B(_04373_),
    .Y(_04374_));
 sky130_fd_sc_hd__xnor2_2 _25025_ (.A(_04368_),
    .B(_04374_),
    .Y(_04375_));
 sky130_fd_sc_hd__xnor2_1 _25026_ (.A(_04363_),
    .B(_04375_),
    .Y(_04376_));
 sky130_fd_sc_hd__xnor2_1 _25027_ (.A(_04361_),
    .B(_04376_),
    .Y(_04377_));
 sky130_fd_sc_hd__a21bo_1 _25028_ (.A1(_04287_),
    .A2(_04299_),
    .B1_N(_04285_),
    .X(_04378_));
 sky130_fd_sc_hd__o21a_1 _25029_ (.A1(_04287_),
    .A2(_04299_),
    .B1(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__xor2_1 _25030_ (.A(_04377_),
    .B(_04379_),
    .X(_04380_));
 sky130_fd_sc_hd__xnor2_2 _25031_ (.A(_04347_),
    .B(_04380_),
    .Y(_04381_));
 sky130_fd_sc_hd__buf_4 _25032_ (.A(_04177_),
    .X(_04382_));
 sky130_fd_sc_hd__a21o_1 _25033_ (.A1(_04262_),
    .A2(_04266_),
    .B1(_04264_),
    .X(_04383_));
 sky130_fd_sc_hd__o21a_1 _25034_ (.A1(_04262_),
    .A2(_04266_),
    .B1(_04383_),
    .X(_04384_));
 sky130_fd_sc_hd__or2_1 _25035_ (.A(_04382_),
    .B(_04384_),
    .X(_04385_));
 sky130_fd_sc_hd__nand2_1 _25036_ (.A(_04382_),
    .B(_04384_),
    .Y(_04386_));
 sky130_fd_sc_hd__and2_1 _25037_ (.A(_04385_),
    .B(_04386_),
    .X(_04387_));
 sky130_fd_sc_hd__o21ba_1 _25038_ (.A1(_04268_),
    .A2(_04301_),
    .B1_N(_04270_),
    .X(_04388_));
 sky130_fd_sc_hd__a21o_1 _25039_ (.A1(_04268_),
    .A2(_04301_),
    .B1(_04388_),
    .X(_04389_));
 sky130_fd_sc_hd__xor2_1 _25040_ (.A(_04387_),
    .B(_04389_),
    .X(_04390_));
 sky130_fd_sc_hd__xnor2_2 _25041_ (.A(_04381_),
    .B(_04390_),
    .Y(_04391_));
 sky130_fd_sc_hd__or2_1 _25042_ (.A(_04305_),
    .B(_04312_),
    .X(_04392_));
 sky130_fd_sc_hd__nand2_1 _25043_ (.A(_04305_),
    .B(_04312_),
    .Y(_04393_));
 sky130_fd_sc_hd__nand2_1 _25044_ (.A(_04303_),
    .B(_04393_),
    .Y(_04394_));
 sky130_fd_sc_hd__nand2_1 _25045_ (.A(_04382_),
    .B(_04303_),
    .Y(_04395_));
 sky130_fd_sc_hd__nor2_1 _25046_ (.A(_04303_),
    .B(_04393_),
    .Y(_04396_));
 sky130_fd_sc_hd__o21bai_1 _25047_ (.A1(_04395_),
    .A2(_04392_),
    .B1_N(_04396_),
    .Y(_04397_));
 sky130_fd_sc_hd__a31o_1 _25048_ (.A1(_04306_),
    .A2(_04392_),
    .A3(_04394_),
    .B1(_04397_),
    .X(_04398_));
 sky130_fd_sc_hd__xor2_2 _25049_ (.A(_04391_),
    .B(_04398_),
    .X(_04399_));
 sky130_fd_sc_hd__xor2_1 _25050_ (.A(_04334_),
    .B(_04399_),
    .X(_04400_));
 sky130_fd_sc_hd__xnor2_1 _25051_ (.A(_04331_),
    .B(_04400_),
    .Y(_04401_));
 sky130_fd_sc_hd__mux2_1 _25052_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[8] ),
    .A1(_04401_),
    .S(_03642_),
    .X(_04402_));
 sky130_fd_sc_hd__clkbuf_1 _25053_ (.A(_04402_),
    .X(_00609_));
 sky130_fd_sc_hd__a221o_1 _25054_ (.A1(_04251_),
    .A2(_04325_),
    .B1(_04334_),
    .B2(_04399_),
    .C1(_04330_),
    .X(_04403_));
 sky130_fd_sc_hd__o21ai_1 _25055_ (.A1(_04334_),
    .A2(_04399_),
    .B1(_04403_),
    .Y(_04404_));
 sky130_fd_sc_hd__a21o_1 _25056_ (.A1(_04395_),
    .A2(_04391_),
    .B1(_04392_),
    .X(_04405_));
 sky130_fd_sc_hd__buf_4 _25057_ (.A(_04306_),
    .X(_04406_));
 sky130_fd_sc_hd__o21a_1 _25058_ (.A1(_04406_),
    .A2(_04396_),
    .B1(_04394_),
    .X(_04407_));
 sky130_fd_sc_hd__or2_1 _25059_ (.A(_04391_),
    .B(_04407_),
    .X(_04408_));
 sky130_fd_sc_hd__a21o_1 _25060_ (.A1(_04370_),
    .A2(_04373_),
    .B1(_04368_),
    .X(_04409_));
 sky130_fd_sc_hd__o21ai_2 _25061_ (.A1(_04370_),
    .A2(_04373_),
    .B1(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hd__and4_2 _25062_ (.A(_04252_),
    .B(_03305_),
    .C(_03829_),
    .D(_04258_),
    .X(_04411_));
 sky130_fd_sc_hd__nor2_1 _25063_ (.A(_03355_),
    .B(_04252_),
    .Y(_04412_));
 sky130_fd_sc_hd__and3_1 _25064_ (.A(_03355_),
    .B(_04252_),
    .C(_04131_),
    .X(_04413_));
 sky130_fd_sc_hd__mux2_1 _25065_ (.A0(_04412_),
    .A1(_04413_),
    .S(_04258_),
    .X(_04414_));
 sky130_fd_sc_hd__and3_1 _25066_ (.A(_03234_),
    .B(_03502_),
    .C(_04131_),
    .X(_04415_));
 sky130_fd_sc_hd__a31o_1 _25067_ (.A1(_04252_),
    .A2(_04258_),
    .A3(_04415_),
    .B1(_04039_),
    .X(_04416_));
 sky130_fd_sc_hd__a21o_1 _25068_ (.A1(_03765_),
    .A2(_04414_),
    .B1(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__nor2_1 _25069_ (.A(_04411_),
    .B(_04417_),
    .Y(_04418_));
 sky130_fd_sc_hd__xnor2_2 _25070_ (.A(_04410_),
    .B(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__nand2_1 _25071_ (.A(_03474_),
    .B(_03936_),
    .Y(_04420_));
 sky130_fd_sc_hd__nor2_1 _25072_ (.A(_03343_),
    .B(_04272_),
    .Y(_04421_));
 sky130_fd_sc_hd__nor2_1 _25073_ (.A(_02982_),
    .B(_04182_),
    .Y(_04422_));
 sky130_fd_sc_hd__xnor2_1 _25074_ (.A(_04421_),
    .B(_04422_),
    .Y(_04423_));
 sky130_fd_sc_hd__xnor2_1 _25075_ (.A(_04420_),
    .B(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__o21ai_1 _25076_ (.A1(_03474_),
    .A2(_04182_),
    .B1(_04348_),
    .Y(_04425_));
 sky130_fd_sc_hd__and3_1 _25077_ (.A(_03496_),
    .B(_03826_),
    .C(_04350_),
    .X(_04426_));
 sky130_fd_sc_hd__a21o_1 _25078_ (.A1(_04349_),
    .A2(_04425_),
    .B1(_04426_),
    .X(_04427_));
 sky130_fd_sc_hd__nor2_2 _25079_ (.A(net1017),
    .B(_04097_),
    .Y(_04428_));
 sky130_fd_sc_hd__nor2_1 _25080_ (.A(_03900_),
    .B(_03200_),
    .Y(_04429_));
 sky130_fd_sc_hd__nor2_1 _25081_ (.A(_03280_),
    .B(_04190_),
    .Y(_04430_));
 sky130_fd_sc_hd__xnor2_1 _25082_ (.A(_04429_),
    .B(_04430_),
    .Y(_04431_));
 sky130_fd_sc_hd__xnor2_2 _25083_ (.A(_04428_),
    .B(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__xnor2_1 _25084_ (.A(_04427_),
    .B(_04432_),
    .Y(_04433_));
 sky130_fd_sc_hd__xnor2_1 _25085_ (.A(_04424_),
    .B(_04433_),
    .Y(_04434_));
 sky130_fd_sc_hd__a21bo_1 _25086_ (.A1(_04354_),
    .A2(_04359_),
    .B1_N(_04352_),
    .X(_04435_));
 sky130_fd_sc_hd__o21a_1 _25087_ (.A1(_04354_),
    .A2(_04359_),
    .B1(_04435_),
    .X(_04436_));
 sky130_fd_sc_hd__nor2_2 _25088_ (.A(_03325_),
    .B(_03908_),
    .Y(_04437_));
 sky130_fd_sc_hd__nor2_1 _25089_ (.A(_03112_),
    .B(_04288_),
    .Y(_04438_));
 sky130_fd_sc_hd__nor2_1 _25090_ (.A(_03254_),
    .B(_03743_),
    .Y(_04439_));
 sky130_fd_sc_hd__xnor2_1 _25091_ (.A(_04438_),
    .B(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__xnor2_2 _25092_ (.A(_04437_),
    .B(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__a21o_1 _25093_ (.A1(_04355_),
    .A2(_04357_),
    .B1(_04356_),
    .X(_04442_));
 sky130_fd_sc_hd__o21a_1 _25094_ (.A1(_04355_),
    .A2(_04357_),
    .B1(_04442_),
    .X(_04443_));
 sky130_fd_sc_hd__a21o_1 _25095_ (.A1(_04364_),
    .A2(_04366_),
    .B1(_04365_),
    .X(_04444_));
 sky130_fd_sc_hd__o21a_1 _25096_ (.A1(_04364_),
    .A2(_04366_),
    .B1(_04444_),
    .X(_04445_));
 sky130_fd_sc_hd__xnor2_1 _25097_ (.A(_04443_),
    .B(_04445_),
    .Y(_04446_));
 sky130_fd_sc_hd__xnor2_2 _25098_ (.A(_04441_),
    .B(_04446_),
    .Y(_04447_));
 sky130_fd_sc_hd__xnor2_1 _25099_ (.A(_04436_),
    .B(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__xnor2_1 _25100_ (.A(_04434_),
    .B(_04448_),
    .Y(_04449_));
 sky130_fd_sc_hd__o21ba_1 _25101_ (.A1(_04363_),
    .A2(_04375_),
    .B1_N(_04361_),
    .X(_04450_));
 sky130_fd_sc_hd__a21oi_1 _25102_ (.A1(_04363_),
    .A2(_04375_),
    .B1(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__nor2_1 _25103_ (.A(_04449_),
    .B(_04451_),
    .Y(_04452_));
 sky130_fd_sc_hd__nand2_1 _25104_ (.A(_04449_),
    .B(_04451_),
    .Y(_04453_));
 sky130_fd_sc_hd__and2b_1 _25105_ (.A_N(_04452_),
    .B(_04453_),
    .X(_04454_));
 sky130_fd_sc_hd__xnor2_2 _25106_ (.A(_04419_),
    .B(_04454_),
    .Y(_04455_));
 sky130_fd_sc_hd__o21ba_1 _25107_ (.A1(_04347_),
    .A2(_04379_),
    .B1_N(_04377_),
    .X(_04456_));
 sky130_fd_sc_hd__a21oi_1 _25108_ (.A1(_04347_),
    .A2(_04379_),
    .B1(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__o21ba_1 _25109_ (.A1(_04336_),
    .A2(_04344_),
    .B1_N(_04345_),
    .X(_04458_));
 sky130_fd_sc_hd__xnor2_1 _25110_ (.A(_04382_),
    .B(_04458_),
    .Y(_04459_));
 sky130_fd_sc_hd__xnor2_1 _25111_ (.A(_04457_),
    .B(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__xnor2_1 _25112_ (.A(_04455_),
    .B(_04460_),
    .Y(_04461_));
 sky130_fd_sc_hd__a21o_1 _25113_ (.A1(_04387_),
    .A2(_04389_),
    .B1(_04381_),
    .X(_04462_));
 sky130_fd_sc_hd__o21a_1 _25114_ (.A1(_04387_),
    .A2(_04389_),
    .B1(_04462_),
    .X(_04463_));
 sky130_fd_sc_hd__xnor2_1 _25115_ (.A(_04386_),
    .B(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__xnor2_1 _25116_ (.A(_04461_),
    .B(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__a21o_1 _25117_ (.A1(_04405_),
    .A2(_04408_),
    .B1(_04465_),
    .X(_04466_));
 sky130_fd_sc_hd__inv_2 _25118_ (.A(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__and3_1 _25119_ (.A(_04405_),
    .B(_04408_),
    .C(_04465_),
    .X(_04468_));
 sky130_fd_sc_hd__nor2_1 _25120_ (.A(_04467_),
    .B(_04468_),
    .Y(_04469_));
 sky130_fd_sc_hd__xnor2_1 _25121_ (.A(_04404_),
    .B(_04469_),
    .Y(_04470_));
 sky130_fd_sc_hd__mux2_1 _25122_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[9] ),
    .A1(_04470_),
    .S(_03642_),
    .X(_04471_));
 sky130_fd_sc_hd__clkbuf_1 _25123_ (.A(_04471_),
    .X(_00610_));
 sky130_fd_sc_hd__o21a_1 _25124_ (.A1(_04387_),
    .A2(_04389_),
    .B1(_04381_),
    .X(_04472_));
 sky130_fd_sc_hd__nand2_1 _25125_ (.A(_04461_),
    .B(_04463_),
    .Y(_04473_));
 sky130_fd_sc_hd__a2bb2o_1 _25126_ (.A1_N(_04461_),
    .A2_N(_04472_),
    .B1(_04473_),
    .B2(_04386_),
    .X(_04474_));
 sky130_fd_sc_hd__o21a_2 _25127_ (.A1(_04419_),
    .A2(_04452_),
    .B1(_04453_),
    .X(_04475_));
 sky130_fd_sc_hd__nand2_1 _25128_ (.A(_02982_),
    .B(_03936_),
    .Y(_04476_));
 sky130_fd_sc_hd__nor2_1 _25129_ (.A(net1017),
    .B(_04272_),
    .Y(_04477_));
 sky130_fd_sc_hd__nor2_1 _25130_ (.A(_03343_),
    .B(_04182_),
    .Y(_04478_));
 sky130_fd_sc_hd__xnor2_1 _25131_ (.A(_04477_),
    .B(_04478_),
    .Y(_04479_));
 sky130_fd_sc_hd__xnor2_2 _25132_ (.A(_04476_),
    .B(_04479_),
    .Y(_04480_));
 sky130_fd_sc_hd__o21ai_1 _25133_ (.A1(_03343_),
    .A2(_04272_),
    .B1(_04420_),
    .Y(_04481_));
 sky130_fd_sc_hd__and3_1 _25134_ (.A(_03474_),
    .B(_03936_),
    .C(_04421_),
    .X(_04482_));
 sky130_fd_sc_hd__a21o_1 _25135_ (.A1(_04422_),
    .A2(_04481_),
    .B1(_04482_),
    .X(_04483_));
 sky130_fd_sc_hd__nor2_1 _25136_ (.A(_03200_),
    .B(_04288_),
    .Y(_04484_));
 sky130_fd_sc_hd__o211a_1 _25137_ (.A1(_03280_),
    .A2(_04097_),
    .B1(_03123_),
    .C1(_03981_),
    .X(_04485_));
 sky130_fd_sc_hd__o211a_1 _25138_ (.A1(_03900_),
    .A2(_04190_),
    .B1(_03889_),
    .C1(_03758_),
    .X(_04486_));
 sky130_fd_sc_hd__nor2_1 _25139_ (.A(_04485_),
    .B(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__xnor2_2 _25140_ (.A(_04484_),
    .B(_04487_),
    .Y(_04488_));
 sky130_fd_sc_hd__xnor2_1 _25141_ (.A(_04483_),
    .B(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__xnor2_2 _25142_ (.A(_04480_),
    .B(_04489_),
    .Y(_04490_));
 sky130_fd_sc_hd__a21bo_1 _25143_ (.A1(_04427_),
    .A2(_04432_),
    .B1_N(_04424_),
    .X(_04491_));
 sky130_fd_sc_hd__o21ai_2 _25144_ (.A1(_04427_),
    .A2(_04432_),
    .B1(_04491_),
    .Y(_04492_));
 sky130_fd_sc_hd__xnor2_1 _25145_ (.A(_03325_),
    .B(_03254_),
    .Y(_04493_));
 sky130_fd_sc_hd__o211a_1 _25146_ (.A1(_04039_),
    .A2(_04493_),
    .B1(_04371_),
    .C1(_04174_),
    .X(_04494_));
 sky130_fd_sc_hd__a211o_1 _25147_ (.A1(_04371_),
    .A2(_04174_),
    .B1(_04039_),
    .C1(_04493_),
    .X(_04495_));
 sky130_fd_sc_hd__and2b_1 _25148_ (.A_N(_04494_),
    .B(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__a21o_1 _25149_ (.A1(_04428_),
    .A2(_04430_),
    .B1(_04429_),
    .X(_04497_));
 sky130_fd_sc_hd__o21a_1 _25150_ (.A1(_04428_),
    .A2(_04430_),
    .B1(_04497_),
    .X(_04498_));
 sky130_fd_sc_hd__o211a_1 _25151_ (.A1(_04437_),
    .A2(_04439_),
    .B1(_04371_),
    .C1(_03687_),
    .X(_04499_));
 sky130_fd_sc_hd__a21o_1 _25152_ (.A1(_04437_),
    .A2(_04439_),
    .B1(_04499_),
    .X(_04500_));
 sky130_fd_sc_hd__nor2_1 _25153_ (.A(_04498_),
    .B(_04500_),
    .Y(_04501_));
 sky130_fd_sc_hd__nand2_1 _25154_ (.A(_04498_),
    .B(_04500_),
    .Y(_04502_));
 sky130_fd_sc_hd__or2b_1 _25155_ (.A(_04501_),
    .B_N(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__xnor2_2 _25156_ (.A(_04496_),
    .B(_04503_),
    .Y(_04504_));
 sky130_fd_sc_hd__xnor2_1 _25157_ (.A(_04492_),
    .B(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__xnor2_2 _25158_ (.A(_04490_),
    .B(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__a21bo_1 _25159_ (.A1(_04436_),
    .A2(_04447_),
    .B1_N(_04434_),
    .X(_04507_));
 sky130_fd_sc_hd__o21a_1 _25160_ (.A1(_04436_),
    .A2(_04447_),
    .B1(_04507_),
    .X(_04508_));
 sky130_fd_sc_hd__a31o_2 _25161_ (.A1(_03355_),
    .A2(_04252_),
    .A3(_03502_),
    .B1(_04339_),
    .X(_04509_));
 sky130_fd_sc_hd__xnor2_4 _25162_ (.A(_04069_),
    .B(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__a21o_1 _25163_ (.A1(_04443_),
    .A2(_04445_),
    .B1(_04441_),
    .X(_04511_));
 sky130_fd_sc_hd__o21ai_2 _25164_ (.A1(_04443_),
    .A2(_04445_),
    .B1(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hd__xnor2_1 _25165_ (.A(_04510_),
    .B(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__xnor2_1 _25166_ (.A(_04508_),
    .B(_04513_),
    .Y(_04514_));
 sky130_fd_sc_hd__xnor2_2 _25167_ (.A(_04506_),
    .B(_04514_),
    .Y(_04515_));
 sky130_fd_sc_hd__or4b_4 _25168_ (.A(_03007_),
    .B(_04039_),
    .C(_04067_),
    .D_N(_03305_),
    .X(_04516_));
 sky130_fd_sc_hd__a21oi_2 _25169_ (.A1(_04410_),
    .A2(_04516_),
    .B1(_04417_),
    .Y(_04517_));
 sky130_fd_sc_hd__buf_4 _25170_ (.A(_04039_),
    .X(_04518_));
 sky130_fd_sc_hd__a21oi_1 _25171_ (.A1(_03355_),
    .A2(_04252_),
    .B1(_04258_),
    .Y(_04519_));
 sky130_fd_sc_hd__o22a_1 _25172_ (.A1(_04069_),
    .A2(_04412_),
    .B1(_04519_),
    .B2(_03765_),
    .X(_04520_));
 sky130_fd_sc_hd__nor2_4 _25173_ (.A(_04518_),
    .B(_04520_),
    .Y(_04521_));
 sky130_fd_sc_hd__xnor2_4 _25174_ (.A(_04177_),
    .B(_04521_),
    .Y(_04522_));
 sky130_fd_sc_hd__xnor2_1 _25175_ (.A(_04517_),
    .B(_04522_),
    .Y(_04523_));
 sky130_fd_sc_hd__xnor2_1 _25176_ (.A(_04515_),
    .B(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__xnor2_2 _25177_ (.A(_04475_),
    .B(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__and2_1 _25178_ (.A(_04457_),
    .B(_04458_),
    .X(_04526_));
 sky130_fd_sc_hd__or2_1 _25179_ (.A(_04457_),
    .B(_04458_),
    .X(_04527_));
 sky130_fd_sc_hd__o21ai_1 _25180_ (.A1(_04455_),
    .A2(_04526_),
    .B1(_04527_),
    .Y(_04528_));
 sky130_fd_sc_hd__or3_1 _25181_ (.A(_04306_),
    .B(_04455_),
    .C(_04527_),
    .X(_04529_));
 sky130_fd_sc_hd__nand2_1 _25182_ (.A(_04455_),
    .B(_04526_),
    .Y(_04530_));
 sky130_fd_sc_hd__o211a_1 _25183_ (.A1(_04382_),
    .A2(_04528_),
    .B1(_04529_),
    .C1(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__xnor2_1 _25184_ (.A(_04525_),
    .B(_04531_),
    .Y(_04532_));
 sky130_fd_sc_hd__xor2_1 _25185_ (.A(_04474_),
    .B(_04532_),
    .X(_04533_));
 sky130_fd_sc_hd__a21o_1 _25186_ (.A1(_04404_),
    .A2(_04466_),
    .B1(_04468_),
    .X(_04534_));
 sky130_fd_sc_hd__xnor2_1 _25187_ (.A(_04533_),
    .B(_04534_),
    .Y(_04535_));
 sky130_fd_sc_hd__mux2_1 _25188_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[10] ),
    .A1(_04535_),
    .S(_03146_),
    .X(_04536_));
 sky130_fd_sc_hd__clkbuf_1 _25189_ (.A(_04536_),
    .X(_00611_));
 sky130_fd_sc_hd__and2_1 _25190_ (.A(_04474_),
    .B(_04532_),
    .X(_04537_));
 sky130_fd_sc_hd__or2_1 _25191_ (.A(_04474_),
    .B(_04532_),
    .X(_04538_));
 sky130_fd_sc_hd__o21a_1 _25192_ (.A1(_04534_),
    .A2(_04537_),
    .B1(_04538_),
    .X(_04539_));
 sky130_fd_sc_hd__nor2_1 _25193_ (.A(_03200_),
    .B(_04131_),
    .Y(_04540_));
 sky130_fd_sc_hd__nor2_1 _25194_ (.A(_03900_),
    .B(_04097_),
    .Y(_04541_));
 sky130_fd_sc_hd__nor2_1 _25195_ (.A(_04190_),
    .B(_04288_),
    .Y(_04542_));
 sky130_fd_sc_hd__xor2_1 _25196_ (.A(_04541_),
    .B(_04542_),
    .X(_04543_));
 sky130_fd_sc_hd__xnor2_2 _25197_ (.A(_04540_),
    .B(_04543_),
    .Y(_04544_));
 sky130_fd_sc_hd__a21bo_1 _25198_ (.A1(_04477_),
    .A2(_04478_),
    .B1_N(_04476_),
    .X(_04545_));
 sky130_fd_sc_hd__o21a_1 _25199_ (.A1(_04477_),
    .A2(_04478_),
    .B1(_04545_),
    .X(_04546_));
 sky130_fd_sc_hd__nand2_1 _25200_ (.A(_03343_),
    .B(_03936_),
    .Y(_04547_));
 sky130_fd_sc_hd__nor2_1 _25201_ (.A(_03280_),
    .B(_04272_),
    .Y(_04548_));
 sky130_fd_sc_hd__nor2_1 _25202_ (.A(net1017),
    .B(_04182_),
    .Y(_04549_));
 sky130_fd_sc_hd__xor2_1 _25203_ (.A(_04548_),
    .B(_04549_),
    .X(_04550_));
 sky130_fd_sc_hd__xnor2_2 _25204_ (.A(_04547_),
    .B(_04550_),
    .Y(_04551_));
 sky130_fd_sc_hd__xnor2_1 _25205_ (.A(_04546_),
    .B(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__xnor2_2 _25206_ (.A(_04544_),
    .B(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__a21bo_1 _25207_ (.A1(_04483_),
    .A2(_04488_),
    .B1_N(_04480_),
    .X(_04554_));
 sky130_fd_sc_hd__o21ai_1 _25208_ (.A1(_04483_),
    .A2(_04488_),
    .B1(_04554_),
    .Y(_04555_));
 sky130_fd_sc_hd__a22o_1 _25209_ (.A1(_03981_),
    .A2(_03123_),
    .B1(_03889_),
    .B2(_03758_),
    .X(_04556_));
 sky130_fd_sc_hd__and4_1 _25210_ (.A(_03758_),
    .B(_03981_),
    .C(_03123_),
    .D(_03889_),
    .X(_04557_));
 sky130_fd_sc_hd__a21o_1 _25211_ (.A1(_04484_),
    .A2(_04556_),
    .B1(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__a21oi_1 _25212_ (.A1(_03254_),
    .A2(_04174_),
    .B1(_03325_),
    .Y(_04559_));
 sky130_fd_sc_hd__a21o_1 _25213_ (.A1(_03363_),
    .A2(_04131_),
    .B1(_04559_),
    .X(_04560_));
 sky130_fd_sc_hd__nand2_2 _25214_ (.A(_03325_),
    .B(_03254_),
    .Y(_04561_));
 sky130_fd_sc_hd__nor2_1 _25215_ (.A(_04371_),
    .B(_04561_),
    .Y(_04562_));
 sky130_fd_sc_hd__a211o_1 _25216_ (.A1(_04371_),
    .A2(_04560_),
    .B1(_04562_),
    .C1(_04518_),
    .X(_04563_));
 sky130_fd_sc_hd__xor2_1 _25217_ (.A(_04558_),
    .B(_04563_),
    .X(_04564_));
 sky130_fd_sc_hd__and2_1 _25218_ (.A(_04555_),
    .B(_04564_),
    .X(_04565_));
 sky130_fd_sc_hd__or2_1 _25219_ (.A(_04555_),
    .B(_04564_),
    .X(_04566_));
 sky130_fd_sc_hd__and2b_1 _25220_ (.A_N(_04565_),
    .B(_04566_),
    .X(_04567_));
 sky130_fd_sc_hd__xor2_2 _25221_ (.A(_04553_),
    .B(_04567_),
    .X(_04568_));
 sky130_fd_sc_hd__a21o_1 _25222_ (.A1(_04492_),
    .A2(_04504_),
    .B1(_04490_),
    .X(_04569_));
 sky130_fd_sc_hd__o21a_1 _25223_ (.A1(_04492_),
    .A2(_04504_),
    .B1(_04569_),
    .X(_04570_));
 sky130_fd_sc_hd__and2_2 _25224_ (.A(_04069_),
    .B(_04339_),
    .X(_04571_));
 sky130_fd_sc_hd__nor2_4 _25225_ (.A(_04411_),
    .B(_04571_),
    .Y(_04572_));
 sky130_fd_sc_hd__a21oi_2 _25226_ (.A1(_04496_),
    .A2(_04502_),
    .B1(_04501_),
    .Y(_04573_));
 sky130_fd_sc_hd__xnor2_2 _25227_ (.A(_04572_),
    .B(_04573_),
    .Y(_04574_));
 sky130_fd_sc_hd__xnor2_1 _25228_ (.A(_04570_),
    .B(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__xnor2_1 _25229_ (.A(_04568_),
    .B(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hd__xnor2_1 _25230_ (.A(_04512_),
    .B(_04572_),
    .Y(_04577_));
 sky130_fd_sc_hd__o21ba_1 _25231_ (.A1(_04508_),
    .A2(_04577_),
    .B1_N(_04506_),
    .X(_04578_));
 sky130_fd_sc_hd__a21oi_1 _25232_ (.A1(_04508_),
    .A2(_04577_),
    .B1(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__a21oi_2 _25233_ (.A1(_04516_),
    .A2(_04512_),
    .B1(_04571_),
    .Y(_04580_));
 sky130_fd_sc_hd__xnor2_1 _25234_ (.A(_04382_),
    .B(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__and2_1 _25235_ (.A(_04579_),
    .B(_04581_),
    .X(_04582_));
 sky130_fd_sc_hd__or2_1 _25236_ (.A(_04579_),
    .B(_04581_),
    .X(_04583_));
 sky130_fd_sc_hd__and2b_1 _25237_ (.A_N(_04582_),
    .B(_04583_),
    .X(_04584_));
 sky130_fd_sc_hd__xnor2_1 _25238_ (.A(_04576_),
    .B(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__inv_2 _25239_ (.A(_04585_),
    .Y(_04586_));
 sky130_fd_sc_hd__xor2_1 _25240_ (.A(_04515_),
    .B(_04521_),
    .X(_04587_));
 sky130_fd_sc_hd__nor2_1 _25241_ (.A(_04517_),
    .B(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hd__a21oi_1 _25242_ (.A1(_04517_),
    .A2(_04587_),
    .B1(_04475_),
    .Y(_04589_));
 sky130_fd_sc_hd__or2_1 _25243_ (.A(_04588_),
    .B(_04589_),
    .X(_04590_));
 sky130_fd_sc_hd__or2_1 _25244_ (.A(_04475_),
    .B(_04588_),
    .X(_04591_));
 sky130_fd_sc_hd__nand2_1 _25245_ (.A(_04517_),
    .B(_04587_),
    .Y(_04592_));
 sky130_fd_sc_hd__o21ai_1 _25246_ (.A1(_04406_),
    .A2(_04592_),
    .B1(_04475_),
    .Y(_04593_));
 sky130_fd_sc_hd__a22o_1 _25247_ (.A1(_04406_),
    .A2(_04590_),
    .B1(_04591_),
    .B2(_04593_),
    .X(_04594_));
 sky130_fd_sc_hd__xnor2_1 _25248_ (.A(_04586_),
    .B(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__nand2_1 _25249_ (.A(_04525_),
    .B(_04528_),
    .Y(_04596_));
 sky130_fd_sc_hd__inv_2 _25250_ (.A(_04525_),
    .Y(_04597_));
 sky130_fd_sc_hd__a21o_1 _25251_ (.A1(_04597_),
    .A2(_04527_),
    .B1(_04455_),
    .X(_04598_));
 sky130_fd_sc_hd__o21a_1 _25252_ (.A1(_04597_),
    .A2(_04526_),
    .B1(_04598_),
    .X(_04599_));
 sky130_fd_sc_hd__or2_1 _25253_ (.A(_04406_),
    .B(_04599_),
    .X(_04600_));
 sky130_fd_sc_hd__and3_1 _25254_ (.A(_04595_),
    .B(_04596_),
    .C(_04600_),
    .X(_04601_));
 sky130_fd_sc_hd__a21o_1 _25255_ (.A1(_04596_),
    .A2(_04600_),
    .B1(_04595_),
    .X(_04602_));
 sky130_fd_sc_hd__and2b_1 _25256_ (.A_N(_04601_),
    .B(_04602_),
    .X(_04603_));
 sky130_fd_sc_hd__xnor2_1 _25257_ (.A(_04539_),
    .B(_04603_),
    .Y(_04604_));
 sky130_fd_sc_hd__mux2_1 _25258_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[11] ),
    .A1(_04604_),
    .S(_03146_),
    .X(_04605_));
 sky130_fd_sc_hd__clkbuf_1 _25259_ (.A(_04605_),
    .X(_00612_));
 sky130_fd_sc_hd__a21o_1 _25260_ (.A1(_04537_),
    .A2(_04602_),
    .B1(_04601_),
    .X(_04606_));
 sky130_fd_sc_hd__a31o_1 _25261_ (.A1(_04534_),
    .A2(_04538_),
    .A3(_04602_),
    .B1(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__nand2_1 _25262_ (.A(_04586_),
    .B(_04592_),
    .Y(_04608_));
 sky130_fd_sc_hd__o2bb2a_1 _25263_ (.A1_N(_04475_),
    .A2_N(_04608_),
    .B1(_04588_),
    .B2(_04586_),
    .X(_04609_));
 sky130_fd_sc_hd__o22a_1 _25264_ (.A1(_04586_),
    .A2(_04590_),
    .B1(_04609_),
    .B2(_04406_),
    .X(_04610_));
 sky130_fd_sc_hd__a21o_1 _25265_ (.A1(_04570_),
    .A2(_04574_),
    .B1(_04568_),
    .X(_04611_));
 sky130_fd_sc_hd__o21ai_2 _25266_ (.A1(_04570_),
    .A2(_04574_),
    .B1(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hd__nor2_2 _25267_ (.A(_03200_),
    .B(_04518_),
    .Y(_04613_));
 sky130_fd_sc_hd__nor2_2 _25268_ (.A(_04097_),
    .B(_04288_),
    .Y(_04614_));
 sky130_fd_sc_hd__nor2_2 _25269_ (.A(_04190_),
    .B(_04131_),
    .Y(_04615_));
 sky130_fd_sc_hd__xnor2_2 _25270_ (.A(_04614_),
    .B(_04615_),
    .Y(_04616_));
 sky130_fd_sc_hd__xnor2_4 _25271_ (.A(_04613_),
    .B(_04616_),
    .Y(_04617_));
 sky130_fd_sc_hd__a21bo_1 _25272_ (.A1(_04548_),
    .A2(_04549_),
    .B1_N(_04547_),
    .X(_04618_));
 sky130_fd_sc_hd__o21a_1 _25273_ (.A1(_04548_),
    .A2(_04549_),
    .B1(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__nand2_1 _25274_ (.A(net1017),
    .B(_03936_),
    .Y(_04620_));
 sky130_fd_sc_hd__nor2_1 _25275_ (.A(_03900_),
    .B(_04272_),
    .Y(_04621_));
 sky130_fd_sc_hd__nor2_1 _25276_ (.A(_03280_),
    .B(_04182_),
    .Y(_04622_));
 sky130_fd_sc_hd__xor2_1 _25277_ (.A(_04621_),
    .B(_04622_),
    .X(_04623_));
 sky130_fd_sc_hd__xnor2_2 _25278_ (.A(_04620_),
    .B(_04623_),
    .Y(_04624_));
 sky130_fd_sc_hd__xor2_2 _25279_ (.A(_04619_),
    .B(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__xnor2_4 _25280_ (.A(_04617_),
    .B(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__a21bo_1 _25281_ (.A1(_04546_),
    .A2(_04551_),
    .B1_N(_04544_),
    .X(_04627_));
 sky130_fd_sc_hd__o21a_1 _25282_ (.A1(_04546_),
    .A2(_04551_),
    .B1(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__a21o_1 _25283_ (.A1(_04541_),
    .A2(_04542_),
    .B1(_04540_),
    .X(_04629_));
 sky130_fd_sc_hd__o21a_1 _25284_ (.A1(_04541_),
    .A2(_04542_),
    .B1(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__and3_1 _25285_ (.A(_04371_),
    .B(_03056_),
    .C(_03363_),
    .X(_04631_));
 sky130_fd_sc_hd__or3_1 _25286_ (.A(_04039_),
    .B(_04562_),
    .C(_04631_),
    .X(_04632_));
 sky130_fd_sc_hd__clkbuf_2 _25287_ (.A(_04632_),
    .X(_04633_));
 sky130_fd_sc_hd__xor2_1 _25288_ (.A(_04630_),
    .B(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__and2b_1 _25289_ (.A_N(_04628_),
    .B(_04634_),
    .X(_04635_));
 sky130_fd_sc_hd__or2b_1 _25290_ (.A(_04634_),
    .B_N(_04628_),
    .X(_04636_));
 sky130_fd_sc_hd__or2b_2 _25291_ (.A(_04635_),
    .B_N(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__xnor2_4 _25292_ (.A(_04626_),
    .B(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__a21o_1 _25293_ (.A1(_04553_),
    .A2(_04566_),
    .B1(_04565_),
    .X(_04639_));
 sky130_fd_sc_hd__or3b_1 _25294_ (.A(_03112_),
    .B(_04174_),
    .C_N(_04561_),
    .X(_04640_));
 sky130_fd_sc_hd__and3b_1 _25295_ (.A_N(_04562_),
    .B(_04640_),
    .C(_04558_),
    .X(_04641_));
 sky130_fd_sc_hd__o21ai_2 _25296_ (.A1(_04631_),
    .A2(_04641_),
    .B1(_03829_),
    .Y(_04642_));
 sky130_fd_sc_hd__xor2_2 _25297_ (.A(_04510_),
    .B(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__xor2_1 _25298_ (.A(_04639_),
    .B(_04643_),
    .X(_04644_));
 sky130_fd_sc_hd__xnor2_2 _25299_ (.A(_04638_),
    .B(_04644_),
    .Y(_04645_));
 sky130_fd_sc_hd__nand2_1 _25300_ (.A(_04069_),
    .B(_04339_),
    .Y(_04646_));
 sky130_fd_sc_hd__o21a_1 _25301_ (.A1(_04411_),
    .A2(_04573_),
    .B1(_04646_),
    .X(_04647_));
 sky130_fd_sc_hd__xnor2_1 _25302_ (.A(_04522_),
    .B(_04647_),
    .Y(_04648_));
 sky130_fd_sc_hd__xnor2_1 _25303_ (.A(_04645_),
    .B(_04648_),
    .Y(_04649_));
 sky130_fd_sc_hd__xnor2_1 _25304_ (.A(_04612_),
    .B(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__o21a_1 _25305_ (.A1(_04576_),
    .A2(_04582_),
    .B1(_04583_),
    .X(_04651_));
 sky130_fd_sc_hd__nand2_1 _25306_ (.A(_04382_),
    .B(_04580_),
    .Y(_04652_));
 sky130_fd_sc_hd__xnor2_1 _25307_ (.A(_04651_),
    .B(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__xnor2_1 _25308_ (.A(_04650_),
    .B(_04653_),
    .Y(_04654_));
 sky130_fd_sc_hd__or2_1 _25309_ (.A(_04610_),
    .B(_04654_),
    .X(_04655_));
 sky130_fd_sc_hd__and2_1 _25310_ (.A(_04610_),
    .B(_04654_),
    .X(_04656_));
 sky130_fd_sc_hd__inv_2 _25311_ (.A(_04656_),
    .Y(_04657_));
 sky130_fd_sc_hd__nand2_1 _25312_ (.A(_04655_),
    .B(_04657_),
    .Y(_04658_));
 sky130_fd_sc_hd__xor2_1 _25313_ (.A(_04607_),
    .B(_04658_),
    .X(_04659_));
 sky130_fd_sc_hd__mux2_1 _25314_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[12] ),
    .A1(_04659_),
    .S(_03146_),
    .X(_04660_));
 sky130_fd_sc_hd__clkbuf_1 _25315_ (.A(_04660_),
    .X(_00613_));
 sky130_fd_sc_hd__o21a_2 _25316_ (.A1(_04607_),
    .A2(_04656_),
    .B1(_04655_),
    .X(_04661_));
 sky130_fd_sc_hd__o21a_1 _25317_ (.A1(_04651_),
    .A2(_04652_),
    .B1(_04650_),
    .X(_04662_));
 sky130_fd_sc_hd__a21oi_2 _25318_ (.A1(_04651_),
    .A2(_04652_),
    .B1(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__nand2_2 _25319_ (.A(_04382_),
    .B(_04647_),
    .Y(_04664_));
 sky130_fd_sc_hd__and2_1 _25320_ (.A(_04521_),
    .B(_04643_),
    .X(_04665_));
 sky130_fd_sc_hd__nor2_1 _25321_ (.A(_04521_),
    .B(_04643_),
    .Y(_04666_));
 sky130_fd_sc_hd__o22a_1 _25322_ (.A1(_04639_),
    .A2(_04638_),
    .B1(_04665_),
    .B2(_04666_),
    .X(_04667_));
 sky130_fd_sc_hd__a21oi_2 _25323_ (.A1(_04639_),
    .A2(_04638_),
    .B1(_04667_),
    .Y(_04668_));
 sky130_fd_sc_hd__nand2_1 _25324_ (.A(_03280_),
    .B(_03936_),
    .Y(_04669_));
 sky130_fd_sc_hd__nor2_1 _25325_ (.A(_04272_),
    .B(_04288_),
    .Y(_04670_));
 sky130_fd_sc_hd__nor2_1 _25326_ (.A(_03900_),
    .B(_04182_),
    .Y(_04671_));
 sky130_fd_sc_hd__xnor2_1 _25327_ (.A(_04670_),
    .B(_04671_),
    .Y(_04672_));
 sky130_fd_sc_hd__xnor2_2 _25328_ (.A(_04669_),
    .B(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__o21ba_1 _25329_ (.A1(_04621_),
    .A2(_04622_),
    .B1_N(_04620_),
    .X(_04674_));
 sky130_fd_sc_hd__a21oi_1 _25330_ (.A1(_04621_),
    .A2(_04622_),
    .B1(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__nor2_1 _25331_ (.A(_04097_),
    .B(_04131_),
    .Y(_04676_));
 sky130_fd_sc_hd__xnor2_1 _25332_ (.A(_03123_),
    .B(_03200_),
    .Y(_04677_));
 sky130_fd_sc_hd__nand2_1 _25333_ (.A(_03829_),
    .B(_04677_),
    .Y(_04678_));
 sky130_fd_sc_hd__xor2_1 _25334_ (.A(_04676_),
    .B(_04678_),
    .X(_04679_));
 sky130_fd_sc_hd__and2_1 _25335_ (.A(_04675_),
    .B(_04679_),
    .X(_04680_));
 sky130_fd_sc_hd__or2_1 _25336_ (.A(_04675_),
    .B(_04679_),
    .X(_04681_));
 sky130_fd_sc_hd__and2b_1 _25337_ (.A_N(_04680_),
    .B(_04681_),
    .X(_04682_));
 sky130_fd_sc_hd__xnor2_2 _25338_ (.A(_04673_),
    .B(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__a21o_1 _25339_ (.A1(_04619_),
    .A2(_04624_),
    .B1(_04617_),
    .X(_04684_));
 sky130_fd_sc_hd__o21a_1 _25340_ (.A1(_04619_),
    .A2(_04624_),
    .B1(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__a21oi_1 _25341_ (.A1(_04614_),
    .A2(_04615_),
    .B1(_04613_),
    .Y(_04686_));
 sky130_fd_sc_hd__o21ba_1 _25342_ (.A1(_04614_),
    .A2(_04615_),
    .B1_N(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__xnor2_1 _25343_ (.A(_04633_),
    .B(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__xor2_1 _25344_ (.A(_04685_),
    .B(_04688_),
    .X(_04689_));
 sky130_fd_sc_hd__xnor2_2 _25345_ (.A(_04683_),
    .B(_04689_),
    .Y(_04690_));
 sky130_fd_sc_hd__a21o_1 _25346_ (.A1(_04626_),
    .A2(_04636_),
    .B1(_04635_),
    .X(_04691_));
 sky130_fd_sc_hd__o21ai_1 _25347_ (.A1(_03326_),
    .A2(_04630_),
    .B1(_04371_),
    .Y(_04692_));
 sky130_fd_sc_hd__nand2_1 _25348_ (.A(_04561_),
    .B(_04630_),
    .Y(_04693_));
 sky130_fd_sc_hd__a21oi_2 _25349_ (.A1(_04692_),
    .A2(_04693_),
    .B1(_04518_),
    .Y(_04694_));
 sky130_fd_sc_hd__xnor2_1 _25350_ (.A(_04510_),
    .B(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__xnor2_1 _25351_ (.A(_04691_),
    .B(_04695_),
    .Y(_04696_));
 sky130_fd_sc_hd__xnor2_2 _25352_ (.A(_04690_),
    .B(_04696_),
    .Y(_04697_));
 sky130_fd_sc_hd__a21o_1 _25353_ (.A1(_04516_),
    .A2(_04642_),
    .B1(_04571_),
    .X(_04698_));
 sky130_fd_sc_hd__xor2_1 _25354_ (.A(_04522_),
    .B(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__xnor2_1 _25355_ (.A(_04697_),
    .B(_04699_),
    .Y(_04700_));
 sky130_fd_sc_hd__xnor2_2 _25356_ (.A(_04668_),
    .B(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__xnor2_1 _25357_ (.A(_04664_),
    .B(_04701_),
    .Y(_04702_));
 sky130_fd_sc_hd__or2_1 _25358_ (.A(_04382_),
    .B(_04647_),
    .X(_04703_));
 sky130_fd_sc_hd__xnor2_1 _25359_ (.A(_04521_),
    .B(_04645_),
    .Y(_04704_));
 sky130_fd_sc_hd__or2_1 _25360_ (.A(_04612_),
    .B(_04704_),
    .X(_04705_));
 sky130_fd_sc_hd__and2_1 _25361_ (.A(_04612_),
    .B(_04704_),
    .X(_04706_));
 sky130_fd_sc_hd__a31o_1 _25362_ (.A1(_04664_),
    .A2(_04703_),
    .A3(_04705_),
    .B1(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__xnor2_1 _25363_ (.A(_04702_),
    .B(_04707_),
    .Y(_04708_));
 sky130_fd_sc_hd__xnor2_1 _25364_ (.A(_04663_),
    .B(_04708_),
    .Y(_04709_));
 sky130_fd_sc_hd__xnor2_1 _25365_ (.A(_04661_),
    .B(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__mux2_1 _25366_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[13] ),
    .A1(_04710_),
    .S(_03146_),
    .X(_04711_));
 sky130_fd_sc_hd__clkbuf_1 _25367_ (.A(_04711_),
    .X(_00614_));
 sky130_fd_sc_hd__nor2_2 _25368_ (.A(_04406_),
    .B(_04698_),
    .Y(_04712_));
 sky130_fd_sc_hd__and2_1 _25369_ (.A(_04406_),
    .B(_04698_),
    .X(_04713_));
 sky130_fd_sc_hd__xor2_1 _25370_ (.A(_04521_),
    .B(_04697_),
    .X(_04714_));
 sky130_fd_sc_hd__nor2_1 _25371_ (.A(_04668_),
    .B(_04714_),
    .Y(_04715_));
 sky130_fd_sc_hd__nand2_1 _25372_ (.A(_04668_),
    .B(_04714_),
    .Y(_04716_));
 sky130_fd_sc_hd__o31ai_4 _25373_ (.A1(_04712_),
    .A2(_04713_),
    .A3(_04715_),
    .B1(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__and2_1 _25374_ (.A(_04572_),
    .B(_04694_),
    .X(_04718_));
 sky130_fd_sc_hd__nor2_1 _25375_ (.A(_04572_),
    .B(_04694_),
    .Y(_04719_));
 sky130_fd_sc_hd__o22a_1 _25376_ (.A1(_04691_),
    .A2(_04690_),
    .B1(_04718_),
    .B2(_04719_),
    .X(_04720_));
 sky130_fd_sc_hd__a21o_1 _25377_ (.A1(_04691_),
    .A2(_04690_),
    .B1(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__nand2_2 _25378_ (.A(_03900_),
    .B(_03936_),
    .Y(_04722_));
 sky130_fd_sc_hd__nor2_2 _25379_ (.A(_04272_),
    .B(_04131_),
    .Y(_04723_));
 sky130_fd_sc_hd__nor2_1 _25380_ (.A(_04288_),
    .B(_04182_),
    .Y(_04724_));
 sky130_fd_sc_hd__xnor2_2 _25381_ (.A(_04723_),
    .B(_04724_),
    .Y(_04725_));
 sky130_fd_sc_hd__xnor2_4 _25382_ (.A(_04722_),
    .B(_04725_),
    .Y(_04726_));
 sky130_fd_sc_hd__a21bo_1 _25383_ (.A1(_04670_),
    .A2(_04671_),
    .B1_N(_04669_),
    .X(_04727_));
 sky130_fd_sc_hd__o21a_1 _25384_ (.A1(_04670_),
    .A2(_04671_),
    .B1(_04727_),
    .X(_04728_));
 sky130_fd_sc_hd__xnor2_1 _25385_ (.A(_03889_),
    .B(_04677_),
    .Y(_04729_));
 sky130_fd_sc_hd__nor2_1 _25386_ (.A(_04518_),
    .B(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__xnor2_2 _25387_ (.A(_04728_),
    .B(_04730_),
    .Y(_04731_));
 sky130_fd_sc_hd__xnor2_4 _25388_ (.A(_04726_),
    .B(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__o21a_1 _25389_ (.A1(_04673_),
    .A2(_04680_),
    .B1(_04681_),
    .X(_04733_));
 sky130_fd_sc_hd__o21ai_1 _25390_ (.A1(_03123_),
    .A2(_04676_),
    .B1(_03124_),
    .Y(_04734_));
 sky130_fd_sc_hd__nand2_1 _25391_ (.A(_03123_),
    .B(_04676_),
    .Y(_04735_));
 sky130_fd_sc_hd__a21oi_2 _25392_ (.A1(_04734_),
    .A2(_04735_),
    .B1(_04518_),
    .Y(_04736_));
 sky130_fd_sc_hd__xnor2_2 _25393_ (.A(_04633_),
    .B(_04736_),
    .Y(_04737_));
 sky130_fd_sc_hd__xnor2_2 _25394_ (.A(_04733_),
    .B(_04737_),
    .Y(_04738_));
 sky130_fd_sc_hd__xnor2_4 _25395_ (.A(_04732_),
    .B(_04738_),
    .Y(_04739_));
 sky130_fd_sc_hd__and2_1 _25396_ (.A(_04685_),
    .B(_04688_),
    .X(_04740_));
 sky130_fd_sc_hd__or2_1 _25397_ (.A(_04685_),
    .B(_04688_),
    .X(_04741_));
 sky130_fd_sc_hd__o21ai_2 _25398_ (.A1(_04683_),
    .A2(_04740_),
    .B1(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__o21ai_1 _25399_ (.A1(_03326_),
    .A2(_04687_),
    .B1(_04371_),
    .Y(_04743_));
 sky130_fd_sc_hd__nand2_1 _25400_ (.A(_04561_),
    .B(_04687_),
    .Y(_04744_));
 sky130_fd_sc_hd__a21oi_2 _25401_ (.A1(_04743_),
    .A2(_04744_),
    .B1(_04518_),
    .Y(_04745_));
 sky130_fd_sc_hd__xnor2_1 _25402_ (.A(_04572_),
    .B(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__xnor2_1 _25403_ (.A(_04742_),
    .B(_04746_),
    .Y(_04747_));
 sky130_fd_sc_hd__xnor2_2 _25404_ (.A(_04739_),
    .B(_04747_),
    .Y(_04748_));
 sky130_fd_sc_hd__o21a_1 _25405_ (.A1(_04411_),
    .A2(_04694_),
    .B1(_04646_),
    .X(_04749_));
 sky130_fd_sc_hd__xnor2_2 _25406_ (.A(_04382_),
    .B(_04749_),
    .Y(_04750_));
 sky130_fd_sc_hd__xnor2_1 _25407_ (.A(_04712_),
    .B(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__xnor2_1 _25408_ (.A(_04748_),
    .B(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__xnor2_1 _25409_ (.A(_04721_),
    .B(_04752_),
    .Y(_04753_));
 sky130_fd_sc_hd__xnor2_2 _25410_ (.A(_04717_),
    .B(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__nor2_1 _25411_ (.A(_04701_),
    .B(_04707_),
    .Y(_04755_));
 sky130_fd_sc_hd__nand2_1 _25412_ (.A(_04701_),
    .B(_04707_),
    .Y(_04756_));
 sky130_fd_sc_hd__o21ai_1 _25413_ (.A1(_04664_),
    .A2(_04755_),
    .B1(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__nand2_1 _25414_ (.A(_04664_),
    .B(_04755_),
    .Y(_04758_));
 sky130_fd_sc_hd__o211a_1 _25415_ (.A1(_04663_),
    .A2(_04757_),
    .B1(_04758_),
    .C1(_04661_),
    .X(_04759_));
 sky130_fd_sc_hd__a2bb2o_1 _25416_ (.A1_N(_04664_),
    .A2_N(_04756_),
    .B1(_04757_),
    .B2(_04663_),
    .X(_04760_));
 sky130_fd_sc_hd__nor2_1 _25417_ (.A(_04661_),
    .B(_04760_),
    .Y(_04761_));
 sky130_fd_sc_hd__inv_2 _25418_ (.A(_04663_),
    .Y(_04762_));
 sky130_fd_sc_hd__nor2_1 _25419_ (.A(_04762_),
    .B(_04664_),
    .Y(_04763_));
 sky130_fd_sc_hd__inv_2 _25420_ (.A(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__o22a_1 _25421_ (.A1(_04663_),
    .A2(_04758_),
    .B1(_04756_),
    .B2(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__o21ai_1 _25422_ (.A1(_04759_),
    .A2(_04761_),
    .B1(_04765_),
    .Y(_04766_));
 sky130_fd_sc_hd__xnor2_1 _25423_ (.A(_04754_),
    .B(_04766_),
    .Y(_04767_));
 sky130_fd_sc_hd__mux2_1 _25424_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[14] ),
    .A1(_04767_),
    .S(_03146_),
    .X(_04768_));
 sky130_fd_sc_hd__clkbuf_1 _25425_ (.A(_04768_),
    .X(_00615_));
 sky130_fd_sc_hd__nor2_1 _25426_ (.A(_04406_),
    .B(_04745_),
    .Y(_04769_));
 sky130_fd_sc_hd__mux2_1 _25427_ (.A0(_04745_),
    .A1(_04769_),
    .S(_04694_),
    .X(_04770_));
 sky130_fd_sc_hd__a21o_1 _25428_ (.A1(_04743_),
    .A2(_04744_),
    .B1(_04518_),
    .X(_04771_));
 sky130_fd_sc_hd__nand2_1 _25429_ (.A(_04516_),
    .B(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__a22o_1 _25430_ (.A1(_04516_),
    .A2(_04770_),
    .B1(_04772_),
    .B2(_04406_),
    .X(_04773_));
 sky130_fd_sc_hd__nand2_1 _25431_ (.A(_04646_),
    .B(_04773_),
    .Y(_04774_));
 sky130_fd_sc_hd__a21o_1 _25432_ (.A1(_03363_),
    .A2(_04437_),
    .B1(_04736_),
    .X(_04775_));
 sky130_fd_sc_hd__a22o_1 _25433_ (.A1(_04561_),
    .A2(_04736_),
    .B1(_04775_),
    .B2(_04371_),
    .X(_04776_));
 sky130_fd_sc_hd__nand2_1 _25434_ (.A(_04726_),
    .B(_04730_),
    .Y(_04777_));
 sky130_fd_sc_hd__or2_1 _25435_ (.A(_04726_),
    .B(_04730_),
    .X(_04778_));
 sky130_fd_sc_hd__mux2_1 _25436_ (.A0(_04777_),
    .A1(_04778_),
    .S(_04728_),
    .X(_04779_));
 sky130_fd_sc_hd__xor2_1 _25437_ (.A(_04776_),
    .B(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__a21oi_1 _25438_ (.A1(_03123_),
    .A2(_03889_),
    .B1(_03124_),
    .Y(_04781_));
 sky130_fd_sc_hd__a21oi_1 _25439_ (.A1(_04190_),
    .A2(_04097_),
    .B1(_04781_),
    .Y(_04782_));
 sky130_fd_sc_hd__nor2_1 _25440_ (.A(_04562_),
    .B(_04631_),
    .Y(_04783_));
 sky130_fd_sc_hd__xnor2_1 _25441_ (.A(_04782_),
    .B(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__nor2_1 _25442_ (.A(_04518_),
    .B(_04784_),
    .Y(_04785_));
 sky130_fd_sc_hd__xnor2_1 _25443_ (.A(_04406_),
    .B(_04785_),
    .Y(_04786_));
 sky130_fd_sc_hd__a211o_1 _25444_ (.A1(_03720_),
    .A2(_03829_),
    .B1(_04131_),
    .C1(_04182_),
    .X(_04787_));
 sky130_fd_sc_hd__a211o_1 _25445_ (.A1(_03722_),
    .A2(_04174_),
    .B1(_04518_),
    .C1(_04272_),
    .X(_04788_));
 sky130_fd_sc_hd__and4_1 _25446_ (.A(_04288_),
    .B(_03936_),
    .C(_04787_),
    .D(_04788_),
    .X(_04789_));
 sky130_fd_sc_hd__a22o_1 _25447_ (.A1(_04288_),
    .A2(_03936_),
    .B1(_04787_),
    .B2(_04788_),
    .X(_04790_));
 sky130_fd_sc_hd__or2b_1 _25448_ (.A(_04789_),
    .B_N(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__a21bo_1 _25449_ (.A1(_04723_),
    .A2(_04724_),
    .B1_N(_04722_),
    .X(_04792_));
 sky130_fd_sc_hd__o21a_1 _25450_ (.A1(_04723_),
    .A2(_04724_),
    .B1(_04792_),
    .X(_04793_));
 sky130_fd_sc_hd__xnor2_1 _25451_ (.A(_04791_),
    .B(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__xnor2_1 _25452_ (.A(_04786_),
    .B(_04794_),
    .Y(_04795_));
 sky130_fd_sc_hd__xnor2_1 _25453_ (.A(_04780_),
    .B(_04795_),
    .Y(_04796_));
 sky130_fd_sc_hd__inv_2 _25454_ (.A(_04737_),
    .Y(_04797_));
 sky130_fd_sc_hd__o21a_1 _25455_ (.A1(_04733_),
    .A2(_04797_),
    .B1(_04732_),
    .X(_04798_));
 sky130_fd_sc_hd__a21oi_1 _25456_ (.A1(_04733_),
    .A2(_04797_),
    .B1(_04798_),
    .Y(_04799_));
 sky130_fd_sc_hd__xnor2_1 _25457_ (.A(_04796_),
    .B(_04799_),
    .Y(_04800_));
 sky130_fd_sc_hd__xnor2_1 _25458_ (.A(_04774_),
    .B(_04800_),
    .Y(_04801_));
 sky130_fd_sc_hd__and3_1 _25459_ (.A(_04742_),
    .B(_04739_),
    .C(_04771_),
    .X(_04802_));
 sky130_fd_sc_hd__nor3_1 _25460_ (.A(_04742_),
    .B(_04739_),
    .C(_04745_),
    .Y(_04803_));
 sky130_fd_sc_hd__and3b_1 _25461_ (.A_N(_04742_),
    .B(_04739_),
    .C(_04572_),
    .X(_04804_));
 sky130_fd_sc_hd__or3b_1 _25462_ (.A(_04572_),
    .B(_04739_),
    .C_N(_04742_),
    .X(_04805_));
 sky130_fd_sc_hd__or4b_2 _25463_ (.A(_04802_),
    .B(_04803_),
    .C(_04804_),
    .D_N(_04805_),
    .X(_04806_));
 sky130_fd_sc_hd__xnor2_2 _25464_ (.A(_04801_),
    .B(_04806_),
    .Y(_04807_));
 sky130_fd_sc_hd__inv_2 _25465_ (.A(_04748_),
    .Y(_04808_));
 sky130_fd_sc_hd__and2_1 _25466_ (.A(_04808_),
    .B(_04750_),
    .X(_04809_));
 sky130_fd_sc_hd__nand2_1 _25467_ (.A(_04721_),
    .B(_04809_),
    .Y(_04810_));
 sky130_fd_sc_hd__o21a_1 _25468_ (.A1(_04808_),
    .A2(_04750_),
    .B1(_04721_),
    .X(_04811_));
 sky130_fd_sc_hd__nor2_1 _25469_ (.A(_04809_),
    .B(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__o21a_1 _25470_ (.A1(_04717_),
    .A2(_04812_),
    .B1(_04810_),
    .X(_04813_));
 sky130_fd_sc_hd__nor2_1 _25471_ (.A(_04721_),
    .B(_04750_),
    .Y(_04814_));
 sky130_fd_sc_hd__nand2_1 _25472_ (.A(_04721_),
    .B(_04750_),
    .Y(_04815_));
 sky130_fd_sc_hd__a21o_1 _25473_ (.A1(_04717_),
    .A2(_04815_),
    .B1(_04814_),
    .X(_04816_));
 sky130_fd_sc_hd__a22o_1 _25474_ (.A1(_04717_),
    .A2(_04814_),
    .B1(_04816_),
    .B2(_04712_),
    .X(_04817_));
 sky130_fd_sc_hd__nand2_1 _25475_ (.A(_04748_),
    .B(_04817_),
    .Y(_04818_));
 sky130_fd_sc_hd__o221a_1 _25476_ (.A1(_04717_),
    .A2(_04810_),
    .B1(_04813_),
    .B2(_04712_),
    .C1(_04818_),
    .X(_04819_));
 sky130_fd_sc_hd__xnor2_2 _25477_ (.A(_04807_),
    .B(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__inv_2 _25478_ (.A(_04754_),
    .Y(_04821_));
 sky130_fd_sc_hd__a21o_1 _25479_ (.A1(_04762_),
    .A2(_04664_),
    .B1(_04821_),
    .X(_04822_));
 sky130_fd_sc_hd__a32o_1 _25480_ (.A1(_04762_),
    .A2(_04664_),
    .A3(_04821_),
    .B1(_04755_),
    .B2(_04822_),
    .X(_04823_));
 sky130_fd_sc_hd__o21a_1 _25481_ (.A1(_04821_),
    .A2(_04755_),
    .B1(_04764_),
    .X(_04824_));
 sky130_fd_sc_hd__a32o_1 _25482_ (.A1(_04821_),
    .A2(_04756_),
    .A3(_04764_),
    .B1(_04824_),
    .B2(_04661_),
    .X(_04825_));
 sky130_fd_sc_hd__a311o_1 _25483_ (.A1(_04661_),
    .A2(_04756_),
    .A3(_04822_),
    .B1(_04823_),
    .C1(_04825_),
    .X(_04826_));
 sky130_fd_sc_hd__xnor2_1 _25484_ (.A(_04820_),
    .B(_04826_),
    .Y(_04827_));
 sky130_fd_sc_hd__mux2_1 _25485_ (.A0(\top0.matmul0.matmul_stage_inst.mult2[15] ),
    .A1(_04827_),
    .S(_03146_),
    .X(_04828_));
 sky130_fd_sc_hd__clkbuf_1 _25486_ (.A(_04828_),
    .X(_00616_));
 sky130_fd_sc_hd__buf_4 _25487_ (.A(_03148_),
    .X(_04829_));
 sky130_fd_sc_hd__mux2_1 _25488_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[0] ),
    .A1(_03641_),
    .S(_04829_),
    .X(_04830_));
 sky130_fd_sc_hd__clkbuf_1 _25489_ (.A(_04830_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _25490_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[1] ),
    .A1(_03756_),
    .S(_04829_),
    .X(_04831_));
 sky130_fd_sc_hd__clkbuf_1 _25491_ (.A(_04831_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _25492_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[2] ),
    .A1(_03855_),
    .S(_04829_),
    .X(_04832_));
 sky130_fd_sc_hd__clkbuf_1 _25493_ (.A(_04832_),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _25494_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[3] ),
    .A1(_03960_),
    .S(_04829_),
    .X(_04833_));
 sky130_fd_sc_hd__clkbuf_1 _25495_ (.A(_04833_),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _25496_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[4] ),
    .A1(_04062_),
    .S(_04829_),
    .X(_04834_));
 sky130_fd_sc_hd__clkbuf_1 _25497_ (.A(_04834_),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _25498_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[5] ),
    .A1(_04154_),
    .S(_04829_),
    .X(_04835_));
 sky130_fd_sc_hd__clkbuf_1 _25499_ (.A(_04835_),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _25500_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[6] ),
    .A1(_04243_),
    .S(_04829_),
    .X(_04836_));
 sky130_fd_sc_hd__clkbuf_1 _25501_ (.A(_04836_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _25502_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[7] ),
    .A1(_04328_),
    .S(_04829_),
    .X(_04837_));
 sky130_fd_sc_hd__clkbuf_1 _25503_ (.A(_04837_),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _25504_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[8] ),
    .A1(_04401_),
    .S(_04829_),
    .X(_04838_));
 sky130_fd_sc_hd__clkbuf_1 _25505_ (.A(_04838_),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _25506_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[9] ),
    .A1(_04470_),
    .S(_04829_),
    .X(_04839_));
 sky130_fd_sc_hd__clkbuf_1 _25507_ (.A(_04839_),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_1 _25508_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[10] ),
    .A1(_04535_),
    .S(_03148_),
    .X(_04840_));
 sky130_fd_sc_hd__clkbuf_1 _25509_ (.A(_04840_),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _25510_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[11] ),
    .A1(_04604_),
    .S(_03148_),
    .X(_04841_));
 sky130_fd_sc_hd__clkbuf_1 _25511_ (.A(_04841_),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _25512_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[12] ),
    .A1(_04659_),
    .S(_03148_),
    .X(_04842_));
 sky130_fd_sc_hd__clkbuf_1 _25513_ (.A(_04842_),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _25514_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[13] ),
    .A1(_04710_),
    .S(_03148_),
    .X(_04843_));
 sky130_fd_sc_hd__clkbuf_1 _25515_ (.A(_04843_),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _25516_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[14] ),
    .A1(_04767_),
    .S(_03148_),
    .X(_04844_));
 sky130_fd_sc_hd__clkbuf_1 _25517_ (.A(_04844_),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _25518_ (.A0(\top0.matmul0.matmul_stage_inst.mult1[15] ),
    .A1(_04827_),
    .S(_03148_),
    .X(_04845_));
 sky130_fd_sc_hd__clkbuf_1 _25519_ (.A(_04845_),
    .X(_00632_));
 sky130_fd_sc_hd__buf_4 _25520_ (.A(_05456_),
    .X(_04846_));
 sky130_fd_sc_hd__mux2_1 _25521_ (.A0(\top0.matmul0.b[0] ),
    .A1(\top0.matmul0.matmul_stage_inst.f[0] ),
    .S(_04846_),
    .X(_04847_));
 sky130_fd_sc_hd__clkbuf_1 _25522_ (.A(_04847_),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _25523_ (.A0(\top0.matmul0.b[1] ),
    .A1(\top0.matmul0.matmul_stage_inst.f[1] ),
    .S(_04846_),
    .X(_04848_));
 sky130_fd_sc_hd__clkbuf_1 _25524_ (.A(_04848_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _25525_ (.A0(\top0.matmul0.b[2] ),
    .A1(\top0.matmul0.matmul_stage_inst.f[2] ),
    .S(_04846_),
    .X(_04849_));
 sky130_fd_sc_hd__clkbuf_1 _25526_ (.A(_04849_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _25527_ (.A0(\top0.matmul0.b[3] ),
    .A1(\top0.matmul0.matmul_stage_inst.f[3] ),
    .S(_04846_),
    .X(_04850_));
 sky130_fd_sc_hd__clkbuf_1 _25528_ (.A(_04850_),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _25529_ (.A0(\top0.matmul0.b[4] ),
    .A1(\top0.matmul0.matmul_stage_inst.f[4] ),
    .S(_04846_),
    .X(_04851_));
 sky130_fd_sc_hd__clkbuf_1 _25530_ (.A(_04851_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _25531_ (.A0(\top0.matmul0.b[5] ),
    .A1(\top0.matmul0.matmul_stage_inst.f[5] ),
    .S(_04846_),
    .X(_04852_));
 sky130_fd_sc_hd__clkbuf_1 _25532_ (.A(_04852_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _25533_ (.A0(\top0.matmul0.b[6] ),
    .A1(\top0.matmul0.matmul_stage_inst.f[6] ),
    .S(_04846_),
    .X(_04853_));
 sky130_fd_sc_hd__clkbuf_1 _25534_ (.A(_04853_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _25535_ (.A0(\top0.matmul0.b[7] ),
    .A1(\top0.matmul0.matmul_stage_inst.f[7] ),
    .S(_04846_),
    .X(_04854_));
 sky130_fd_sc_hd__clkbuf_1 _25536_ (.A(_04854_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _25537_ (.A0(\top0.matmul0.b[8] ),
    .A1(\top0.matmul0.matmul_stage_inst.f[8] ),
    .S(_04846_),
    .X(_04855_));
 sky130_fd_sc_hd__clkbuf_1 _25538_ (.A(_04855_),
    .X(_00641_));
 sky130_fd_sc_hd__clkbuf_4 _25539_ (.A(_05456_),
    .X(_04856_));
 sky130_fd_sc_hd__mux2_1 _25540_ (.A0(\top0.matmul0.b[9] ),
    .A1(\top0.matmul0.matmul_stage_inst.f[9] ),
    .S(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__clkbuf_1 _25541_ (.A(_04857_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _25542_ (.A0(net951),
    .A1(\top0.matmul0.matmul_stage_inst.f[10] ),
    .S(_04856_),
    .X(_04858_));
 sky130_fd_sc_hd__clkbuf_1 _25543_ (.A(_04858_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _25544_ (.A0(\top0.matmul0.b[11] ),
    .A1(\top0.matmul0.matmul_stage_inst.f[11] ),
    .S(_04856_),
    .X(_04859_));
 sky130_fd_sc_hd__clkbuf_1 _25545_ (.A(_04859_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _25546_ (.A0(\top0.matmul0.b[12] ),
    .A1(\top0.matmul0.matmul_stage_inst.f[12] ),
    .S(_04856_),
    .X(_04860_));
 sky130_fd_sc_hd__clkbuf_1 _25547_ (.A(_04860_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _25548_ (.A0(\top0.matmul0.b[13] ),
    .A1(\top0.matmul0.matmul_stage_inst.f[13] ),
    .S(_04856_),
    .X(_04861_));
 sky130_fd_sc_hd__clkbuf_1 _25549_ (.A(_04861_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _25550_ (.A0(\top0.matmul0.b[14] ),
    .A1(\top0.matmul0.matmul_stage_inst.f[14] ),
    .S(_04856_),
    .X(_04862_));
 sky130_fd_sc_hd__clkbuf_1 _25551_ (.A(_04862_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _25552_ (.A0(net943),
    .A1(\top0.matmul0.matmul_stage_inst.f[15] ),
    .S(_04856_),
    .X(_04863_));
 sky130_fd_sc_hd__clkbuf_1 _25553_ (.A(_04863_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _25554_ (.A0(\top0.matmul0.a[0] ),
    .A1(\top0.matmul0.matmul_stage_inst.e[0] ),
    .S(_04856_),
    .X(_04864_));
 sky130_fd_sc_hd__clkbuf_1 _25555_ (.A(_04864_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _25556_ (.A0(\top0.matmul0.a[1] ),
    .A1(\top0.matmul0.matmul_stage_inst.e[1] ),
    .S(_04856_),
    .X(_04865_));
 sky130_fd_sc_hd__clkbuf_1 _25557_ (.A(_04865_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _25558_ (.A0(\top0.matmul0.a[2] ),
    .A1(\top0.matmul0.matmul_stage_inst.e[2] ),
    .S(_04856_),
    .X(_04866_));
 sky130_fd_sc_hd__clkbuf_1 _25559_ (.A(_04866_),
    .X(_00651_));
 sky130_fd_sc_hd__clkbuf_4 _25560_ (.A(_05456_),
    .X(_04867_));
 sky130_fd_sc_hd__mux2_1 _25561_ (.A0(net987),
    .A1(\top0.matmul0.matmul_stage_inst.e[3] ),
    .S(_04867_),
    .X(_04868_));
 sky130_fd_sc_hd__clkbuf_1 _25562_ (.A(_04868_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _25563_ (.A0(\top0.matmul0.a[4] ),
    .A1(\top0.matmul0.matmul_stage_inst.e[4] ),
    .S(_04867_),
    .X(_04869_));
 sky130_fd_sc_hd__clkbuf_1 _25564_ (.A(_04869_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _25565_ (.A0(\top0.matmul0.a[5] ),
    .A1(\top0.matmul0.matmul_stage_inst.e[5] ),
    .S(_04867_),
    .X(_04870_));
 sky130_fd_sc_hd__clkbuf_1 _25566_ (.A(_04870_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _25567_ (.A0(\top0.matmul0.a[6] ),
    .A1(\top0.matmul0.matmul_stage_inst.e[6] ),
    .S(_04867_),
    .X(_04871_));
 sky130_fd_sc_hd__clkbuf_1 _25568_ (.A(_04871_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _25569_ (.A0(\top0.matmul0.a[7] ),
    .A1(\top0.matmul0.matmul_stage_inst.e[7] ),
    .S(_04867_),
    .X(_04872_));
 sky130_fd_sc_hd__clkbuf_1 _25570_ (.A(_04872_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _25571_ (.A0(\top0.matmul0.a[8] ),
    .A1(\top0.matmul0.matmul_stage_inst.e[8] ),
    .S(_04867_),
    .X(_04873_));
 sky130_fd_sc_hd__clkbuf_1 _25572_ (.A(_04873_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _25573_ (.A0(\top0.matmul0.a[9] ),
    .A1(\top0.matmul0.matmul_stage_inst.e[9] ),
    .S(_04867_),
    .X(_04874_));
 sky130_fd_sc_hd__clkbuf_1 _25574_ (.A(_04874_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _25575_ (.A0(\top0.matmul0.a[10] ),
    .A1(\top0.matmul0.matmul_stage_inst.e[10] ),
    .S(_04867_),
    .X(_04875_));
 sky130_fd_sc_hd__clkbuf_1 _25576_ (.A(_04875_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _25577_ (.A0(\top0.matmul0.a[11] ),
    .A1(\top0.matmul0.matmul_stage_inst.e[11] ),
    .S(_04867_),
    .X(_04876_));
 sky130_fd_sc_hd__clkbuf_1 _25578_ (.A(_04876_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _25579_ (.A0(\top0.matmul0.a[12] ),
    .A1(\top0.matmul0.matmul_stage_inst.e[12] ),
    .S(_04867_),
    .X(_04877_));
 sky130_fd_sc_hd__clkbuf_1 _25580_ (.A(_04877_),
    .X(_00661_));
 sky130_fd_sc_hd__clkbuf_4 _25581_ (.A(_05456_),
    .X(_04878_));
 sky130_fd_sc_hd__mux2_1 _25582_ (.A0(\top0.matmul0.a[13] ),
    .A1(\top0.matmul0.matmul_stage_inst.e[13] ),
    .S(_04878_),
    .X(_04879_));
 sky130_fd_sc_hd__clkbuf_1 _25583_ (.A(_04879_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _25584_ (.A0(\top0.matmul0.a[14] ),
    .A1(\top0.matmul0.matmul_stage_inst.e[14] ),
    .S(_04878_),
    .X(_04880_));
 sky130_fd_sc_hd__clkbuf_1 _25585_ (.A(_04880_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _25586_ (.A0(\top0.matmul0.a[15] ),
    .A1(\top0.matmul0.matmul_stage_inst.e[15] ),
    .S(_04878_),
    .X(_04881_));
 sky130_fd_sc_hd__clkbuf_1 _25587_ (.A(_04881_),
    .X(_00664_));
 sky130_fd_sc_hd__and2_1 _25588_ (.A(net70),
    .B(\top0.matmul0.cos[0] ),
    .X(_04882_));
 sky130_fd_sc_hd__inv_2 _25589_ (.A(net73),
    .Y(_04883_));
 sky130_fd_sc_hd__buf_2 _25590_ (.A(_04883_),
    .X(_04884_));
 sky130_fd_sc_hd__inv_2 _25591_ (.A(net69),
    .Y(_04885_));
 sky130_fd_sc_hd__buf_2 _25592_ (.A(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__a21o_1 _25593_ (.A1(_04884_),
    .A2(_04886_),
    .B1(_04846_),
    .X(_04887_));
 sky130_fd_sc_hd__o22a_1 _25594_ (.A1(net759),
    .A2(_00000_),
    .B1(_04882_),
    .B2(_04887_),
    .X(_00665_));
 sky130_fd_sc_hd__or3_1 _25595_ (.A(_04886_),
    .B(\top0.matmul0.cos[1] ),
    .C(_04878_),
    .X(_04888_));
 sky130_fd_sc_hd__o21a_1 _25596_ (.A1(net846),
    .A2(_00000_),
    .B1(_04888_),
    .X(_00666_));
 sky130_fd_sc_hd__and2_1 _25597_ (.A(net71),
    .B(\top0.matmul0.cos[2] ),
    .X(_04889_));
 sky130_fd_sc_hd__buf_2 _25598_ (.A(_05456_),
    .X(_04890_));
 sky130_fd_sc_hd__a21o_2 _25599_ (.A1(net73),
    .A2(_04886_),
    .B1(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__o22a_1 _25600_ (.A1(net750),
    .A2(_00000_),
    .B1(_04889_),
    .B2(_04891_),
    .X(_00667_));
 sky130_fd_sc_hd__or3_1 _25601_ (.A(_04886_),
    .B(\top0.matmul0.cos[4] ),
    .C(_04878_),
    .X(_04892_));
 sky130_fd_sc_hd__o21a_1 _25602_ (.A1(net747),
    .A2(_00000_),
    .B1(_04892_),
    .X(_00668_));
 sky130_fd_sc_hd__or3_1 _25603_ (.A(_04886_),
    .B(\top0.matmul0.cos[5] ),
    .C(_04878_),
    .X(_04893_));
 sky130_fd_sc_hd__o21a_1 _25604_ (.A1(net836),
    .A2(_00000_),
    .B1(_04893_),
    .X(_00669_));
 sky130_fd_sc_hd__and2_1 _25605_ (.A(net70),
    .B(\top0.matmul0.cos[6] ),
    .X(_04894_));
 sky130_fd_sc_hd__o22a_1 _25606_ (.A1(net755),
    .A2(_00000_),
    .B1(_04887_),
    .B2(_04894_),
    .X(_00670_));
 sky130_fd_sc_hd__or3_1 _25607_ (.A(_04886_),
    .B(\top0.matmul0.cos[7] ),
    .C(_04878_),
    .X(_04895_));
 sky130_fd_sc_hd__o21a_1 _25608_ (.A1(net725),
    .A2(_00000_),
    .B1(_04895_),
    .X(_00671_));
 sky130_fd_sc_hd__clkbuf_4 _25609_ (.A(_05457_),
    .X(_04896_));
 sky130_fd_sc_hd__and2_1 _25610_ (.A(net70),
    .B(\top0.matmul0.cos[8] ),
    .X(_04897_));
 sky130_fd_sc_hd__o22a_1 _25611_ (.A1(net739),
    .A2(_04896_),
    .B1(_04891_),
    .B2(_04897_),
    .X(_00672_));
 sky130_fd_sc_hd__and2_1 _25612_ (.A(net70),
    .B(\top0.matmul0.cos[9] ),
    .X(_04898_));
 sky130_fd_sc_hd__o22a_1 _25613_ (.A1(net850),
    .A2(_04896_),
    .B1(_04891_),
    .B2(_04898_),
    .X(_00673_));
 sky130_fd_sc_hd__and2_1 _25614_ (.A(net71),
    .B(\top0.matmul0.cos[10] ),
    .X(_04899_));
 sky130_fd_sc_hd__o22a_1 _25615_ (.A1(net753),
    .A2(_04896_),
    .B1(_04887_),
    .B2(_04899_),
    .X(_00674_));
 sky130_fd_sc_hd__and2_1 _25616_ (.A(net70),
    .B(\top0.matmul0.cos[11] ),
    .X(_04900_));
 sky130_fd_sc_hd__o22a_1 _25617_ (.A1(net752),
    .A2(_04896_),
    .B1(_04891_),
    .B2(_04900_),
    .X(_00675_));
 sky130_fd_sc_hd__and2_1 _25618_ (.A(net70),
    .B(\top0.matmul0.cos[12] ),
    .X(_04901_));
 sky130_fd_sc_hd__o22a_1 _25619_ (.A1(net746),
    .A2(_04896_),
    .B1(_04891_),
    .B2(_04901_),
    .X(_00676_));
 sky130_fd_sc_hd__and2_1 _25620_ (.A(\top0.matmul0.op[1] ),
    .B(\top0.matmul0.cos[13] ),
    .X(_04902_));
 sky130_fd_sc_hd__o22a_1 _25621_ (.A1(net742),
    .A2(_04896_),
    .B1(_04887_),
    .B2(_04902_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _25622_ (.A0(\top0.matmul0.matmul_stage_inst.a[14] ),
    .A1(_04902_),
    .S(_05458_),
    .X(_04903_));
 sky130_fd_sc_hd__clkbuf_1 _25623_ (.A(_04903_),
    .X(_00678_));
 sky130_fd_sc_hd__clkbuf_4 _25624_ (.A(_04890_),
    .X(_04904_));
 sky130_fd_sc_hd__nor2_1 _25625_ (.A(\top0.matmul0.sin[1] ),
    .B(\top0.matmul0.sin[0] ),
    .Y(_04905_));
 sky130_fd_sc_hd__and3_1 _25626_ (.A(_04884_),
    .B(\top0.matmul0.sin[1] ),
    .C(\top0.matmul0.sin[0] ),
    .X(_04906_));
 sky130_fd_sc_hd__o21ai_1 _25627_ (.A1(_04905_),
    .A2(_04906_),
    .B1(net69),
    .Y(_04907_));
 sky130_fd_sc_hd__nand2_1 _25628_ (.A(net69),
    .B(\top0.matmul0.sin[1] ),
    .Y(_04908_));
 sky130_fd_sc_hd__a21oi_1 _25629_ (.A1(net72),
    .A2(_04908_),
    .B1(_04890_),
    .Y(_04909_));
 sky130_fd_sc_hd__a22o_1 _25630_ (.A1(net870),
    .A2(_04904_),
    .B1(_04907_),
    .B2(_04909_),
    .X(_00679_));
 sky130_fd_sc_hd__or2_1 _25631_ (.A(net72),
    .B(_04905_),
    .X(_04910_));
 sky130_fd_sc_hd__xnor2_1 _25632_ (.A(\top0.matmul0.sin[2] ),
    .B(_04910_),
    .Y(_04911_));
 sky130_fd_sc_hd__nor2_1 _25633_ (.A(_04886_),
    .B(_05456_),
    .Y(_04912_));
 sky130_fd_sc_hd__clkbuf_4 _25634_ (.A(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__a22o_1 _25635_ (.A1(net859),
    .A2(_04904_),
    .B1(_04911_),
    .B2(_04913_),
    .X(_00680_));
 sky130_fd_sc_hd__or4_4 _25636_ (.A(\top0.matmul0.sin[1] ),
    .B(\top0.matmul0.sin[0] ),
    .C(\top0.matmul0.sin[2] ),
    .D(\top0.matmul0.sin[3] ),
    .X(_04914_));
 sky130_fd_sc_hd__inv_2 _25637_ (.A(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__o311a_1 _25638_ (.A1(\top0.matmul0.sin[1] ),
    .A2(\top0.matmul0.sin[0] ),
    .A3(\top0.matmul0.sin[2] ),
    .B1(\top0.matmul0.sin[3] ),
    .C1(_04884_),
    .X(_04916_));
 sky130_fd_sc_hd__o21ai_1 _25639_ (.A1(_04915_),
    .A2(_04916_),
    .B1(net69),
    .Y(_04917_));
 sky130_fd_sc_hd__nand2_1 _25640_ (.A(net69),
    .B(\top0.matmul0.sin[3] ),
    .Y(_04918_));
 sky130_fd_sc_hd__a21oi_1 _25641_ (.A1(net72),
    .A2(_04918_),
    .B1(_04890_),
    .Y(_04919_));
 sky130_fd_sc_hd__a22o_1 _25642_ (.A1(net847),
    .A2(_04904_),
    .B1(_04917_),
    .B2(_04919_),
    .X(_00681_));
 sky130_fd_sc_hd__nor2_1 _25643_ (.A(\top0.matmul0.sin[4] ),
    .B(_04914_),
    .Y(_04920_));
 sky130_fd_sc_hd__and3_1 _25644_ (.A(_04884_),
    .B(\top0.matmul0.sin[4] ),
    .C(_04914_),
    .X(_04921_));
 sky130_fd_sc_hd__o21ai_1 _25645_ (.A1(_04920_),
    .A2(_04921_),
    .B1(net69),
    .Y(_04922_));
 sky130_fd_sc_hd__nand2_1 _25646_ (.A(net69),
    .B(\top0.matmul0.sin[4] ),
    .Y(_04923_));
 sky130_fd_sc_hd__a21oi_1 _25647_ (.A1(net72),
    .A2(_04923_),
    .B1(_04890_),
    .Y(_04924_));
 sky130_fd_sc_hd__a22o_1 _25648_ (.A1(net822),
    .A2(_04904_),
    .B1(_04922_),
    .B2(_04924_),
    .X(_00682_));
 sky130_fd_sc_hd__clkbuf_4 _25649_ (.A(_04890_),
    .X(_04925_));
 sky130_fd_sc_hd__or3_2 _25650_ (.A(\top0.matmul0.sin[4] ),
    .B(\top0.matmul0.sin[5] ),
    .C(_04914_),
    .X(_04926_));
 sky130_fd_sc_hd__or3b_1 _25651_ (.A(net73),
    .B(_04920_),
    .C_N(\top0.matmul0.sin[5] ),
    .X(_04927_));
 sky130_fd_sc_hd__nand2_1 _25652_ (.A(_04926_),
    .B(_04927_),
    .Y(_04928_));
 sky130_fd_sc_hd__nand2_1 _25653_ (.A(net71),
    .B(\top0.matmul0.sin[5] ),
    .Y(_04929_));
 sky130_fd_sc_hd__a221o_1 _25654_ (.A1(net71),
    .A2(_04928_),
    .B1(_04929_),
    .B2(net73),
    .C1(_04878_),
    .X(_04930_));
 sky130_fd_sc_hd__a21bo_1 _25655_ (.A1(net799),
    .A2(_04925_),
    .B1_N(_04930_),
    .X(_00683_));
 sky130_fd_sc_hd__or2_2 _25656_ (.A(\top0.matmul0.sin[6] ),
    .B(_04926_),
    .X(_04931_));
 sky130_fd_sc_hd__nand3_1 _25657_ (.A(_04883_),
    .B(\top0.matmul0.sin[6] ),
    .C(_04926_),
    .Y(_04932_));
 sky130_fd_sc_hd__nand2_1 _25658_ (.A(_04931_),
    .B(_04932_),
    .Y(_04933_));
 sky130_fd_sc_hd__nand2_1 _25659_ (.A(net71),
    .B(\top0.matmul0.sin[6] ),
    .Y(_04934_));
 sky130_fd_sc_hd__a221o_1 _25660_ (.A1(net71),
    .A2(_04933_),
    .B1(_04934_),
    .B2(net74),
    .C1(_04878_),
    .X(_04935_));
 sky130_fd_sc_hd__a21bo_1 _25661_ (.A1(net735),
    .A2(_04904_),
    .B1_N(_04935_),
    .X(_00684_));
 sky130_fd_sc_hd__clkbuf_4 _25662_ (.A(_04913_),
    .X(_04936_));
 sky130_fd_sc_hd__and2_1 _25663_ (.A(_04884_),
    .B(_04931_),
    .X(_04937_));
 sky130_fd_sc_hd__xor2_1 _25664_ (.A(\top0.matmul0.sin[7] ),
    .B(_04937_),
    .X(_04938_));
 sky130_fd_sc_hd__a22o_1 _25665_ (.A1(net779),
    .A2(_04904_),
    .B1(_04936_),
    .B2(_04938_),
    .X(_00685_));
 sky130_fd_sc_hd__o21a_1 _25666_ (.A1(\top0.matmul0.sin[7] ),
    .A2(_04931_),
    .B1(_04884_),
    .X(_04939_));
 sky130_fd_sc_hd__xor2_1 _25667_ (.A(\top0.matmul0.sin[8] ),
    .B(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__a22o_1 _25668_ (.A1(net791),
    .A2(_04904_),
    .B1(_04936_),
    .B2(_04940_),
    .X(_00686_));
 sky130_fd_sc_hd__or3_1 _25669_ (.A(\top0.matmul0.sin[7] ),
    .B(\top0.matmul0.sin[8] ),
    .C(_04931_),
    .X(_04941_));
 sky130_fd_sc_hd__or2_2 _25670_ (.A(\top0.matmul0.sin[9] ),
    .B(_04941_),
    .X(_04942_));
 sky130_fd_sc_hd__nand3_1 _25671_ (.A(_04883_),
    .B(\top0.matmul0.sin[9] ),
    .C(_04941_),
    .Y(_04943_));
 sky130_fd_sc_hd__nand2_1 _25672_ (.A(_04942_),
    .B(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__nand2_1 _25673_ (.A(net71),
    .B(\top0.matmul0.sin[9] ),
    .Y(_04945_));
 sky130_fd_sc_hd__a221o_1 _25674_ (.A1(net71),
    .A2(_04944_),
    .B1(_04945_),
    .B2(net74),
    .C1(_05456_),
    .X(_04946_));
 sky130_fd_sc_hd__a21bo_1 _25675_ (.A1(net805),
    .A2(_04904_),
    .B1_N(_04946_),
    .X(_00687_));
 sky130_fd_sc_hd__and2_1 _25676_ (.A(_04884_),
    .B(_04942_),
    .X(_04947_));
 sky130_fd_sc_hd__xor2_1 _25677_ (.A(\top0.matmul0.sin[10] ),
    .B(_04947_),
    .X(_04948_));
 sky130_fd_sc_hd__a22o_1 _25678_ (.A1(net854),
    .A2(_04904_),
    .B1(_04936_),
    .B2(_04948_),
    .X(_00688_));
 sky130_fd_sc_hd__o21a_1 _25679_ (.A1(\top0.matmul0.sin[10] ),
    .A2(_04942_),
    .B1(_04884_),
    .X(_04949_));
 sky130_fd_sc_hd__xor2_1 _25680_ (.A(\top0.matmul0.sin[11] ),
    .B(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__a22o_1 _25681_ (.A1(net825),
    .A2(_04904_),
    .B1(_04936_),
    .B2(_04950_),
    .X(_00689_));
 sky130_fd_sc_hd__or3_1 _25682_ (.A(\top0.matmul0.sin[10] ),
    .B(\top0.matmul0.sin[11] ),
    .C(_04942_),
    .X(_04951_));
 sky130_fd_sc_hd__and2_1 _25683_ (.A(_04884_),
    .B(_04951_),
    .X(_04952_));
 sky130_fd_sc_hd__xnor2_1 _25684_ (.A(\top0.matmul0.sin[12] ),
    .B(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__o2bb2a_1 _25685_ (.A1_N(_04913_),
    .A2_N(_04953_),
    .B1(net841),
    .B2(_00000_),
    .X(_00690_));
 sky130_fd_sc_hd__or2_1 _25686_ (.A(\top0.matmul0.sin[12] ),
    .B(_04951_),
    .X(_04954_));
 sky130_fd_sc_hd__mux2_1 _25687_ (.A0(_04885_),
    .A1(_04954_),
    .S(_04883_),
    .X(_04955_));
 sky130_fd_sc_hd__a21oi_1 _25688_ (.A1(\top0.matmul0.sin[13] ),
    .A2(_04954_),
    .B1(_04886_),
    .Y(_04956_));
 sky130_fd_sc_hd__o221a_1 _25689_ (.A1(\top0.matmul0.sin[13] ),
    .A2(_04955_),
    .B1(_04956_),
    .B2(net72),
    .C1(_04896_),
    .X(_04957_));
 sky130_fd_sc_hd__a21o_1 _25690_ (.A1(net714),
    .A2(_04925_),
    .B1(_04957_),
    .X(_00691_));
 sky130_fd_sc_hd__or4b_1 _25691_ (.A(net72),
    .B(_04885_),
    .C(\top0.matmul0.sin[13] ),
    .D_N(_04954_),
    .X(_04958_));
 sky130_fd_sc_hd__o21ai_1 _25692_ (.A1(_04886_),
    .A2(\top0.matmul0.sin[13] ),
    .B1(net73),
    .Y(_04959_));
 sky130_fd_sc_hd__and3_1 _25693_ (.A(_05457_),
    .B(_04958_),
    .C(_04959_),
    .X(_04960_));
 sky130_fd_sc_hd__o21ba_1 _25694_ (.A1(\top0.matmul0.matmul_stage_inst.c[14] ),
    .A2(_04896_),
    .B1_N(_04960_),
    .X(_04961_));
 sky130_fd_sc_hd__clkbuf_1 _25695_ (.A(_04961_),
    .X(_00692_));
 sky130_fd_sc_hd__o21ba_1 _25696_ (.A1(\top0.matmul0.matmul_stage_inst.c[15] ),
    .A2(_04896_),
    .B1_N(_04960_),
    .X(_04962_));
 sky130_fd_sc_hd__clkbuf_1 _25697_ (.A(_04962_),
    .X(_00693_));
 sky130_fd_sc_hd__and3_1 _25698_ (.A(net69),
    .B(\top0.matmul0.sin[0] ),
    .C(_04896_),
    .X(_04963_));
 sky130_fd_sc_hd__a21o_1 _25699_ (.A1(net862),
    .A2(_04925_),
    .B1(_04963_),
    .X(_00694_));
 sky130_fd_sc_hd__clkbuf_4 _25700_ (.A(_04890_),
    .X(_04964_));
 sky130_fd_sc_hd__nand2_1 _25701_ (.A(net72),
    .B(\top0.matmul0.sin[0] ),
    .Y(_04965_));
 sky130_fd_sc_hd__xnor2_1 _25702_ (.A(\top0.matmul0.sin[1] ),
    .B(_04965_),
    .Y(_04966_));
 sky130_fd_sc_hd__a22o_1 _25703_ (.A1(net887),
    .A2(_04964_),
    .B1(_04936_),
    .B2(_04966_),
    .X(_00695_));
 sky130_fd_sc_hd__or2_1 _25704_ (.A(_04884_),
    .B(_04905_),
    .X(_04967_));
 sky130_fd_sc_hd__xnor2_1 _25705_ (.A(\top0.matmul0.sin[2] ),
    .B(_04967_),
    .Y(_04968_));
 sky130_fd_sc_hd__a22o_1 _25706_ (.A1(net871),
    .A2(_04964_),
    .B1(_04936_),
    .B2(_04968_),
    .X(_00696_));
 sky130_fd_sc_hd__o31a_1 _25707_ (.A1(\top0.matmul0.sin[1] ),
    .A2(\top0.matmul0.sin[0] ),
    .A3(\top0.matmul0.sin[2] ),
    .B1(net72),
    .X(_04969_));
 sky130_fd_sc_hd__xor2_1 _25708_ (.A(\top0.matmul0.sin[3] ),
    .B(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__a22o_1 _25709_ (.A1(net819),
    .A2(_04964_),
    .B1(_04936_),
    .B2(_04970_),
    .X(_00697_));
 sky130_fd_sc_hd__nand2_1 _25710_ (.A(net72),
    .B(_04914_),
    .Y(_04971_));
 sky130_fd_sc_hd__xnor2_1 _25711_ (.A(\top0.matmul0.sin[4] ),
    .B(_04971_),
    .Y(_04972_));
 sky130_fd_sc_hd__a22o_1 _25712_ (.A1(net784),
    .A2(_04964_),
    .B1(_04936_),
    .B2(_04972_),
    .X(_00698_));
 sky130_fd_sc_hd__or2_1 _25713_ (.A(_04883_),
    .B(_04920_),
    .X(_04973_));
 sky130_fd_sc_hd__xnor2_1 _25714_ (.A(\top0.matmul0.sin[5] ),
    .B(_04973_),
    .Y(_04974_));
 sky130_fd_sc_hd__a22o_1 _25715_ (.A1(net866),
    .A2(_04964_),
    .B1(_04936_),
    .B2(_04974_),
    .X(_00699_));
 sky130_fd_sc_hd__nand2_1 _25716_ (.A(net73),
    .B(_04926_),
    .Y(_04975_));
 sky130_fd_sc_hd__xnor2_1 _25717_ (.A(\top0.matmul0.sin[6] ),
    .B(_04975_),
    .Y(_04976_));
 sky130_fd_sc_hd__a22o_1 _25718_ (.A1(net764),
    .A2(_04964_),
    .B1(_04936_),
    .B2(_04976_),
    .X(_00700_));
 sky130_fd_sc_hd__nand2_1 _25719_ (.A(net74),
    .B(_04931_),
    .Y(_04977_));
 sky130_fd_sc_hd__xnor2_1 _25720_ (.A(\top0.matmul0.sin[7] ),
    .B(_04977_),
    .Y(_04978_));
 sky130_fd_sc_hd__a22o_1 _25721_ (.A1(net792),
    .A2(_04964_),
    .B1(_04913_),
    .B2(_04978_),
    .X(_00701_));
 sky130_fd_sc_hd__o21ai_1 _25722_ (.A1(\top0.matmul0.sin[7] ),
    .A2(_04931_),
    .B1(net74),
    .Y(_04979_));
 sky130_fd_sc_hd__xnor2_1 _25723_ (.A(\top0.matmul0.sin[8] ),
    .B(_04979_),
    .Y(_04980_));
 sky130_fd_sc_hd__a22o_1 _25724_ (.A1(net856),
    .A2(_04964_),
    .B1(_04913_),
    .B2(_04980_),
    .X(_00702_));
 sky130_fd_sc_hd__nand2_1 _25725_ (.A(net74),
    .B(_04941_),
    .Y(_04981_));
 sky130_fd_sc_hd__xnor2_1 _25726_ (.A(\top0.matmul0.sin[9] ),
    .B(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__a22o_1 _25727_ (.A1(net906),
    .A2(_04964_),
    .B1(_04913_),
    .B2(_04982_),
    .X(_00703_));
 sky130_fd_sc_hd__nand2_1 _25728_ (.A(net74),
    .B(_04942_),
    .Y(_04983_));
 sky130_fd_sc_hd__xnor2_1 _25729_ (.A(\top0.matmul0.sin[10] ),
    .B(_04983_),
    .Y(_04984_));
 sky130_fd_sc_hd__a22o_1 _25730_ (.A1(net808),
    .A2(_04964_),
    .B1(_04913_),
    .B2(_04984_),
    .X(_00704_));
 sky130_fd_sc_hd__o21ai_1 _25731_ (.A1(\top0.matmul0.sin[10] ),
    .A2(_04942_),
    .B1(net73),
    .Y(_04985_));
 sky130_fd_sc_hd__xnor2_1 _25732_ (.A(\top0.matmul0.sin[11] ),
    .B(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__a22o_1 _25733_ (.A1(net891),
    .A2(_04890_),
    .B1(_04913_),
    .B2(_04986_),
    .X(_00705_));
 sky130_fd_sc_hd__nand2_1 _25734_ (.A(net72),
    .B(_04951_),
    .Y(_04987_));
 sky130_fd_sc_hd__xnor2_1 _25735_ (.A(\top0.matmul0.sin[12] ),
    .B(_04987_),
    .Y(_04988_));
 sky130_fd_sc_hd__a22o_1 _25736_ (.A1(net813),
    .A2(_04890_),
    .B1(_04913_),
    .B2(_04988_),
    .X(_00706_));
 sky130_fd_sc_hd__nand2_1 _25737_ (.A(net73),
    .B(_04954_),
    .Y(_04989_));
 sky130_fd_sc_hd__xnor2_1 _25738_ (.A(\top0.matmul0.sin[13] ),
    .B(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__a22o_1 _25739_ (.A1(net786),
    .A2(_04890_),
    .B1(_04913_),
    .B2(_04990_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _25740_ (.A0(_04989_),
    .A1(net73),
    .S(\top0.matmul0.sin[13] ),
    .X(_04991_));
 sky130_fd_sc_hd__and2b_1 _25741_ (.A_N(_04991_),
    .B(_04912_),
    .X(_04992_));
 sky130_fd_sc_hd__a21o_1 _25742_ (.A1(net778),
    .A2(_04925_),
    .B1(_04992_),
    .X(_00708_));
 sky130_fd_sc_hd__a21o_1 _25743_ (.A1(net711),
    .A2(_04925_),
    .B1(_04992_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _25744_ (.A0(net993),
    .A1(_04882_),
    .S(_05458_),
    .X(_04993_));
 sky130_fd_sc_hd__clkbuf_1 _25745_ (.A(_04993_),
    .X(_00710_));
 sky130_fd_sc_hd__and3_1 _25746_ (.A(net69),
    .B(\top0.matmul0.cos[1] ),
    .C(_05458_),
    .X(_04994_));
 sky130_fd_sc_hd__a21o_1 _25747_ (.A1(net768),
    .A2(_04925_),
    .B1(_04994_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _25748_ (.A0(\top0.matmul0.matmul_stage_inst.a[2] ),
    .A1(_04889_),
    .S(_05458_),
    .X(_04995_));
 sky130_fd_sc_hd__clkbuf_1 _25749_ (.A(_04995_),
    .X(_00712_));
 sky130_fd_sc_hd__and3_1 _25750_ (.A(net70),
    .B(\top0.matmul0.cos[3] ),
    .C(_05458_),
    .X(_04996_));
 sky130_fd_sc_hd__a21o_1 _25751_ (.A1(net770),
    .A2(_04925_),
    .B1(_04996_),
    .X(_00713_));
 sky130_fd_sc_hd__and3_1 _25752_ (.A(net69),
    .B(\top0.matmul0.cos[4] ),
    .C(_05458_),
    .X(_04997_));
 sky130_fd_sc_hd__a21o_1 _25753_ (.A1(net717),
    .A2(_04925_),
    .B1(_04997_),
    .X(_00714_));
 sky130_fd_sc_hd__and3_1 _25754_ (.A(net70),
    .B(\top0.matmul0.cos[5] ),
    .C(_05458_),
    .X(_04998_));
 sky130_fd_sc_hd__a21o_1 _25755_ (.A1(net767),
    .A2(_04925_),
    .B1(_04998_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _25756_ (.A0(\top0.matmul0.matmul_stage_inst.a[6] ),
    .A1(_04894_),
    .S(_05458_),
    .X(_04999_));
 sky130_fd_sc_hd__clkbuf_1 _25757_ (.A(_04999_),
    .X(_00716_));
 sky130_fd_sc_hd__and3_1 _25758_ (.A(net70),
    .B(\top0.matmul0.cos[7] ),
    .C(_05458_),
    .X(_05000_));
 sky130_fd_sc_hd__a21o_1 _25759_ (.A1(net716),
    .A2(_04925_),
    .B1(_05000_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _25760_ (.A0(\top0.matmul0.matmul_stage_inst.a[8] ),
    .A1(_04897_),
    .S(_05457_),
    .X(_05001_));
 sky130_fd_sc_hd__clkbuf_1 _25761_ (.A(_05001_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _25762_ (.A0(\top0.matmul0.matmul_stage_inst.a[9] ),
    .A1(_04898_),
    .S(_05457_),
    .X(_05002_));
 sky130_fd_sc_hd__clkbuf_1 _25763_ (.A(_05002_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _25764_ (.A0(\top0.matmul0.matmul_stage_inst.a[10] ),
    .A1(_04899_),
    .S(_05457_),
    .X(_05003_));
 sky130_fd_sc_hd__clkbuf_1 _25765_ (.A(_05003_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _25766_ (.A0(\top0.matmul0.matmul_stage_inst.a[11] ),
    .A1(_04900_),
    .S(_05457_),
    .X(_05004_));
 sky130_fd_sc_hd__clkbuf_1 _25767_ (.A(_05004_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _25768_ (.A0(\top0.matmul0.matmul_stage_inst.a[12] ),
    .A1(_04901_),
    .S(_05457_),
    .X(_05005_));
 sky130_fd_sc_hd__clkbuf_1 _25769_ (.A(_05005_),
    .X(_00722_));
 sky130_fd_sc_hd__or3_1 _25770_ (.A(_04886_),
    .B(\top0.matmul0.cos[13] ),
    .C(_04878_),
    .X(_05006_));
 sky130_fd_sc_hd__o21a_1 _25771_ (.A1(net730),
    .A2(_00000_),
    .B1(_05006_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _25772_ (.A0(\top0.matmul0.op_in[0] ),
    .A1(net74),
    .S(_05460_),
    .X(_05007_));
 sky130_fd_sc_hd__clkbuf_1 _25773_ (.A(_05007_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _25774_ (.A0(\top0.matmul0.op_in[1] ),
    .A1(net70),
    .S(_05460_),
    .X(_05008_));
 sky130_fd_sc_hd__clkbuf_1 _25775_ (.A(_05008_),
    .X(_00725_));
 sky130_fd_sc_hd__or2_1 _25776_ (.A(_12009_),
    .B(net205),
    .X(_05009_));
 sky130_fd_sc_hd__o21a_1 _25777_ (.A1(_02282_),
    .A2(_05009_),
    .B1(_05427_),
    .X(_05010_));
 sky130_fd_sc_hd__a21oi_1 _25778_ (.A1(net207),
    .A2(net209),
    .B1(_05010_),
    .Y(_00726_));
 sky130_fd_sc_hd__a21o_1 _25779_ (.A1(net205),
    .A2(_02282_),
    .B1(_12019_),
    .X(_05011_));
 sky130_fd_sc_hd__o21ai_1 _25780_ (.A1(_12030_),
    .A2(_12023_),
    .B1(_05011_),
    .Y(_05012_));
 sky130_fd_sc_hd__nor2_2 _25781_ (.A(net205),
    .B(_12019_),
    .Y(_05013_));
 sky130_fd_sc_hd__clkbuf_4 _25782_ (.A(_05013_),
    .X(_05014_));
 sky130_fd_sc_hd__or2b_2 _25783_ (.A(net208),
    .B_N(net205),
    .X(_05015_));
 sky130_fd_sc_hd__o21ai_1 _25784_ (.A1(\top0.pid_d.out_valid ),
    .A2(_12030_),
    .B1(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__a22o_1 _25785_ (.A1(_05425_),
    .A2(_05014_),
    .B1(_05016_),
    .B2(net207),
    .X(_05017_));
 sky130_fd_sc_hd__mux2_1 _25786_ (.A0(_05012_),
    .A1(\top0.matmul0.start ),
    .S(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__clkbuf_1 _25787_ (.A(_05018_),
    .X(_00727_));
 sky130_fd_sc_hd__a2bb2o_1 _25788_ (.A1_N(net208),
    .A2_N(_12017_),
    .B1(\top0.cordic0.in_valid ),
    .B2(net205),
    .X(_05019_));
 sky130_fd_sc_hd__nand2_1 _25789_ (.A(net208),
    .B(_05009_),
    .Y(_05020_));
 sky130_fd_sc_hd__a22o_1 _25790_ (.A1(_12009_),
    .A2(_05019_),
    .B1(_05020_),
    .B2(\top0.cordic0.in_valid ),
    .X(_00728_));
 sky130_fd_sc_hd__nand2_1 _25791_ (.A(_12009_),
    .B(net205),
    .Y(_05021_));
 sky130_fd_sc_hd__and3_1 _25792_ (.A(net208),
    .B(_05009_),
    .C(_05021_),
    .X(_05022_));
 sky130_fd_sc_hd__a21o_1 _25793_ (.A1(_05439_),
    .A2(_05022_),
    .B1(\top0.clarke_done ),
    .X(_05023_));
 sky130_fd_sc_hd__nand2_1 _25794_ (.A(_12024_),
    .B(_05022_),
    .Y(_05024_));
 sky130_fd_sc_hd__and2_1 _25795_ (.A(_05023_),
    .B(_05024_),
    .X(_05025_));
 sky130_fd_sc_hd__clkbuf_1 _25796_ (.A(_05025_),
    .X(_00729_));
 sky130_fd_sc_hd__a21o_1 _25797_ (.A1(\top0.cordic0.out_valid ),
    .A2(_05022_),
    .B1(\top0.cordic_done ),
    .X(_05026_));
 sky130_fd_sc_hd__and2_1 _25798_ (.A(_05024_),
    .B(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__clkbuf_1 _25799_ (.A(_05027_),
    .X(_00730_));
 sky130_fd_sc_hd__a21o_2 _25800_ (.A1(_12009_),
    .A2(_02282_),
    .B1(_12012_),
    .X(_05028_));
 sky130_fd_sc_hd__buf_2 _25801_ (.A(_05028_),
    .X(_05029_));
 sky130_fd_sc_hd__nor2_1 _25802_ (.A(_02282_),
    .B(_12014_),
    .Y(_05030_));
 sky130_fd_sc_hd__clkbuf_4 _25803_ (.A(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__xor2_1 _25804_ (.A(\top0.matmul0.alpha_pass[0] ),
    .B(\top0.matmul0.beta_pass[0] ),
    .X(_05032_));
 sky130_fd_sc_hd__a22o_1 _25805_ (.A1(net833),
    .A2(_05029_),
    .B1(_05031_),
    .B2(_05032_),
    .X(_00731_));
 sky130_fd_sc_hd__or2_1 _25806_ (.A(\top0.matmul0.alpha_pass[1] ),
    .B(\top0.matmul0.beta_pass[1] ),
    .X(_05033_));
 sky130_fd_sc_hd__nand2_1 _25807_ (.A(\top0.matmul0.alpha_pass[1] ),
    .B(\top0.matmul0.beta_pass[1] ),
    .Y(_05034_));
 sky130_fd_sc_hd__nor2_1 _25808_ (.A(\top0.matmul0.alpha_pass[0] ),
    .B(\top0.matmul0.beta_pass[0] ),
    .Y(_05035_));
 sky130_fd_sc_hd__a21oi_1 _25809_ (.A1(_05033_),
    .A2(_05034_),
    .B1(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__and3_1 _25810_ (.A(_05035_),
    .B(_05033_),
    .C(_05034_),
    .X(_05037_));
 sky130_fd_sc_hd__or2_1 _25811_ (.A(_05036_),
    .B(_05037_),
    .X(_05038_));
 sky130_fd_sc_hd__a22o_1 _25812_ (.A1(\top0.c_out_calc[1] ),
    .A2(_05029_),
    .B1(_05031_),
    .B2(_05038_),
    .X(_00732_));
 sky130_fd_sc_hd__xnor2_2 _25813_ (.A(\top0.matmul0.alpha_pass[2] ),
    .B(\top0.matmul0.beta_pass[2] ),
    .Y(_05039_));
 sky130_fd_sc_hd__mux2_1 _25814_ (.A0(_05034_),
    .A1(_05033_),
    .S(_05035_),
    .X(_05040_));
 sky130_fd_sc_hd__xnor2_1 _25815_ (.A(_05039_),
    .B(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__a22o_1 _25816_ (.A1(net798),
    .A2(_05029_),
    .B1(_05031_),
    .B2(_05041_),
    .X(_00733_));
 sky130_fd_sc_hd__and2_1 _25817_ (.A(\top0.matmul0.alpha_pass[1] ),
    .B(\top0.matmul0.beta_pass[1] ),
    .X(_05042_));
 sky130_fd_sc_hd__o21bai_2 _25818_ (.A1(_05042_),
    .A2(_05039_),
    .B1_N(_05035_),
    .Y(_05043_));
 sky130_fd_sc_hd__nand2_1 _25819_ (.A(_05033_),
    .B(_05039_),
    .Y(_05044_));
 sky130_fd_sc_hd__nand2_1 _25820_ (.A(_05043_),
    .B(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__nor2_1 _25821_ (.A(\top0.matmul0.alpha_pass[2] ),
    .B(\top0.matmul0.beta_pass[2] ),
    .Y(_05046_));
 sky130_fd_sc_hd__xor2_2 _25822_ (.A(\top0.matmul0.alpha_pass[3] ),
    .B(\top0.matmul0.beta_pass[3] ),
    .X(_05047_));
 sky130_fd_sc_hd__xor2_1 _25823_ (.A(_05046_),
    .B(_05047_),
    .X(_05048_));
 sky130_fd_sc_hd__xnor2_1 _25824_ (.A(_05045_),
    .B(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__a22o_1 _25825_ (.A1(\top0.c_out_calc[3] ),
    .A2(_05029_),
    .B1(_05031_),
    .B2(_05049_),
    .X(_00734_));
 sky130_fd_sc_hd__a31o_1 _25826_ (.A1(_05043_),
    .A2(_05044_),
    .A3(_05047_),
    .B1(_05046_),
    .X(_05050_));
 sky130_fd_sc_hd__a21o_1 _25827_ (.A1(_05043_),
    .A2(_05044_),
    .B1(_05047_),
    .X(_05051_));
 sky130_fd_sc_hd__and2_1 _25828_ (.A(_05050_),
    .B(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__nor2_1 _25829_ (.A(\top0.matmul0.alpha_pass[3] ),
    .B(\top0.matmul0.beta_pass[3] ),
    .Y(_05053_));
 sky130_fd_sc_hd__xor2_2 _25830_ (.A(\top0.matmul0.alpha_pass[4] ),
    .B(\top0.matmul0.beta_pass[4] ),
    .X(_05054_));
 sky130_fd_sc_hd__xnor2_1 _25831_ (.A(_05053_),
    .B(_05054_),
    .Y(_05055_));
 sky130_fd_sc_hd__xnor2_1 _25832_ (.A(_05052_),
    .B(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__a22o_1 _25833_ (.A1(\top0.c_out_calc[4] ),
    .A2(_05029_),
    .B1(_05031_),
    .B2(_05056_),
    .X(_00735_));
 sky130_fd_sc_hd__a31o_1 _25834_ (.A1(_05050_),
    .A2(_05051_),
    .A3(_05054_),
    .B1(_05053_),
    .X(_05057_));
 sky130_fd_sc_hd__o21ai_2 _25835_ (.A1(_05052_),
    .A2(_05054_),
    .B1(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__or2_2 _25836_ (.A(\top0.matmul0.alpha_pass[4] ),
    .B(\top0.matmul0.beta_pass[4] ),
    .X(_05059_));
 sky130_fd_sc_hd__xor2_1 _25837_ (.A(net76),
    .B(\top0.matmul0.beta_pass[5] ),
    .X(_05060_));
 sky130_fd_sc_hd__xnor2_1 _25838_ (.A(_05059_),
    .B(_05060_),
    .Y(_05061_));
 sky130_fd_sc_hd__xnor2_1 _25839_ (.A(_05058_),
    .B(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__a22o_1 _25840_ (.A1(net743),
    .A2(_05029_),
    .B1(_05031_),
    .B2(_05062_),
    .X(_00736_));
 sky130_fd_sc_hd__or2_1 _25841_ (.A(\top0.matmul0.beta_pass[5] ),
    .B(_05058_),
    .X(_05063_));
 sky130_fd_sc_hd__o211a_1 _25842_ (.A1(net76),
    .A2(_05059_),
    .B1(_05058_),
    .C1(\top0.matmul0.beta_pass[5] ),
    .X(_05064_));
 sky130_fd_sc_hd__a31o_1 _25843_ (.A1(net76),
    .A2(_05059_),
    .A3(_05063_),
    .B1(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__nor4_1 _25844_ (.A(net76),
    .B(\top0.matmul0.beta_pass[5] ),
    .C(_05058_),
    .D(_05059_),
    .Y(_05066_));
 sky130_fd_sc_hd__xnor2_1 _25845_ (.A(\top0.matmul0.alpha_pass[6] ),
    .B(\top0.matmul0.beta_pass[6] ),
    .Y(_05067_));
 sky130_fd_sc_hd__o21ai_1 _25846_ (.A1(_05065_),
    .A2(_05066_),
    .B1(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hd__or3_1 _25847_ (.A(_05067_),
    .B(_05065_),
    .C(net12),
    .X(_05069_));
 sky130_fd_sc_hd__a32o_1 _25848_ (.A1(_05031_),
    .A2(_05068_),
    .A3(_05069_),
    .B1(_05028_),
    .B2(net867),
    .X(_00737_));
 sky130_fd_sc_hd__xnor2_2 _25849_ (.A(\top0.matmul0.alpha_pass[7] ),
    .B(\top0.matmul0.beta_pass[7] ),
    .Y(_05070_));
 sky130_fd_sc_hd__or4_1 _25850_ (.A(\top0.matmul0.alpha_pass[4] ),
    .B(\top0.matmul0.alpha_pass[5] ),
    .C(\top0.matmul0.beta_pass[4] ),
    .D(_05063_),
    .X(_05071_));
 sky130_fd_sc_hd__a21o_1 _25851_ (.A1(\top0.matmul0.beta_pass[6] ),
    .A2(_05071_),
    .B1(_05065_),
    .X(_05072_));
 sky130_fd_sc_hd__a22oi_2 _25852_ (.A1(\top0.matmul0.beta_pass[6] ),
    .A2(_05065_),
    .B1(_05072_),
    .B2(\top0.matmul0.alpha_pass[6] ),
    .Y(_05073_));
 sky130_fd_sc_hd__nor2_1 _25853_ (.A(\top0.matmul0.alpha_pass[6] ),
    .B(\top0.matmul0.beta_pass[6] ),
    .Y(_05074_));
 sky130_fd_sc_hd__a21oi_1 _25854_ (.A1(_05071_),
    .A2(_05074_),
    .B1(_05070_),
    .Y(_05075_));
 sky130_fd_sc_hd__a211o_1 _25855_ (.A1(_05070_),
    .A2(_05073_),
    .B1(_05075_),
    .C1(_02282_),
    .X(_05076_));
 sky130_fd_sc_hd__mux2_1 _25856_ (.A0(\top0.matmul0.alpha_pass[6] ),
    .A1(_05074_),
    .S(_05070_),
    .X(_05077_));
 sky130_fd_sc_hd__o31a_1 _25857_ (.A1(\top0.matmul0.alpha_pass[5] ),
    .A2(\top0.matmul0.beta_pass[5] ),
    .A3(_05438_),
    .B1(_05070_),
    .X(_05078_));
 sky130_fd_sc_hd__a211oi_1 _25858_ (.A1(_05439_),
    .A2(_05065_),
    .B1(_05078_),
    .C1(_05067_),
    .Y(_05079_));
 sky130_fd_sc_hd__a2111oi_1 _25859_ (.A1(net11),
    .A2(_05077_),
    .B1(_05079_),
    .C1(_02282_),
    .D1(_12014_),
    .Y(_05080_));
 sky130_fd_sc_hd__a22o_1 _25860_ (.A1(net888),
    .A2(_05029_),
    .B1(_05076_),
    .B2(_05080_),
    .X(_00738_));
 sky130_fd_sc_hd__inv_2 _25861_ (.A(_05070_),
    .Y(_05081_));
 sky130_fd_sc_hd__a221o_2 _25862_ (.A1(_05081_),
    .A2(_05073_),
    .B1(_05074_),
    .B2(net11),
    .C1(_05601_),
    .X(_05082_));
 sky130_fd_sc_hd__nor2_2 _25863_ (.A(\top0.matmul0.alpha_pass[7] ),
    .B(\top0.matmul0.beta_pass[7] ),
    .Y(_05083_));
 sky130_fd_sc_hd__xor2_1 _25864_ (.A(net1024),
    .B(\top0.matmul0.beta_pass[8] ),
    .X(_05084_));
 sky130_fd_sc_hd__xor2_1 _25865_ (.A(_05083_),
    .B(_05084_),
    .X(_05085_));
 sky130_fd_sc_hd__nand2_1 _25866_ (.A(_05082_),
    .B(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__or2_1 _25867_ (.A(_05082_),
    .B(_05085_),
    .X(_05087_));
 sky130_fd_sc_hd__a32o_1 _25868_ (.A1(_05031_),
    .A2(_05086_),
    .A3(_05087_),
    .B1(_05028_),
    .B2(net801),
    .X(_00739_));
 sky130_fd_sc_hd__xnor2_4 _25869_ (.A(\top0.matmul0.alpha_pass[9] ),
    .B(\top0.matmul0.beta_pass[9] ),
    .Y(_05088_));
 sky130_fd_sc_hd__nor2_1 _25870_ (.A(net1024),
    .B(\top0.matmul0.beta_pass[8] ),
    .Y(_05089_));
 sky130_fd_sc_hd__o211a_1 _25871_ (.A1(\top0.matmul0.alpha_pass[7] ),
    .A2(\top0.matmul0.beta_pass[7] ),
    .B1(\top0.matmul0.beta_pass[8] ),
    .C1(net1024),
    .X(_05090_));
 sky130_fd_sc_hd__nor3_1 _25872_ (.A(_05088_),
    .B(_05090_),
    .C(_05089_),
    .Y(_05091_));
 sky130_fd_sc_hd__a311o_1 _25873_ (.A1(_05083_),
    .A2(_05088_),
    .A3(_05089_),
    .B1(_05091_),
    .C1(_08900_),
    .X(_05092_));
 sky130_fd_sc_hd__nand2_1 _25874_ (.A(_05082_),
    .B(_05083_),
    .Y(_05093_));
 sky130_fd_sc_hd__a22o_1 _25875_ (.A1(_05083_),
    .A2(_05084_),
    .B1(_05089_),
    .B2(_05093_),
    .X(_05094_));
 sky130_fd_sc_hd__nor2_1 _25876_ (.A(_05082_),
    .B(_05083_),
    .Y(_05095_));
 sky130_fd_sc_hd__o21a_1 _25877_ (.A1(\top0.matmul0.beta_pass[8] ),
    .A2(_05095_),
    .B1(_05093_),
    .X(_05096_));
 sky130_fd_sc_hd__a22o_1 _25878_ (.A1(\top0.matmul0.beta_pass[8] ),
    .A2(_05095_),
    .B1(_05096_),
    .B2(net1024),
    .X(_05097_));
 sky130_fd_sc_hd__mux2_1 _25879_ (.A0(_05094_),
    .A1(_05097_),
    .S(_05088_),
    .X(_05098_));
 sky130_fd_sc_hd__a221o_1 _25880_ (.A1(_05082_),
    .A2(_05092_),
    .B1(_05098_),
    .B2(_05439_),
    .C1(_12014_),
    .X(_05099_));
 sky130_fd_sc_hd__a21bo_1 _25881_ (.A1(\top0.c_out_calc[9] ),
    .A2(_05029_),
    .B1_N(_05099_),
    .X(_00740_));
 sky130_fd_sc_hd__a21o_1 _25882_ (.A1(_05088_),
    .A2(_05093_),
    .B1(\top0.matmul0.beta_pass[8] ),
    .X(_05100_));
 sky130_fd_sc_hd__o21a_1 _25883_ (.A1(_05088_),
    .A2(_05095_),
    .B1(_05100_),
    .X(_05101_));
 sky130_fd_sc_hd__o221ai_4 _25884_ (.A1(_05088_),
    .A2(_05096_),
    .B1(_05101_),
    .B2(\top0.matmul0.alpha_pass[8] ),
    .C1(_05436_),
    .Y(_05102_));
 sky130_fd_sc_hd__or2_1 _25885_ (.A(\top0.matmul0.alpha_pass[9] ),
    .B(\top0.matmul0.beta_pass[9] ),
    .X(_05103_));
 sky130_fd_sc_hd__clkbuf_2 _25886_ (.A(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__xnor2_1 _25887_ (.A(\top0.matmul0.alpha_pass[10] ),
    .B(net429),
    .Y(_05105_));
 sky130_fd_sc_hd__nand2_1 _25888_ (.A(_05104_),
    .B(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__or2_1 _25889_ (.A(_05104_),
    .B(_05105_),
    .X(_05107_));
 sky130_fd_sc_hd__a21o_1 _25890_ (.A1(_05106_),
    .A2(_05107_),
    .B1(_02282_),
    .X(_05108_));
 sky130_fd_sc_hd__xnor2_1 _25891_ (.A(_05102_),
    .B(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__a2bb2o_1 _25892_ (.A1_N(_05109_),
    .A2_N(_12014_),
    .B1(net840),
    .B2(_05029_),
    .X(_00741_));
 sky130_fd_sc_hd__xor2_4 _25893_ (.A(\top0.matmul0.alpha_pass[11] ),
    .B(\top0.matmul0.beta_pass[11] ),
    .X(_05110_));
 sky130_fd_sc_hd__nand4_1 _25894_ (.A(net430),
    .B(_05438_),
    .C(_05104_),
    .D(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__o31a_1 _25895_ (.A1(\top0.matmul0.alpha_pass[10] ),
    .A2(net429),
    .A3(_05110_),
    .B1(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__or2b_1 _25896_ (.A(_05104_),
    .B_N(_05102_),
    .X(_05113_));
 sky130_fd_sc_hd__and2b_1 _25897_ (.A_N(_05102_),
    .B(_05104_),
    .X(_05114_));
 sky130_fd_sc_hd__a21o_1 _25898_ (.A1(net429),
    .A2(_05113_),
    .B1(_05114_),
    .X(_05115_));
 sky130_fd_sc_hd__a21bo_1 _25899_ (.A1(_05437_),
    .A2(_05104_),
    .B1_N(_05102_),
    .X(_05116_));
 sky130_fd_sc_hd__a21o_1 _25900_ (.A1(net429),
    .A2(_05116_),
    .B1(_05114_),
    .X(_05117_));
 sky130_fd_sc_hd__nand2_1 _25901_ (.A(_05110_),
    .B(_05117_),
    .Y(_05118_));
 sky130_fd_sc_hd__o31a_1 _25902_ (.A1(_08900_),
    .A2(_05110_),
    .A3(_05115_),
    .B1(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__inv_2 _25903_ (.A(\top0.matmul0.alpha_pass[10] ),
    .Y(_05120_));
 sky130_fd_sc_hd__nor2_1 _25904_ (.A(net429),
    .B(_05104_),
    .Y(_05121_));
 sky130_fd_sc_hd__nand3_1 _25905_ (.A(_05102_),
    .B(_05110_),
    .C(_05121_),
    .Y(_05122_));
 sky130_fd_sc_hd__a211o_1 _25906_ (.A1(net429),
    .A2(_05114_),
    .B1(_05121_),
    .C1(_05110_),
    .X(_05123_));
 sky130_fd_sc_hd__a211o_1 _25907_ (.A1(_05122_),
    .A2(_05123_),
    .B1(\top0.matmul0.alpha_pass[10] ),
    .C1(_02282_),
    .X(_05124_));
 sky130_fd_sc_hd__o221a_1 _25908_ (.A1(_05102_),
    .A2(_05112_),
    .B1(_05119_),
    .B2(_05120_),
    .C1(_05124_),
    .X(_05125_));
 sky130_fd_sc_hd__a2bb2o_1 _25909_ (.A1_N(_05125_),
    .A2_N(_12014_),
    .B1(net844),
    .B2(_05029_),
    .X(_00742_));
 sky130_fd_sc_hd__a21o_1 _25910_ (.A1(_05120_),
    .A2(_05121_),
    .B1(_05601_),
    .X(_05126_));
 sky130_fd_sc_hd__a22oi_2 _25911_ (.A1(net429),
    .A2(_05114_),
    .B1(_05115_),
    .B2(\top0.matmul0.alpha_pass[10] ),
    .Y(_05127_));
 sky130_fd_sc_hd__a22o_1 _25912_ (.A1(_05102_),
    .A2(_05126_),
    .B1(_05127_),
    .B2(_05110_),
    .X(_05128_));
 sky130_fd_sc_hd__xnor2_2 _25913_ (.A(\top0.matmul0.alpha_pass[12] ),
    .B(\top0.matmul0.beta_pass[12] ),
    .Y(_05129_));
 sky130_fd_sc_hd__nor2_1 _25914_ (.A(\top0.matmul0.alpha_pass[11] ),
    .B(\top0.matmul0.beta_pass[11] ),
    .Y(_05130_));
 sky130_fd_sc_hd__xnor2_1 _25915_ (.A(_05129_),
    .B(_05130_),
    .Y(_05131_));
 sky130_fd_sc_hd__nand2_1 _25916_ (.A(_05128_),
    .B(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__or2_1 _25917_ (.A(_05128_),
    .B(_05131_),
    .X(_05133_));
 sky130_fd_sc_hd__a32o_1 _25918_ (.A1(_05030_),
    .A2(_05132_),
    .A3(_05133_),
    .B1(_05028_),
    .B2(net939),
    .X(_00743_));
 sky130_fd_sc_hd__nor2_1 _25919_ (.A(_08899_),
    .B(_05129_),
    .Y(_05134_));
 sky130_fd_sc_hd__nand2_1 _25920_ (.A(_05436_),
    .B(_05129_),
    .Y(_05135_));
 sky130_fd_sc_hd__a31o_1 _25921_ (.A1(_05102_),
    .A2(_05126_),
    .A3(_05135_),
    .B1(_05130_),
    .X(_05136_));
 sky130_fd_sc_hd__a31o_1 _25922_ (.A1(_05110_),
    .A2(_05127_),
    .A3(_05135_),
    .B1(_05136_),
    .X(_05137_));
 sky130_fd_sc_hd__o21a_1 _25923_ (.A1(_05128_),
    .A2(_05134_),
    .B1(_05137_),
    .X(_05138_));
 sky130_fd_sc_hd__or2_1 _25924_ (.A(\top0.matmul0.alpha_pass[12] ),
    .B(\top0.matmul0.beta_pass[12] ),
    .X(_05139_));
 sky130_fd_sc_hd__xnor2_2 _25925_ (.A(\top0.matmul0.alpha_pass[13] ),
    .B(\top0.matmul0.beta_pass[13] ),
    .Y(_05140_));
 sky130_fd_sc_hd__xnor2_1 _25926_ (.A(_05139_),
    .B(_05140_),
    .Y(_05141_));
 sky130_fd_sc_hd__xnor2_1 _25927_ (.A(_05138_),
    .B(_05141_),
    .Y(_05142_));
 sky130_fd_sc_hd__a22o_1 _25928_ (.A1(net936),
    .A2(_05028_),
    .B1(_05031_),
    .B2(_05142_),
    .X(_00744_));
 sky130_fd_sc_hd__a21bo_1 _25929_ (.A1(_05437_),
    .A2(_05140_),
    .B1_N(_05138_),
    .X(_05143_));
 sky130_fd_sc_hd__nor2_1 _25930_ (.A(_08899_),
    .B(_05140_),
    .Y(_05144_));
 sky130_fd_sc_hd__o2bb2a_1 _25931_ (.A1_N(_05139_),
    .A2_N(_05143_),
    .B1(_05144_),
    .B2(_05138_),
    .X(_05145_));
 sky130_fd_sc_hd__nor2_2 _25932_ (.A(\top0.matmul0.alpha_pass[13] ),
    .B(\top0.matmul0.beta_pass[13] ),
    .Y(_05146_));
 sky130_fd_sc_hd__xor2_1 _25933_ (.A(\top0.matmul0.alpha_pass[14] ),
    .B(net428),
    .X(_05147_));
 sky130_fd_sc_hd__xnor2_1 _25934_ (.A(_05146_),
    .B(_05147_),
    .Y(_05148_));
 sky130_fd_sc_hd__xnor2_1 _25935_ (.A(_05145_),
    .B(_05148_),
    .Y(_05149_));
 sky130_fd_sc_hd__a22o_1 _25936_ (.A1(net916),
    .A2(_05028_),
    .B1(_05031_),
    .B2(_05149_),
    .X(_00745_));
 sky130_fd_sc_hd__xnor2_1 _25937_ (.A(\top0.matmul0.alpha_pass[15] ),
    .B(\top0.matmul0.beta_pass[15] ),
    .Y(_05150_));
 sky130_fd_sc_hd__nor2_1 _25938_ (.A(\top0.matmul0.alpha_pass[14] ),
    .B(net428),
    .Y(_05151_));
 sky130_fd_sc_hd__a31o_1 _25939_ (.A1(_05146_),
    .A2(_05150_),
    .A3(_05151_),
    .B1(_02282_),
    .X(_05152_));
 sky130_fd_sc_hd__a21oi_1 _25940_ (.A1(_05145_),
    .A2(_05152_),
    .B1(_12014_),
    .Y(_05153_));
 sky130_fd_sc_hd__nand2_1 _25941_ (.A(_05439_),
    .B(_05150_),
    .Y(_05154_));
 sky130_fd_sc_hd__nand2_1 _25942_ (.A(_05145_),
    .B(_05146_),
    .Y(_05155_));
 sky130_fd_sc_hd__nand2_1 _25943_ (.A(_05439_),
    .B(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__a21o_1 _25944_ (.A1(_05151_),
    .A2(_05156_),
    .B1(_05150_),
    .X(_05157_));
 sky130_fd_sc_hd__nor2_1 _25945_ (.A(_05145_),
    .B(_05146_),
    .Y(_05158_));
 sky130_fd_sc_hd__a21o_1 _25946_ (.A1(net428),
    .A2(_05155_),
    .B1(_05158_),
    .X(_05159_));
 sky130_fd_sc_hd__a22oi_1 _25947_ (.A1(net428),
    .A2(_05158_),
    .B1(_05159_),
    .B2(\top0.matmul0.alpha_pass[14] ),
    .Y(_05160_));
 sky130_fd_sc_hd__mux2_1 _25948_ (.A0(_05154_),
    .A1(_05157_),
    .S(_05160_),
    .X(_05161_));
 sky130_fd_sc_hd__a22o_1 _25949_ (.A1(net921),
    .A2(_05028_),
    .B1(_05153_),
    .B2(_05161_),
    .X(_00746_));
 sky130_fd_sc_hd__o21ai_1 _25950_ (.A1(net207),
    .A2(_05015_),
    .B1(_12016_),
    .Y(_05162_));
 sky130_fd_sc_hd__and3_1 _25951_ (.A(_12025_),
    .B(_12010_),
    .C(_12014_),
    .X(_05163_));
 sky130_fd_sc_hd__buf_2 _25952_ (.A(_05163_),
    .X(_05164_));
 sky130_fd_sc_hd__clkbuf_4 _25953_ (.A(_05164_),
    .X(_05165_));
 sky130_fd_sc_hd__mux2_1 _25954_ (.A0(\top0.matmul0.op_in[0] ),
    .A1(_05162_),
    .S(_05165_),
    .X(_05166_));
 sky130_fd_sc_hd__clkbuf_1 _25955_ (.A(_05166_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _25956_ (.A0(\top0.matmul0.op_in[1] ),
    .A1(_12015_),
    .S(_05165_),
    .X(_05167_));
 sky130_fd_sc_hd__clkbuf_1 _25957_ (.A(_05167_),
    .X(_00748_));
 sky130_fd_sc_hd__a211oi_4 _25958_ (.A1(_12030_),
    .A2(_05015_),
    .B1(net207),
    .C1(_08900_),
    .Y(_05168_));
 sky130_fd_sc_hd__buf_2 _25959_ (.A(_05168_),
    .X(_05169_));
 sky130_fd_sc_hd__a22o_1 _25960_ (.A1(\top0.pid_q.out[0] ),
    .A2(_12032_),
    .B1(_05014_),
    .B2(\spi0.data_packed[48] ),
    .X(_05170_));
 sky130_fd_sc_hd__a21o_1 _25961_ (.A1(\top0.matmul0.beta_pass[0] ),
    .A2(_05169_),
    .B1(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__mux2_1 _25962_ (.A0(\top0.b_in_matmul[0] ),
    .A1(_05171_),
    .S(_05165_),
    .X(_05172_));
 sky130_fd_sc_hd__clkbuf_1 _25963_ (.A(_05172_),
    .X(_00749_));
 sky130_fd_sc_hd__a22o_1 _25964_ (.A1(\top0.pid_q.out[1] ),
    .A2(_12032_),
    .B1(_05014_),
    .B2(\spi0.data_packed[49] ),
    .X(_05173_));
 sky130_fd_sc_hd__a21o_1 _25965_ (.A1(\top0.matmul0.beta_pass[1] ),
    .A2(_05169_),
    .B1(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__mux2_1 _25966_ (.A0(net998),
    .A1(_05174_),
    .S(_05165_),
    .X(_05175_));
 sky130_fd_sc_hd__clkbuf_1 _25967_ (.A(_05175_),
    .X(_00750_));
 sky130_fd_sc_hd__a22o_1 _25968_ (.A1(\top0.pid_q.out[2] ),
    .A2(_12032_),
    .B1(_05014_),
    .B2(\spi0.data_packed[50] ),
    .X(_05176_));
 sky130_fd_sc_hd__a21o_1 _25969_ (.A1(\top0.matmul0.beta_pass[2] ),
    .A2(_05169_),
    .B1(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__mux2_1 _25970_ (.A0(\top0.b_in_matmul[2] ),
    .A1(_05177_),
    .S(_05165_),
    .X(_05178_));
 sky130_fd_sc_hd__clkbuf_1 _25971_ (.A(_05178_),
    .X(_00751_));
 sky130_fd_sc_hd__a22o_1 _25972_ (.A1(\top0.pid_q.out[3] ),
    .A2(_12032_),
    .B1(_05014_),
    .B2(\spi0.data_packed[51] ),
    .X(_05179_));
 sky130_fd_sc_hd__a21o_1 _25973_ (.A1(\top0.matmul0.beta_pass[3] ),
    .A2(_05169_),
    .B1(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__mux2_1 _25974_ (.A0(\top0.b_in_matmul[3] ),
    .A1(_05180_),
    .S(_05165_),
    .X(_05181_));
 sky130_fd_sc_hd__clkbuf_1 _25975_ (.A(_05181_),
    .X(_00752_));
 sky130_fd_sc_hd__a22o_1 _25976_ (.A1(\top0.pid_q.out[4] ),
    .A2(_12032_),
    .B1(_05014_),
    .B2(\spi0.data_packed[52] ),
    .X(_05182_));
 sky130_fd_sc_hd__a21o_1 _25977_ (.A1(\top0.matmul0.beta_pass[4] ),
    .A2(_05169_),
    .B1(_05182_),
    .X(_05183_));
 sky130_fd_sc_hd__mux2_1 _25978_ (.A0(\top0.b_in_matmul[4] ),
    .A1(_05183_),
    .S(_05165_),
    .X(_05184_));
 sky130_fd_sc_hd__clkbuf_1 _25979_ (.A(_05184_),
    .X(_00753_));
 sky130_fd_sc_hd__a22o_1 _25980_ (.A1(\top0.pid_q.out[5] ),
    .A2(_12032_),
    .B1(_05014_),
    .B2(\spi0.data_packed[53] ),
    .X(_05185_));
 sky130_fd_sc_hd__a21o_1 _25981_ (.A1(\top0.matmul0.beta_pass[5] ),
    .A2(_05169_),
    .B1(_05185_),
    .X(_05186_));
 sky130_fd_sc_hd__mux2_1 _25982_ (.A0(net1004),
    .A1(_05186_),
    .S(_05165_),
    .X(_05187_));
 sky130_fd_sc_hd__clkbuf_1 _25983_ (.A(_05187_),
    .X(_00754_));
 sky130_fd_sc_hd__a22o_1 _25984_ (.A1(\top0.pid_q.out[6] ),
    .A2(_12032_),
    .B1(_05014_),
    .B2(\spi0.data_packed[54] ),
    .X(_05188_));
 sky130_fd_sc_hd__a21o_1 _25985_ (.A1(\top0.matmul0.beta_pass[6] ),
    .A2(_05169_),
    .B1(_05188_),
    .X(_05189_));
 sky130_fd_sc_hd__mux2_1 _25986_ (.A0(net966),
    .A1(_05189_),
    .S(_05165_),
    .X(_05190_));
 sky130_fd_sc_hd__clkbuf_1 _25987_ (.A(_05190_),
    .X(_00755_));
 sky130_fd_sc_hd__a22o_1 _25988_ (.A1(\top0.pid_q.out[7] ),
    .A2(_12032_),
    .B1(_05014_),
    .B2(\spi0.data_packed[55] ),
    .X(_05191_));
 sky130_fd_sc_hd__a21o_1 _25989_ (.A1(\top0.matmul0.beta_pass[7] ),
    .A2(_05169_),
    .B1(_05191_),
    .X(_05192_));
 sky130_fd_sc_hd__mux2_1 _25990_ (.A0(\top0.b_in_matmul[7] ),
    .A1(_05192_),
    .S(_05165_),
    .X(_05193_));
 sky130_fd_sc_hd__clkbuf_1 _25991_ (.A(_05193_),
    .X(_00756_));
 sky130_fd_sc_hd__a22o_1 _25992_ (.A1(\top0.pid_q.out[8] ),
    .A2(_12032_),
    .B1(_05014_),
    .B2(\spi0.data_packed[56] ),
    .X(_05194_));
 sky130_fd_sc_hd__a21o_1 _25993_ (.A1(\top0.matmul0.beta_pass[8] ),
    .A2(_05169_),
    .B1(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__buf_4 _25994_ (.A(_05164_),
    .X(_05196_));
 sky130_fd_sc_hd__mux2_1 _25995_ (.A0(\top0.b_in_matmul[8] ),
    .A1(_05195_),
    .S(_05196_),
    .X(_05197_));
 sky130_fd_sc_hd__clkbuf_1 _25996_ (.A(_05197_),
    .X(_00757_));
 sky130_fd_sc_hd__clkbuf_4 _25997_ (.A(_12031_),
    .X(_05198_));
 sky130_fd_sc_hd__clkbuf_4 _25998_ (.A(_05013_),
    .X(_05199_));
 sky130_fd_sc_hd__a22o_1 _25999_ (.A1(\top0.pid_q.out[9] ),
    .A2(_05198_),
    .B1(_05199_),
    .B2(\spi0.data_packed[57] ),
    .X(_05200_));
 sky130_fd_sc_hd__a21o_1 _26000_ (.A1(\top0.matmul0.beta_pass[9] ),
    .A2(_05169_),
    .B1(_05200_),
    .X(_05201_));
 sky130_fd_sc_hd__mux2_1 _26001_ (.A0(\top0.b_in_matmul[9] ),
    .A1(_05201_),
    .S(_05196_),
    .X(_05202_));
 sky130_fd_sc_hd__clkbuf_1 _26002_ (.A(_05202_),
    .X(_00758_));
 sky130_fd_sc_hd__buf_2 _26003_ (.A(_05168_),
    .X(_05203_));
 sky130_fd_sc_hd__a22o_1 _26004_ (.A1(\top0.pid_q.out[10] ),
    .A2(_05198_),
    .B1(_05199_),
    .B2(\spi0.data_packed[58] ),
    .X(_05204_));
 sky130_fd_sc_hd__a21o_1 _26005_ (.A1(net430),
    .A2(_05203_),
    .B1(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__mux2_1 _26006_ (.A0(\top0.b_in_matmul[10] ),
    .A1(_05205_),
    .S(_05196_),
    .X(_05206_));
 sky130_fd_sc_hd__clkbuf_1 _26007_ (.A(_05206_),
    .X(_00759_));
 sky130_fd_sc_hd__a22o_1 _26008_ (.A1(\top0.pid_q.out[11] ),
    .A2(_05198_),
    .B1(_05199_),
    .B2(\spi0.data_packed[59] ),
    .X(_05207_));
 sky130_fd_sc_hd__a21o_1 _26009_ (.A1(\top0.matmul0.beta_pass[11] ),
    .A2(_05203_),
    .B1(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__mux2_1 _26010_ (.A0(net980),
    .A1(_05208_),
    .S(_05196_),
    .X(_05209_));
 sky130_fd_sc_hd__clkbuf_1 _26011_ (.A(_05209_),
    .X(_00760_));
 sky130_fd_sc_hd__a22o_1 _26012_ (.A1(\top0.pid_q.out[12] ),
    .A2(_05198_),
    .B1(_05199_),
    .B2(\spi0.data_packed[60] ),
    .X(_05210_));
 sky130_fd_sc_hd__a21o_1 _26013_ (.A1(\top0.matmul0.beta_pass[12] ),
    .A2(_05203_),
    .B1(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__mux2_1 _26014_ (.A0(\top0.b_in_matmul[12] ),
    .A1(_05211_),
    .S(_05196_),
    .X(_05212_));
 sky130_fd_sc_hd__clkbuf_1 _26015_ (.A(_05212_),
    .X(_00761_));
 sky130_fd_sc_hd__a22o_1 _26016_ (.A1(\top0.pid_q.out[13] ),
    .A2(_05198_),
    .B1(_05199_),
    .B2(\spi0.data_packed[61] ),
    .X(_05213_));
 sky130_fd_sc_hd__a21o_1 _26017_ (.A1(\top0.matmul0.beta_pass[13] ),
    .A2(_05203_),
    .B1(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__mux2_1 _26018_ (.A0(\top0.b_in_matmul[13] ),
    .A1(_05214_),
    .S(_05196_),
    .X(_05215_));
 sky130_fd_sc_hd__clkbuf_1 _26019_ (.A(_05215_),
    .X(_00762_));
 sky130_fd_sc_hd__a22o_1 _26020_ (.A1(\top0.pid_q.out[14] ),
    .A2(_05198_),
    .B1(_05199_),
    .B2(\spi0.data_packed[62] ),
    .X(_05216_));
 sky130_fd_sc_hd__a21o_1 _26021_ (.A1(net428),
    .A2(_05203_),
    .B1(_05216_),
    .X(_05217_));
 sky130_fd_sc_hd__mux2_1 _26022_ (.A0(net994),
    .A1(_05217_),
    .S(_05196_),
    .X(_05218_));
 sky130_fd_sc_hd__clkbuf_1 _26023_ (.A(_05218_),
    .X(_00763_));
 sky130_fd_sc_hd__a22o_1 _26024_ (.A1(\top0.pid_q.out[15] ),
    .A2(_05198_),
    .B1(_05199_),
    .B2(\spi0.data_packed[63] ),
    .X(_05219_));
 sky130_fd_sc_hd__a21o_1 _26025_ (.A1(\top0.matmul0.beta_pass[15] ),
    .A2(_05203_),
    .B1(_05219_),
    .X(_05220_));
 sky130_fd_sc_hd__mux2_1 _26026_ (.A0(\top0.b_in_matmul[15] ),
    .A1(_05220_),
    .S(_05196_),
    .X(_05221_));
 sky130_fd_sc_hd__clkbuf_1 _26027_ (.A(_05221_),
    .X(_00764_));
 sky130_fd_sc_hd__a22o_1 _26028_ (.A1(\top0.pid_d.out[0] ),
    .A2(_05198_),
    .B1(_05199_),
    .B2(\spi0.data_packed[64] ),
    .X(_05222_));
 sky130_fd_sc_hd__a21o_1 _26029_ (.A1(\top0.matmul0.alpha_pass[0] ),
    .A2(_05203_),
    .B1(_05222_),
    .X(_05223_));
 sky130_fd_sc_hd__mux2_1 _26030_ (.A0(\top0.a_in_matmul[0] ),
    .A1(_05223_),
    .S(_05196_),
    .X(_05224_));
 sky130_fd_sc_hd__clkbuf_1 _26031_ (.A(_05224_),
    .X(_00765_));
 sky130_fd_sc_hd__a22o_1 _26032_ (.A1(\top0.pid_d.out[1] ),
    .A2(_05198_),
    .B1(_05199_),
    .B2(\spi0.data_packed[65] ),
    .X(_05225_));
 sky130_fd_sc_hd__a21o_1 _26033_ (.A1(\top0.matmul0.alpha_pass[1] ),
    .A2(_05203_),
    .B1(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__mux2_1 _26034_ (.A0(\top0.a_in_matmul[1] ),
    .A1(_05226_),
    .S(_05196_),
    .X(_05227_));
 sky130_fd_sc_hd__clkbuf_1 _26035_ (.A(_05227_),
    .X(_00766_));
 sky130_fd_sc_hd__a22o_1 _26036_ (.A1(\top0.pid_d.out[2] ),
    .A2(_05198_),
    .B1(_05199_),
    .B2(\spi0.data_packed[66] ),
    .X(_05228_));
 sky130_fd_sc_hd__a21o_1 _26037_ (.A1(\top0.matmul0.alpha_pass[2] ),
    .A2(_05203_),
    .B1(_05228_),
    .X(_05229_));
 sky130_fd_sc_hd__clkbuf_4 _26038_ (.A(_05164_),
    .X(_05230_));
 sky130_fd_sc_hd__mux2_1 _26039_ (.A0(net979),
    .A1(_05229_),
    .S(_05230_),
    .X(_05231_));
 sky130_fd_sc_hd__clkbuf_1 _26040_ (.A(_05231_),
    .X(_00767_));
 sky130_fd_sc_hd__buf_2 _26041_ (.A(_12031_),
    .X(_05232_));
 sky130_fd_sc_hd__buf_2 _26042_ (.A(_05013_),
    .X(_05233_));
 sky130_fd_sc_hd__a22o_1 _26043_ (.A1(\top0.pid_d.out[3] ),
    .A2(_05232_),
    .B1(_05233_),
    .B2(\spi0.data_packed[67] ),
    .X(_05234_));
 sky130_fd_sc_hd__a21o_1 _26044_ (.A1(\top0.matmul0.alpha_pass[3] ),
    .A2(_05203_),
    .B1(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__mux2_1 _26045_ (.A0(\top0.a_in_matmul[3] ),
    .A1(_05235_),
    .S(_05230_),
    .X(_05236_));
 sky130_fd_sc_hd__clkbuf_1 _26046_ (.A(_05236_),
    .X(_00768_));
 sky130_fd_sc_hd__buf_2 _26047_ (.A(_05168_),
    .X(_05237_));
 sky130_fd_sc_hd__a22o_1 _26048_ (.A1(\top0.pid_d.out[4] ),
    .A2(_05232_),
    .B1(_05233_),
    .B2(\spi0.data_packed[68] ),
    .X(_05238_));
 sky130_fd_sc_hd__a21o_1 _26049_ (.A1(\top0.matmul0.alpha_pass[4] ),
    .A2(_05237_),
    .B1(_05238_),
    .X(_05239_));
 sky130_fd_sc_hd__mux2_1 _26050_ (.A0(\top0.a_in_matmul[4] ),
    .A1(_05239_),
    .S(_05230_),
    .X(_05240_));
 sky130_fd_sc_hd__clkbuf_1 _26051_ (.A(_05240_),
    .X(_00769_));
 sky130_fd_sc_hd__a22o_1 _26052_ (.A1(\top0.pid_d.out[5] ),
    .A2(_05232_),
    .B1(_05233_),
    .B2(\spi0.data_packed[69] ),
    .X(_05241_));
 sky130_fd_sc_hd__a21o_1 _26053_ (.A1(net76),
    .A2(_05237_),
    .B1(_05241_),
    .X(_05242_));
 sky130_fd_sc_hd__mux2_1 _26054_ (.A0(\top0.a_in_matmul[5] ),
    .A1(_05242_),
    .S(_05230_),
    .X(_05243_));
 sky130_fd_sc_hd__clkbuf_1 _26055_ (.A(_05243_),
    .X(_00770_));
 sky130_fd_sc_hd__a22o_1 _26056_ (.A1(\top0.pid_d.out[6] ),
    .A2(_05232_),
    .B1(_05233_),
    .B2(\spi0.data_packed[70] ),
    .X(_05244_));
 sky130_fd_sc_hd__a21o_1 _26057_ (.A1(\top0.matmul0.alpha_pass[6] ),
    .A2(_05237_),
    .B1(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__mux2_1 _26058_ (.A0(\top0.a_in_matmul[6] ),
    .A1(_05245_),
    .S(_05230_),
    .X(_05246_));
 sky130_fd_sc_hd__clkbuf_1 _26059_ (.A(_05246_),
    .X(_00771_));
 sky130_fd_sc_hd__a22o_1 _26060_ (.A1(\top0.pid_d.out[7] ),
    .A2(_05232_),
    .B1(_05233_),
    .B2(\spi0.data_packed[71] ),
    .X(_05247_));
 sky130_fd_sc_hd__a21o_1 _26061_ (.A1(\top0.matmul0.alpha_pass[7] ),
    .A2(_05237_),
    .B1(_05247_),
    .X(_05248_));
 sky130_fd_sc_hd__mux2_1 _26062_ (.A0(\top0.a_in_matmul[7] ),
    .A1(_05248_),
    .S(_05230_),
    .X(_05249_));
 sky130_fd_sc_hd__clkbuf_1 _26063_ (.A(_05249_),
    .X(_00772_));
 sky130_fd_sc_hd__a22o_1 _26064_ (.A1(\top0.pid_d.out[8] ),
    .A2(_05232_),
    .B1(_05233_),
    .B2(\spi0.data_packed[72] ),
    .X(_05250_));
 sky130_fd_sc_hd__a21o_1 _26065_ (.A1(net1024),
    .A2(_05237_),
    .B1(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__mux2_1 _26066_ (.A0(net985),
    .A1(_05251_),
    .S(_05230_),
    .X(_05252_));
 sky130_fd_sc_hd__clkbuf_1 _26067_ (.A(_05252_),
    .X(_00773_));
 sky130_fd_sc_hd__a22o_1 _26068_ (.A1(\top0.pid_d.out[9] ),
    .A2(_05232_),
    .B1(_05233_),
    .B2(\spi0.data_packed[73] ),
    .X(_05253_));
 sky130_fd_sc_hd__a21o_1 _26069_ (.A1(\top0.matmul0.alpha_pass[9] ),
    .A2(_05237_),
    .B1(_05253_),
    .X(_05254_));
 sky130_fd_sc_hd__mux2_1 _26070_ (.A0(\top0.a_in_matmul[9] ),
    .A1(_05254_),
    .S(_05230_),
    .X(_05255_));
 sky130_fd_sc_hd__clkbuf_1 _26071_ (.A(_05255_),
    .X(_00774_));
 sky130_fd_sc_hd__a22o_1 _26072_ (.A1(\top0.pid_d.out[10] ),
    .A2(_05232_),
    .B1(_05233_),
    .B2(\spi0.data_packed[74] ),
    .X(_05256_));
 sky130_fd_sc_hd__a21o_1 _26073_ (.A1(\top0.matmul0.alpha_pass[10] ),
    .A2(_05237_),
    .B1(_05256_),
    .X(_05257_));
 sky130_fd_sc_hd__mux2_1 _26074_ (.A0(\top0.a_in_matmul[10] ),
    .A1(_05257_),
    .S(_05230_),
    .X(_05258_));
 sky130_fd_sc_hd__clkbuf_1 _26075_ (.A(_05258_),
    .X(_00775_));
 sky130_fd_sc_hd__a22o_1 _26076_ (.A1(\top0.pid_d.out[11] ),
    .A2(_05232_),
    .B1(_05233_),
    .B2(\spi0.data_packed[75] ),
    .X(_05259_));
 sky130_fd_sc_hd__a21o_1 _26077_ (.A1(\top0.matmul0.alpha_pass[11] ),
    .A2(_05237_),
    .B1(_05259_),
    .X(_05260_));
 sky130_fd_sc_hd__mux2_1 _26078_ (.A0(\top0.a_in_matmul[11] ),
    .A1(_05260_),
    .S(_05230_),
    .X(_05261_));
 sky130_fd_sc_hd__clkbuf_1 _26079_ (.A(_05261_),
    .X(_00776_));
 sky130_fd_sc_hd__a22o_1 _26080_ (.A1(\top0.pid_d.out[12] ),
    .A2(_05232_),
    .B1(_05233_),
    .B2(\spi0.data_packed[76] ),
    .X(_05262_));
 sky130_fd_sc_hd__a21o_1 _26081_ (.A1(\top0.matmul0.alpha_pass[12] ),
    .A2(_05237_),
    .B1(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__mux2_1 _26082_ (.A0(\top0.a_in_matmul[12] ),
    .A1(_05263_),
    .S(_05164_),
    .X(_05264_));
 sky130_fd_sc_hd__clkbuf_1 _26083_ (.A(_05264_),
    .X(_00777_));
 sky130_fd_sc_hd__a22o_1 _26084_ (.A1(\top0.pid_d.out[13] ),
    .A2(_12031_),
    .B1(_05013_),
    .B2(\spi0.data_packed[77] ),
    .X(_05265_));
 sky130_fd_sc_hd__a21o_1 _26085_ (.A1(\top0.matmul0.alpha_pass[13] ),
    .A2(_05237_),
    .B1(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__mux2_1 _26086_ (.A0(\top0.a_in_matmul[13] ),
    .A1(_05266_),
    .S(_05164_),
    .X(_05267_));
 sky130_fd_sc_hd__clkbuf_1 _26087_ (.A(_05267_),
    .X(_00778_));
 sky130_fd_sc_hd__a22o_1 _26088_ (.A1(\top0.pid_d.out[14] ),
    .A2(_12031_),
    .B1(_05013_),
    .B2(\spi0.data_packed[78] ),
    .X(_05268_));
 sky130_fd_sc_hd__a21o_1 _26089_ (.A1(\top0.matmul0.alpha_pass[14] ),
    .A2(_05168_),
    .B1(_05268_),
    .X(_05269_));
 sky130_fd_sc_hd__mux2_1 _26090_ (.A0(\top0.a_in_matmul[14] ),
    .A1(_05269_),
    .S(_05164_),
    .X(_05270_));
 sky130_fd_sc_hd__clkbuf_1 _26091_ (.A(_05270_),
    .X(_00779_));
 sky130_fd_sc_hd__a22o_1 _26092_ (.A1(\top0.pid_d.out[15] ),
    .A2(_12031_),
    .B1(_05013_),
    .B2(\spi0.data_packed[79] ),
    .X(_05271_));
 sky130_fd_sc_hd__a21o_1 _26093_ (.A1(\top0.matmul0.alpha_pass[15] ),
    .A2(_05168_),
    .B1(_05271_),
    .X(_05272_));
 sky130_fd_sc_hd__mux2_1 _26094_ (.A0(\top0.a_in_matmul[15] ),
    .A1(_05272_),
    .S(_05164_),
    .X(_05273_));
 sky130_fd_sc_hd__clkbuf_1 _26095_ (.A(_05273_),
    .X(_00780_));
 sky130_fd_sc_hd__and2_1 _26096_ (.A(_05426_),
    .B(_05013_),
    .X(_05274_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _26097_ (.A(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__buf_2 _26098_ (.A(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__o22a_2 _26099_ (.A1(_12017_),
    .A2(_12019_),
    .B1(_12012_),
    .B2(_12009_),
    .X(_05277_));
 sky130_fd_sc_hd__buf_2 _26100_ (.A(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__a22o_1 _26101_ (.A1(\top0.periodTop[0] ),
    .A2(_05276_),
    .B1(_05278_),
    .B2(net68),
    .X(_00781_));
 sky130_fd_sc_hd__a22o_1 _26102_ (.A1(\top0.periodTop[1] ),
    .A2(_05276_),
    .B1(_05278_),
    .B2(net62),
    .X(_00782_));
 sky130_fd_sc_hd__a22o_1 _26103_ (.A1(\top0.periodTop[2] ),
    .A2(_05276_),
    .B1(_05278_),
    .B2(net59),
    .X(_00783_));
 sky130_fd_sc_hd__a22o_1 _26104_ (.A1(net782),
    .A2(_05276_),
    .B1(_05278_),
    .B2(net58),
    .X(_00784_));
 sky130_fd_sc_hd__a22o_1 _26105_ (.A1(net741),
    .A2(_05276_),
    .B1(_05278_),
    .B2(net1025),
    .X(_00785_));
 sky130_fd_sc_hd__a22o_1 _26106_ (.A1(net845),
    .A2(_05276_),
    .B1(_05278_),
    .B2(net1027),
    .X(_00786_));
 sky130_fd_sc_hd__a22o_1 _26107_ (.A1(\top0.periodTop[6] ),
    .A2(_05276_),
    .B1(_05278_),
    .B2(net50),
    .X(_00787_));
 sky130_fd_sc_hd__a22o_1 _26108_ (.A1(\top0.periodTop[7] ),
    .A2(_05276_),
    .B1(_05278_),
    .B2(net47),
    .X(_00788_));
 sky130_fd_sc_hd__a22o_1 _26109_ (.A1(\top0.periodTop[8] ),
    .A2(_05276_),
    .B1(_05278_),
    .B2(net43),
    .X(_00789_));
 sky130_fd_sc_hd__a22o_1 _26110_ (.A1(\top0.periodTop[9] ),
    .A2(_05276_),
    .B1(_05278_),
    .B2(net42),
    .X(_00790_));
 sky130_fd_sc_hd__clkbuf_4 _26111_ (.A(_05275_),
    .X(_05279_));
 sky130_fd_sc_hd__clkbuf_4 _26112_ (.A(_05277_),
    .X(_05280_));
 sky130_fd_sc_hd__a22o_1 _26113_ (.A1(net900),
    .A2(_05279_),
    .B1(_05280_),
    .B2(net40),
    .X(_00791_));
 sky130_fd_sc_hd__a22o_1 _26114_ (.A1(net832),
    .A2(_05279_),
    .B1(_05280_),
    .B2(net38),
    .X(_00792_));
 sky130_fd_sc_hd__a22o_1 _26115_ (.A1(net895),
    .A2(_05279_),
    .B1(_05280_),
    .B2(net35),
    .X(_00793_));
 sky130_fd_sc_hd__a22o_1 _26116_ (.A1(net886),
    .A2(_05279_),
    .B1(_05280_),
    .B2(net32),
    .X(_00794_));
 sky130_fd_sc_hd__a22o_1 _26117_ (.A1(net754),
    .A2(_05279_),
    .B1(_05280_),
    .B2(net1030),
    .X(_00795_));
 sky130_fd_sc_hd__a22o_1 _26118_ (.A1(net737),
    .A2(_05279_),
    .B1(_05280_),
    .B2(net24),
    .X(_00796_));
 sky130_fd_sc_hd__a22o_1 _26119_ (.A1(\spi0.data_packed[16] ),
    .A2(_05279_),
    .B1(_05280_),
    .B2(net907),
    .X(_00797_));
 sky130_fd_sc_hd__a22o_1 _26120_ (.A1(\spi0.data_packed[17] ),
    .A2(_05279_),
    .B1(_05280_),
    .B2(net919),
    .X(_00798_));
 sky130_fd_sc_hd__a22o_1 _26121_ (.A1(\spi0.data_packed[18] ),
    .A2(_05279_),
    .B1(_05280_),
    .B2(\top0.currT_r[2] ),
    .X(_00799_));
 sky130_fd_sc_hd__a22o_1 _26122_ (.A1(\spi0.data_packed[19] ),
    .A2(_05279_),
    .B1(_05280_),
    .B2(net934),
    .X(_00800_));
 sky130_fd_sc_hd__clkbuf_4 _26123_ (.A(_05275_),
    .X(_05281_));
 sky130_fd_sc_hd__clkbuf_4 _26124_ (.A(_05277_),
    .X(_05282_));
 sky130_fd_sc_hd__a22o_1 _26125_ (.A1(\spi0.data_packed[20] ),
    .A2(_05281_),
    .B1(_05282_),
    .B2(net918),
    .X(_00801_));
 sky130_fd_sc_hd__a22o_1 _26126_ (.A1(\spi0.data_packed[21] ),
    .A2(_05281_),
    .B1(_05282_),
    .B2(net905),
    .X(_00802_));
 sky130_fd_sc_hd__a22o_1 _26127_ (.A1(\spi0.data_packed[22] ),
    .A2(_05281_),
    .B1(_05282_),
    .B2(net960),
    .X(_00803_));
 sky130_fd_sc_hd__a22o_1 _26128_ (.A1(\spi0.data_packed[23] ),
    .A2(_05281_),
    .B1(_05282_),
    .B2(net962),
    .X(_00804_));
 sky130_fd_sc_hd__a22o_1 _26129_ (.A1(\spi0.data_packed[24] ),
    .A2(_05281_),
    .B1(_05282_),
    .B2(net948),
    .X(_00805_));
 sky130_fd_sc_hd__a22o_1 _26130_ (.A1(\spi0.data_packed[25] ),
    .A2(_05281_),
    .B1(_05282_),
    .B2(net952),
    .X(_00806_));
 sky130_fd_sc_hd__a22o_1 _26131_ (.A1(\spi0.data_packed[26] ),
    .A2(_05281_),
    .B1(_05282_),
    .B2(\top0.currT_r[10] ),
    .X(_00807_));
 sky130_fd_sc_hd__a22o_1 _26132_ (.A1(\spi0.data_packed[27] ),
    .A2(_05281_),
    .B1(_05282_),
    .B2(net935),
    .X(_00808_));
 sky130_fd_sc_hd__a22o_1 _26133_ (.A1(\spi0.data_packed[28] ),
    .A2(_05281_),
    .B1(_05282_),
    .B2(net922),
    .X(_00809_));
 sky130_fd_sc_hd__a22o_1 _26134_ (.A1(\spi0.data_packed[29] ),
    .A2(_05281_),
    .B1(_05282_),
    .B2(\top0.currT_r[13] ),
    .X(_00810_));
 sky130_fd_sc_hd__a22o_1 _26135_ (.A1(\spi0.data_packed[30] ),
    .A2(_05275_),
    .B1(_05277_),
    .B2(\top0.currT_r[14] ),
    .X(_00811_));
 sky130_fd_sc_hd__a22o_1 _26136_ (.A1(\spi0.data_packed[31] ),
    .A2(_05275_),
    .B1(_05277_),
    .B2(net802),
    .X(_00812_));
 sky130_fd_sc_hd__nor2_1 _26137_ (.A(net18),
    .B(\spi0.data_packed[15] ),
    .Y(_05283_));
 sky130_fd_sc_hd__xnor2_1 _26138_ (.A(\spi0.data_packed[0] ),
    .B(_05283_),
    .Y(_05284_));
 sky130_fd_sc_hd__mux2_1 _26139_ (.A0(_05284_),
    .A1(\top0.cordic0.slte0.opB[2] ),
    .S(_12006_),
    .X(_05285_));
 sky130_fd_sc_hd__clkbuf_1 _26140_ (.A(_05285_),
    .X(_00813_));
 sky130_fd_sc_hd__a21oi_1 _26141_ (.A1(\spi0.data_packed[0] ),
    .A2(\spi0.data_packed[15] ),
    .B1(net19),
    .Y(_05286_));
 sky130_fd_sc_hd__xnor2_1 _26142_ (.A(\spi0.data_packed[1] ),
    .B(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__mux2_1 _26143_ (.A0(_05287_),
    .A1(\top0.cordic0.slte0.opB[3] ),
    .S(_12006_),
    .X(_05288_));
 sky130_fd_sc_hd__clkbuf_1 _26144_ (.A(_05288_),
    .X(_00814_));
 sky130_fd_sc_hd__a31o_1 _26145_ (.A1(\spi0.data_packed[0] ),
    .A2(\spi0.data_packed[15] ),
    .A3(\spi0.data_packed[1] ),
    .B1(net19),
    .X(_05289_));
 sky130_fd_sc_hd__xor2_1 _26146_ (.A(\spi0.data_packed[2] ),
    .B(_05289_),
    .X(_05290_));
 sky130_fd_sc_hd__mux2_1 _26147_ (.A0(_05290_),
    .A1(\top0.cordic0.slte0.opB[4] ),
    .S(_12006_),
    .X(_05291_));
 sky130_fd_sc_hd__clkbuf_1 _26148_ (.A(_05291_),
    .X(_00815_));
 sky130_fd_sc_hd__and4_1 _26149_ (.A(\spi0.data_packed[0] ),
    .B(\spi0.data_packed[15] ),
    .C(\spi0.data_packed[1] ),
    .D(\spi0.data_packed[2] ),
    .X(_05292_));
 sky130_fd_sc_hd__nor2_1 _26150_ (.A(net18),
    .B(_05292_),
    .Y(_05293_));
 sky130_fd_sc_hd__xnor2_1 _26151_ (.A(\spi0.data_packed[3] ),
    .B(_05293_),
    .Y(_05294_));
 sky130_fd_sc_hd__mux2_1 _26152_ (.A0(_05294_),
    .A1(\top0.cordic0.slte0.opB[5] ),
    .S(_12006_),
    .X(_05295_));
 sky130_fd_sc_hd__clkbuf_1 _26153_ (.A(_05295_),
    .X(_00816_));
 sky130_fd_sc_hd__a21oi_1 _26154_ (.A1(\spi0.data_packed[3] ),
    .A2(_05292_),
    .B1(net18),
    .Y(_05296_));
 sky130_fd_sc_hd__xnor2_1 _26155_ (.A(\spi0.data_packed[4] ),
    .B(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__mux2_1 _26156_ (.A0(_05297_),
    .A1(\top0.cordic0.slte0.opB[6] ),
    .S(_12006_),
    .X(_05298_));
 sky130_fd_sc_hd__clkbuf_1 _26157_ (.A(_05298_),
    .X(_00817_));
 sky130_fd_sc_hd__and3_1 _26158_ (.A(\spi0.data_packed[3] ),
    .B(\spi0.data_packed[4] ),
    .C(_05292_),
    .X(_05299_));
 sky130_fd_sc_hd__nor2_1 _26159_ (.A(net18),
    .B(_05299_),
    .Y(_05300_));
 sky130_fd_sc_hd__xnor2_1 _26160_ (.A(\spi0.data_packed[5] ),
    .B(_05300_),
    .Y(_05301_));
 sky130_fd_sc_hd__mux2_1 _26161_ (.A0(_05301_),
    .A1(\top0.cordic0.slte0.opB[7] ),
    .S(_12006_),
    .X(_05302_));
 sky130_fd_sc_hd__clkbuf_1 _26162_ (.A(_05302_),
    .X(_00818_));
 sky130_fd_sc_hd__and2_1 _26163_ (.A(\spi0.data_packed[5] ),
    .B(_05299_),
    .X(_05303_));
 sky130_fd_sc_hd__nor2_1 _26164_ (.A(net18),
    .B(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__xnor2_1 _26165_ (.A(\spi0.data_packed[6] ),
    .B(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__mux2_1 _26166_ (.A0(_05305_),
    .A1(\top0.cordic0.slte0.opB[8] ),
    .S(_12006_),
    .X(_05306_));
 sky130_fd_sc_hd__clkbuf_1 _26167_ (.A(_05306_),
    .X(_00819_));
 sky130_fd_sc_hd__a31o_1 _26168_ (.A1(\spi0.data_packed[5] ),
    .A2(\spi0.data_packed[6] ),
    .A3(_05299_),
    .B1(net18),
    .X(_05307_));
 sky130_fd_sc_hd__xor2_1 _26169_ (.A(\spi0.data_packed[7] ),
    .B(_05307_),
    .X(_05308_));
 sky130_fd_sc_hd__mux2_1 _26170_ (.A0(_05308_),
    .A1(\top0.cordic0.slte0.opB[9] ),
    .S(_12006_),
    .X(_05309_));
 sky130_fd_sc_hd__clkbuf_1 _26171_ (.A(_05309_),
    .X(_00820_));
 sky130_fd_sc_hd__and3_1 _26172_ (.A(\spi0.data_packed[6] ),
    .B(\spi0.data_packed[7] ),
    .C(_05303_),
    .X(_05310_));
 sky130_fd_sc_hd__nor2_1 _26173_ (.A(\spi0.data_packed[14] ),
    .B(_05310_),
    .Y(_05311_));
 sky130_fd_sc_hd__xnor2_1 _26174_ (.A(\spi0.data_packed[8] ),
    .B(_05311_),
    .Y(_05312_));
 sky130_fd_sc_hd__mux2_1 _26175_ (.A0(_05312_),
    .A1(\top0.cordic0.slte0.opB[10] ),
    .S(_12006_),
    .X(_05313_));
 sky130_fd_sc_hd__clkbuf_1 _26176_ (.A(_05313_),
    .X(_00821_));
 sky130_fd_sc_hd__and2_1 _26177_ (.A(\spi0.data_packed[8] ),
    .B(_05310_),
    .X(_05314_));
 sky130_fd_sc_hd__nor2_1 _26178_ (.A(net19),
    .B(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__xnor2_1 _26179_ (.A(\spi0.data_packed[9] ),
    .B(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__mux2_1 _26180_ (.A0(_05316_),
    .A1(\top0.cordic0.slte0.opB[11] ),
    .S(_12003_),
    .X(_05317_));
 sky130_fd_sc_hd__clkbuf_1 _26181_ (.A(_05317_),
    .X(_00822_));
 sky130_fd_sc_hd__a31o_1 _26182_ (.A1(\spi0.data_packed[8] ),
    .A2(\spi0.data_packed[9] ),
    .A3(_05310_),
    .B1(net18),
    .X(_05318_));
 sky130_fd_sc_hd__xor2_1 _26183_ (.A(\spi0.data_packed[10] ),
    .B(_05318_),
    .X(_05319_));
 sky130_fd_sc_hd__mux2_1 _26184_ (.A0(_05319_),
    .A1(\top0.cordic0.slte0.opB[12] ),
    .S(_12003_),
    .X(_05320_));
 sky130_fd_sc_hd__clkbuf_1 _26185_ (.A(_05320_),
    .X(_00823_));
 sky130_fd_sc_hd__and3_1 _26186_ (.A(\spi0.data_packed[9] ),
    .B(\spi0.data_packed[10] ),
    .C(_05314_),
    .X(_05321_));
 sky130_fd_sc_hd__nor2_1 _26187_ (.A(net18),
    .B(_05321_),
    .Y(_05322_));
 sky130_fd_sc_hd__xnor2_1 _26188_ (.A(\spi0.data_packed[11] ),
    .B(_05322_),
    .Y(_05323_));
 sky130_fd_sc_hd__mux2_1 _26189_ (.A0(_05323_),
    .A1(\top0.cordic0.slte0.opB[13] ),
    .S(_12003_),
    .X(_05324_));
 sky130_fd_sc_hd__clkbuf_1 _26190_ (.A(_05324_),
    .X(_00824_));
 sky130_fd_sc_hd__a21oi_1 _26191_ (.A1(\spi0.data_packed[11] ),
    .A2(_05321_),
    .B1(net18),
    .Y(_05325_));
 sky130_fd_sc_hd__xnor2_1 _26192_ (.A(\spi0.data_packed[12] ),
    .B(_05325_),
    .Y(_05326_));
 sky130_fd_sc_hd__mux2_1 _26193_ (.A0(_05326_),
    .A1(\top0.cordic0.slte0.opB[14] ),
    .S(_12003_),
    .X(_05327_));
 sky130_fd_sc_hd__clkbuf_1 _26194_ (.A(_05327_),
    .X(_00825_));
 sky130_fd_sc_hd__a31o_1 _26195_ (.A1(\spi0.data_packed[11] ),
    .A2(\spi0.data_packed[12] ),
    .A3(_05321_),
    .B1(net18),
    .X(_05328_));
 sky130_fd_sc_hd__xor2_1 _26196_ (.A(\spi0.data_packed[13] ),
    .B(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__mux2_1 _26197_ (.A0(_05329_),
    .A1(\top0.cordic0.slte0.opB[15] ),
    .S(_12003_),
    .X(_05330_));
 sky130_fd_sc_hd__clkbuf_1 _26198_ (.A(_05330_),
    .X(_00826_));
 sky130_fd_sc_hd__o21a_1 _26199_ (.A1(net209),
    .A2(\top0.svm0.out_valid ),
    .B1(net206),
    .X(_05331_));
 sky130_fd_sc_hd__o21a_1 _26200_ (.A1(net208),
    .A2(_12017_),
    .B1(\top0.ready ),
    .X(_05332_));
 sky130_fd_sc_hd__o22a_1 _26201_ (.A1(\top0.ready ),
    .A2(_05331_),
    .B1(_05332_),
    .B2(net207),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _26202_ (.A0(net3),
    .A1(\spi0.data_packed[0] ),
    .S(net694),
    .X(_05333_));
 sky130_fd_sc_hd__clkbuf_1 _26203_ (.A(_05333_),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _26204_ (.A0(\spi0.data_packed[0] ),
    .A1(\spi0.data_packed[1] ),
    .S(net694),
    .X(_05334_));
 sky130_fd_sc_hd__clkbuf_1 _26205_ (.A(_05334_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _26206_ (.A0(\spi0.data_packed[1] ),
    .A1(\spi0.data_packed[2] ),
    .S(net695),
    .X(_05335_));
 sky130_fd_sc_hd__clkbuf_1 _26207_ (.A(_05335_),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _26208_ (.A0(\spi0.data_packed[2] ),
    .A1(\spi0.data_packed[3] ),
    .S(net694),
    .X(_05336_));
 sky130_fd_sc_hd__clkbuf_1 _26209_ (.A(_05336_),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _26210_ (.A0(\spi0.data_packed[3] ),
    .A1(\spi0.data_packed[4] ),
    .S(net694),
    .X(_05337_));
 sky130_fd_sc_hd__clkbuf_1 _26211_ (.A(_05337_),
    .X(_00832_));
 sky130_fd_sc_hd__mux2_1 _26212_ (.A0(\spi0.data_packed[4] ),
    .A1(\spi0.data_packed[5] ),
    .S(net694),
    .X(_05338_));
 sky130_fd_sc_hd__clkbuf_1 _26213_ (.A(_05338_),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_1 _26214_ (.A0(\spi0.data_packed[5] ),
    .A1(\spi0.data_packed[6] ),
    .S(net694),
    .X(_05339_));
 sky130_fd_sc_hd__clkbuf_1 _26215_ (.A(_05339_),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _26216_ (.A0(\spi0.data_packed[6] ),
    .A1(\spi0.data_packed[7] ),
    .S(net694),
    .X(_05340_));
 sky130_fd_sc_hd__clkbuf_1 _26217_ (.A(_05340_),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _26218_ (.A0(\spi0.data_packed[7] ),
    .A1(\spi0.data_packed[8] ),
    .S(net694),
    .X(_05341_));
 sky130_fd_sc_hd__clkbuf_1 _26219_ (.A(_05341_),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _26220_ (.A0(\spi0.data_packed[8] ),
    .A1(\spi0.data_packed[9] ),
    .S(net694),
    .X(_05342_));
 sky130_fd_sc_hd__clkbuf_1 _26221_ (.A(_05342_),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _26222_ (.A0(\spi0.data_packed[9] ),
    .A1(\spi0.data_packed[10] ),
    .S(net695),
    .X(_05343_));
 sky130_fd_sc_hd__clkbuf_1 _26223_ (.A(_05343_),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _26224_ (.A0(\spi0.data_packed[10] ),
    .A1(\spi0.data_packed[11] ),
    .S(net695),
    .X(_05344_));
 sky130_fd_sc_hd__clkbuf_1 _26225_ (.A(_05344_),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _26226_ (.A0(\spi0.data_packed[11] ),
    .A1(\spi0.data_packed[12] ),
    .S(net695),
    .X(_05345_));
 sky130_fd_sc_hd__clkbuf_1 _26227_ (.A(_05345_),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _26228_ (.A0(\spi0.data_packed[12] ),
    .A1(\spi0.data_packed[13] ),
    .S(net695),
    .X(_05346_));
 sky130_fd_sc_hd__clkbuf_1 _26229_ (.A(_05346_),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _26230_ (.A0(\spi0.data_packed[13] ),
    .A1(net19),
    .S(net694),
    .X(_05347_));
 sky130_fd_sc_hd__clkbuf_1 _26231_ (.A(_05347_),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _26232_ (.A0(net19),
    .A1(\spi0.data_packed[15] ),
    .S(net695),
    .X(_05348_));
 sky130_fd_sc_hd__clkbuf_1 _26233_ (.A(_05348_),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _26234_ (.A0(\spi0.data_packed[15] ),
    .A1(\spi0.data_packed[16] ),
    .S(net695),
    .X(_05349_));
 sky130_fd_sc_hd__clkbuf_1 _26235_ (.A(_05349_),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _26236_ (.A0(\spi0.data_packed[16] ),
    .A1(\spi0.data_packed[17] ),
    .S(net697),
    .X(_05350_));
 sky130_fd_sc_hd__clkbuf_1 _26237_ (.A(_05350_),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _26238_ (.A0(\spi0.data_packed[17] ),
    .A1(\spi0.data_packed[18] ),
    .S(net697),
    .X(_05351_));
 sky130_fd_sc_hd__clkbuf_1 _26239_ (.A(_05351_),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _26240_ (.A0(\spi0.data_packed[18] ),
    .A1(\spi0.data_packed[19] ),
    .S(net697),
    .X(_05352_));
 sky130_fd_sc_hd__clkbuf_1 _26241_ (.A(_05352_),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _26242_ (.A0(\spi0.data_packed[19] ),
    .A1(\spi0.data_packed[20] ),
    .S(net697),
    .X(_05353_));
 sky130_fd_sc_hd__clkbuf_1 _26243_ (.A(_05353_),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _26244_ (.A0(\spi0.data_packed[20] ),
    .A1(\spi0.data_packed[21] ),
    .S(net698),
    .X(_05354_));
 sky130_fd_sc_hd__clkbuf_1 _26245_ (.A(_05354_),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _26246_ (.A0(\spi0.data_packed[21] ),
    .A1(\spi0.data_packed[22] ),
    .S(net698),
    .X(_05355_));
 sky130_fd_sc_hd__clkbuf_1 _26247_ (.A(_05355_),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _26248_ (.A0(\spi0.data_packed[22] ),
    .A1(\spi0.data_packed[23] ),
    .S(net698),
    .X(_05356_));
 sky130_fd_sc_hd__clkbuf_1 _26249_ (.A(_05356_),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _26250_ (.A0(\spi0.data_packed[23] ),
    .A1(\spi0.data_packed[24] ),
    .S(net698),
    .X(_05357_));
 sky130_fd_sc_hd__clkbuf_1 _26251_ (.A(_05357_),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _26252_ (.A0(\spi0.data_packed[24] ),
    .A1(\spi0.data_packed[25] ),
    .S(net698),
    .X(_05358_));
 sky130_fd_sc_hd__clkbuf_1 _26253_ (.A(_05358_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _26254_ (.A0(\spi0.data_packed[25] ),
    .A1(\spi0.data_packed[26] ),
    .S(net698),
    .X(_05359_));
 sky130_fd_sc_hd__clkbuf_1 _26255_ (.A(_05359_),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _26256_ (.A0(\spi0.data_packed[26] ),
    .A1(\spi0.data_packed[27] ),
    .S(net699),
    .X(_05360_));
 sky130_fd_sc_hd__clkbuf_1 _26257_ (.A(_05360_),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _26258_ (.A0(\spi0.data_packed[27] ),
    .A1(\spi0.data_packed[28] ),
    .S(net699),
    .X(_05361_));
 sky130_fd_sc_hd__clkbuf_1 _26259_ (.A(_05361_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _26260_ (.A0(\spi0.data_packed[28] ),
    .A1(\spi0.data_packed[29] ),
    .S(net699),
    .X(_05362_));
 sky130_fd_sc_hd__clkbuf_1 _26261_ (.A(_05362_),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _26262_ (.A0(\spi0.data_packed[29] ),
    .A1(\spi0.data_packed[30] ),
    .S(net696),
    .X(_05363_));
 sky130_fd_sc_hd__clkbuf_1 _26263_ (.A(_05363_),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _26264_ (.A0(\spi0.data_packed[30] ),
    .A1(\spi0.data_packed[31] ),
    .S(net696),
    .X(_05364_));
 sky130_fd_sc_hd__clkbuf_1 _26265_ (.A(_05364_),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _26266_ (.A0(\spi0.data_packed[31] ),
    .A1(\spi0.data_packed[32] ),
    .S(net690),
    .X(_05365_));
 sky130_fd_sc_hd__clkbuf_1 _26267_ (.A(_05365_),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _26268_ (.A0(\spi0.data_packed[32] ),
    .A1(\spi0.data_packed[33] ),
    .S(net688),
    .X(_05366_));
 sky130_fd_sc_hd__clkbuf_1 _26269_ (.A(_05366_),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _26270_ (.A0(net958),
    .A1(net944),
    .S(net688),
    .X(_05367_));
 sky130_fd_sc_hd__clkbuf_1 _26271_ (.A(_05367_),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_1 _26272_ (.A0(net944),
    .A1(\spi0.data_packed[35] ),
    .S(net688),
    .X(_05368_));
 sky130_fd_sc_hd__clkbuf_1 _26273_ (.A(net945),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _26274_ (.A0(net975),
    .A1(\spi0.data_packed[36] ),
    .S(net688),
    .X(_05369_));
 sky130_fd_sc_hd__clkbuf_1 _26275_ (.A(_05369_),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _26276_ (.A0(\spi0.data_packed[36] ),
    .A1(net973),
    .S(net688),
    .X(_05370_));
 sky130_fd_sc_hd__clkbuf_1 _26277_ (.A(net974),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _26278_ (.A0(net973),
    .A1(\spi0.data_packed[38] ),
    .S(net688),
    .X(_05371_));
 sky130_fd_sc_hd__clkbuf_1 _26279_ (.A(_05371_),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _26280_ (.A0(net953),
    .A1(\spi0.data_packed[39] ),
    .S(net688),
    .X(_05372_));
 sky130_fd_sc_hd__clkbuf_1 _26281_ (.A(net954),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _26282_ (.A0(net967),
    .A1(net946),
    .S(net688),
    .X(_05373_));
 sky130_fd_sc_hd__clkbuf_1 _26283_ (.A(_05373_),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _26284_ (.A0(net946),
    .A1(\spi0.data_packed[41] ),
    .S(net688),
    .X(_05374_));
 sky130_fd_sc_hd__clkbuf_1 _26285_ (.A(net947),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _26286_ (.A0(\spi0.data_packed[41] ),
    .A1(net956),
    .S(net688),
    .X(_05375_));
 sky130_fd_sc_hd__clkbuf_1 _26287_ (.A(net957),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _26288_ (.A0(\spi0.data_packed[42] ),
    .A1(net1011),
    .S(net689),
    .X(_05376_));
 sky130_fd_sc_hd__clkbuf_1 _26289_ (.A(_05376_),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _26290_ (.A0(net942),
    .A1(net925),
    .S(net690),
    .X(_05377_));
 sky130_fd_sc_hd__clkbuf_1 _26291_ (.A(_05377_),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _26292_ (.A0(net925),
    .A1(\spi0.data_packed[45] ),
    .S(net693),
    .X(_05378_));
 sky130_fd_sc_hd__clkbuf_1 _26293_ (.A(net926),
    .X(_00873_));
 sky130_fd_sc_hd__mux2_1 _26294_ (.A0(net949),
    .A1(\spi0.data_packed[46] ),
    .S(net693),
    .X(_05379_));
 sky130_fd_sc_hd__clkbuf_1 _26295_ (.A(net950),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _26296_ (.A0(net969),
    .A1(\spi0.data_packed[47] ),
    .S(net693),
    .X(_05380_));
 sky130_fd_sc_hd__clkbuf_1 _26297_ (.A(_05380_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _26298_ (.A0(\spi0.data_packed[47] ),
    .A1(\spi0.data_packed[48] ),
    .S(net697),
    .X(_05381_));
 sky130_fd_sc_hd__clkbuf_1 _26299_ (.A(_05381_),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _26300_ (.A0(\spi0.data_packed[48] ),
    .A1(\spi0.data_packed[49] ),
    .S(net697),
    .X(_05382_));
 sky130_fd_sc_hd__clkbuf_1 _26301_ (.A(_05382_),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _26302_ (.A0(\spi0.data_packed[49] ),
    .A1(\spi0.data_packed[50] ),
    .S(net697),
    .X(_05383_));
 sky130_fd_sc_hd__clkbuf_1 _26303_ (.A(_05383_),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _26304_ (.A0(\spi0.data_packed[50] ),
    .A1(\spi0.data_packed[51] ),
    .S(net697),
    .X(_05384_));
 sky130_fd_sc_hd__clkbuf_1 _26305_ (.A(_05384_),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _26306_ (.A0(\spi0.data_packed[51] ),
    .A1(\spi0.data_packed[52] ),
    .S(net697),
    .X(_05385_));
 sky130_fd_sc_hd__clkbuf_1 _26307_ (.A(_05385_),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _26308_ (.A0(\spi0.data_packed[52] ),
    .A1(\spi0.data_packed[53] ),
    .S(net697),
    .X(_05386_));
 sky130_fd_sc_hd__clkbuf_1 _26309_ (.A(_05386_),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _26310_ (.A0(\spi0.data_packed[53] ),
    .A1(\spi0.data_packed[54] ),
    .S(net700),
    .X(_05387_));
 sky130_fd_sc_hd__clkbuf_1 _26311_ (.A(_05387_),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_1 _26312_ (.A0(\spi0.data_packed[54] ),
    .A1(\spi0.data_packed[55] ),
    .S(net698),
    .X(_05388_));
 sky130_fd_sc_hd__clkbuf_1 _26313_ (.A(_05388_),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_1 _26314_ (.A0(\spi0.data_packed[55] ),
    .A1(\spi0.data_packed[56] ),
    .S(net698),
    .X(_05389_));
 sky130_fd_sc_hd__clkbuf_1 _26315_ (.A(_05389_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _26316_ (.A0(\spi0.data_packed[56] ),
    .A1(\spi0.data_packed[57] ),
    .S(net698),
    .X(_05390_));
 sky130_fd_sc_hd__clkbuf_1 _26317_ (.A(_05390_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _26318_ (.A0(\spi0.data_packed[57] ),
    .A1(\spi0.data_packed[58] ),
    .S(net699),
    .X(_05391_));
 sky130_fd_sc_hd__clkbuf_1 _26319_ (.A(_05391_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _26320_ (.A0(\spi0.data_packed[58] ),
    .A1(\spi0.data_packed[59] ),
    .S(net698),
    .X(_05392_));
 sky130_fd_sc_hd__clkbuf_1 _26321_ (.A(_05392_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _26322_ (.A0(\spi0.data_packed[59] ),
    .A1(\spi0.data_packed[60] ),
    .S(net699),
    .X(_05393_));
 sky130_fd_sc_hd__clkbuf_1 _26323_ (.A(_05393_),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _26324_ (.A0(\spi0.data_packed[60] ),
    .A1(\spi0.data_packed[61] ),
    .S(net699),
    .X(_05394_));
 sky130_fd_sc_hd__clkbuf_1 _26325_ (.A(_05394_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _26326_ (.A0(\spi0.data_packed[61] ),
    .A1(\spi0.data_packed[62] ),
    .S(net699),
    .X(_05395_));
 sky130_fd_sc_hd__clkbuf_1 _26327_ (.A(_05395_),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _26328_ (.A0(\spi0.data_packed[62] ),
    .A1(\spi0.data_packed[63] ),
    .S(net696),
    .X(_05396_));
 sky130_fd_sc_hd__clkbuf_1 _26329_ (.A(_05396_),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _26330_ (.A0(\spi0.data_packed[63] ),
    .A1(\spi0.data_packed[64] ),
    .S(net695),
    .X(_05397_));
 sky130_fd_sc_hd__clkbuf_1 _26331_ (.A(_05397_),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _26332_ (.A0(\spi0.data_packed[64] ),
    .A1(\spi0.data_packed[65] ),
    .S(net693),
    .X(_05398_));
 sky130_fd_sc_hd__clkbuf_1 _26333_ (.A(_05398_),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _26334_ (.A0(\spi0.data_packed[65] ),
    .A1(\spi0.data_packed[66] ),
    .S(net695),
    .X(_05399_));
 sky130_fd_sc_hd__clkbuf_1 _26335_ (.A(_05399_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _26336_ (.A0(\spi0.data_packed[66] ),
    .A1(\spi0.data_packed[67] ),
    .S(net690),
    .X(_05400_));
 sky130_fd_sc_hd__clkbuf_1 _26337_ (.A(_05400_),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_1 _26338_ (.A0(\spi0.data_packed[67] ),
    .A1(\spi0.data_packed[68] ),
    .S(net692),
    .X(_05401_));
 sky130_fd_sc_hd__clkbuf_1 _26339_ (.A(_05401_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _26340_ (.A0(\spi0.data_packed[68] ),
    .A1(\spi0.data_packed[69] ),
    .S(net692),
    .X(_05402_));
 sky130_fd_sc_hd__clkbuf_1 _26341_ (.A(_05402_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _26342_ (.A0(\spi0.data_packed[69] ),
    .A1(\spi0.data_packed[70] ),
    .S(net689),
    .X(_05403_));
 sky130_fd_sc_hd__clkbuf_1 _26343_ (.A(_05403_),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _26344_ (.A0(\spi0.data_packed[70] ),
    .A1(\spi0.data_packed[71] ),
    .S(net689),
    .X(_05404_));
 sky130_fd_sc_hd__clkbuf_1 _26345_ (.A(_05404_),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _26346_ (.A0(\spi0.data_packed[71] ),
    .A1(\spi0.data_packed[72] ),
    .S(net689),
    .X(_05405_));
 sky130_fd_sc_hd__clkbuf_1 _26347_ (.A(_05405_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _26348_ (.A0(\spi0.data_packed[72] ),
    .A1(\spi0.data_packed[73] ),
    .S(net692),
    .X(_05406_));
 sky130_fd_sc_hd__clkbuf_1 _26349_ (.A(_05406_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _26350_ (.A0(\spi0.data_packed[73] ),
    .A1(\spi0.data_packed[74] ),
    .S(net690),
    .X(_05407_));
 sky130_fd_sc_hd__clkbuf_1 _26351_ (.A(_05407_),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _26352_ (.A0(\spi0.data_packed[74] ),
    .A1(\spi0.data_packed[75] ),
    .S(net690),
    .X(_05408_));
 sky130_fd_sc_hd__clkbuf_1 _26353_ (.A(_05408_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _26354_ (.A0(\spi0.data_packed[75] ),
    .A1(\spi0.data_packed[76] ),
    .S(net690),
    .X(_05409_));
 sky130_fd_sc_hd__clkbuf_1 _26355_ (.A(_05409_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _26356_ (.A0(\spi0.data_packed[76] ),
    .A1(\spi0.data_packed[77] ),
    .S(net690),
    .X(_05410_));
 sky130_fd_sc_hd__clkbuf_1 _26357_ (.A(_05410_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _26358_ (.A0(\spi0.data_packed[77] ),
    .A1(\spi0.data_packed[78] ),
    .S(net690),
    .X(_05411_));
 sky130_fd_sc_hd__clkbuf_1 _26359_ (.A(_05411_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _26360_ (.A0(\spi0.data_packed[78] ),
    .A1(\spi0.data_packed[79] ),
    .S(net690),
    .X(_05412_));
 sky130_fd_sc_hd__clkbuf_1 _26361_ (.A(_05412_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _26362_ (.A0(\spi0.data_packed[79] ),
    .A1(\spi0.opcode[0] ),
    .S(net690),
    .X(_05413_));
 sky130_fd_sc_hd__clkbuf_1 _26363_ (.A(_05413_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _26364_ (.A0(\spi0.opcode[0] ),
    .A1(\spi0.opcode[1] ),
    .S(net691),
    .X(_05414_));
 sky130_fd_sc_hd__clkbuf_1 _26365_ (.A(_05414_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _26366_ (.A0(\spi0.opcode[1] ),
    .A1(\spi0.opcode[2] ),
    .S(net691),
    .X(_05415_));
 sky130_fd_sc_hd__clkbuf_1 _26367_ (.A(_05415_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _26368_ (.A0(\spi0.opcode[2] ),
    .A1(\spi0.opcode[3] ),
    .S(net691),
    .X(_05416_));
 sky130_fd_sc_hd__clkbuf_1 _26369_ (.A(_05416_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _26370_ (.A0(\spi0.opcode[3] ),
    .A1(\spi0.opcode[4] ),
    .S(net691),
    .X(_05417_));
 sky130_fd_sc_hd__clkbuf_1 _26371_ (.A(_05417_),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _26372_ (.A0(\spi0.opcode[4] ),
    .A1(\spi0.opcode[5] ),
    .S(net691),
    .X(_05418_));
 sky130_fd_sc_hd__clkbuf_1 _26373_ (.A(_05418_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _26374_ (.A0(\spi0.opcode[5] ),
    .A1(\spi0.opcode[6] ),
    .S(net696),
    .X(_05419_));
 sky130_fd_sc_hd__clkbuf_1 _26375_ (.A(_05419_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _26376_ (.A0(\spi0.opcode[6] ),
    .A1(net963),
    .S(net696),
    .X(_05420_));
 sky130_fd_sc_hd__clkbuf_1 _26377_ (.A(_05420_),
    .X(_00915_));
 sky130_fd_sc_hd__dfrtp_1 _26378_ (.CLK(clknet_leaf_40_clk_sys),
    .D(_00019_),
    .RESET_B(net682),
    .Q(\top0.svm0.tC[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26379_ (.CLK(clknet_leaf_43_clk_sys),
    .D(_00020_),
    .RESET_B(net682),
    .Q(\top0.svm0.tC[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26380_ (.CLK(clknet_leaf_42_clk_sys),
    .D(_00021_),
    .RESET_B(net684),
    .Q(\top0.svm0.tC[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26381_ (.CLK(clknet_leaf_42_clk_sys),
    .D(_00022_),
    .RESET_B(net684),
    .Q(\top0.svm0.tC[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26382_ (.CLK(clknet_leaf_42_clk_sys),
    .D(_00023_),
    .RESET_B(net684),
    .Q(\top0.svm0.tC[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26383_ (.CLK(clknet_leaf_42_clk_sys),
    .D(_00024_),
    .RESET_B(net684),
    .Q(\top0.svm0.tC[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26384_ (.CLK(clknet_leaf_41_clk_sys),
    .D(_00025_),
    .RESET_B(net684),
    .Q(\top0.svm0.tC[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26385_ (.CLK(clknet_leaf_41_clk_sys),
    .D(_00026_),
    .RESET_B(net685),
    .Q(\top0.svm0.tC[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26386_ (.CLK(clknet_leaf_41_clk_sys),
    .D(_00027_),
    .RESET_B(net682),
    .Q(\top0.svm0.tC[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26387_ (.CLK(clknet_leaf_39_clk_sys),
    .D(_00028_),
    .RESET_B(net682),
    .Q(\top0.svm0.tC[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26388_ (.CLK(clknet_leaf_38_clk_sys),
    .D(_00029_),
    .RESET_B(net677),
    .Q(\top0.svm0.tC[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26389_ (.CLK(clknet_leaf_39_clk_sys),
    .D(_00030_),
    .RESET_B(net677),
    .Q(\top0.svm0.tC[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26390_ (.CLK(clknet_leaf_39_clk_sys),
    .D(_00031_),
    .RESET_B(net677),
    .Q(\top0.svm0.tC[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26391_ (.CLK(clknet_leaf_38_clk_sys),
    .D(_00032_),
    .RESET_B(net677),
    .Q(\top0.svm0.tC[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26392_ (.CLK(clknet_leaf_37_clk_sys),
    .D(_00033_),
    .RESET_B(net679),
    .Q(\top0.svm0.tC[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26393_ (.CLK(clknet_leaf_37_clk_sys),
    .D(_00034_),
    .RESET_B(net679),
    .Q(\top0.svm0.tC[15] ));
 sky130_fd_sc_hd__dfstp_2 _26394_ (.CLK(clknet_leaf_86_clk_sys),
    .D(_00035_),
    .SET_B(net640),
    .Q(net7));
 sky130_fd_sc_hd__dfrtp_1 _26395_ (.CLK(clknet_leaf_85_clk_sys),
    .D(_00036_),
    .RESET_B(net640),
    .Q(\top0.kpd[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26396_ (.CLK(clknet_leaf_85_clk_sys),
    .D(_00037_),
    .RESET_B(net640),
    .Q(\top0.kpd[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26397_ (.CLK(clknet_leaf_79_clk_sys),
    .D(_00038_),
    .RESET_B(net632),
    .Q(\top0.kpd[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26398_ (.CLK(clknet_leaf_79_clk_sys),
    .D(_00039_),
    .RESET_B(net588),
    .Q(\top0.kpd[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26399_ (.CLK(clknet_leaf_98_clk_sys),
    .D(_00040_),
    .RESET_B(net588),
    .Q(\top0.kpd[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26400_ (.CLK(clknet_leaf_98_clk_sys),
    .D(_00041_),
    .RESET_B(net588),
    .Q(\top0.kpd[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26401_ (.CLK(clknet_leaf_98_clk_sys),
    .D(_00042_),
    .RESET_B(net588),
    .Q(\top0.kpd[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26402_ (.CLK(clknet_leaf_98_clk_sys),
    .D(_00043_),
    .RESET_B(net589),
    .Q(\top0.kpd[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26403_ (.CLK(clknet_leaf_98_clk_sys),
    .D(_00044_),
    .RESET_B(net588),
    .Q(\top0.kpd[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26404_ (.CLK(clknet_leaf_98_clk_sys),
    .D(_00045_),
    .RESET_B(net589),
    .Q(\top0.kpd[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26405_ (.CLK(clknet_leaf_79_clk_sys),
    .D(_00046_),
    .RESET_B(net632),
    .Q(\top0.kpd[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26406_ (.CLK(clknet_leaf_98_clk_sys),
    .D(_00047_),
    .RESET_B(net632),
    .Q(\top0.kpd[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26407_ (.CLK(clknet_leaf_79_clk_sys),
    .D(_00048_),
    .RESET_B(net632),
    .Q(\top0.kpd[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26408_ (.CLK(clknet_leaf_79_clk_sys),
    .D(_00049_),
    .RESET_B(net634),
    .Q(\top0.kpd[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26409_ (.CLK(clknet_leaf_85_clk_sys),
    .D(_00050_),
    .RESET_B(net634),
    .Q(\top0.kpd[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26410_ (.CLK(clknet_leaf_85_clk_sys),
    .D(_00051_),
    .RESET_B(net640),
    .Q(\top0.kpd[15] ));
 sky130_fd_sc_hd__dfrtp_1 _26411_ (.CLK(clknet_leaf_62_clk_sys),
    .D(_00052_),
    .RESET_B(net650),
    .Q(\top0.kpq[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26412_ (.CLK(clknet_leaf_62_clk_sys),
    .D(_00053_),
    .RESET_B(net646),
    .Q(\top0.kpq[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26413_ (.CLK(clknet_leaf_61_clk_sys),
    .D(_00054_),
    .RESET_B(net650),
    .Q(\top0.kpq[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26414_ (.CLK(clknet_leaf_62_clk_sys),
    .D(_00055_),
    .RESET_B(net650),
    .Q(\top0.kpq[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26415_ (.CLK(clknet_leaf_61_clk_sys),
    .D(_00056_),
    .RESET_B(net650),
    .Q(\top0.kpq[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26416_ (.CLK(clknet_leaf_61_clk_sys),
    .D(_00057_),
    .RESET_B(net650),
    .Q(\top0.kpq[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26417_ (.CLK(clknet_leaf_59_clk_sys),
    .D(_00058_),
    .RESET_B(net650),
    .Q(\top0.kpq[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26418_ (.CLK(clknet_leaf_60_clk_sys),
    .D(_00059_),
    .RESET_B(net650),
    .Q(\top0.kpq[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26419_ (.CLK(clknet_leaf_60_clk_sys),
    .D(_00060_),
    .RESET_B(net650),
    .Q(\top0.kpq[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26420_ (.CLK(clknet_leaf_58_clk_sys),
    .D(_00061_),
    .RESET_B(net650),
    .Q(\top0.kpq[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26421_ (.CLK(clknet_leaf_60_clk_sys),
    .D(_00062_),
    .RESET_B(net650),
    .Q(\top0.kpq[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26422_ (.CLK(clknet_leaf_58_clk_sys),
    .D(_00063_),
    .RESET_B(net653),
    .Q(\top0.kpq[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26423_ (.CLK(clknet_leaf_58_clk_sys),
    .D(_00064_),
    .RESET_B(net644),
    .Q(\top0.kpq[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26424_ (.CLK(clknet_leaf_56_clk_sys),
    .D(_00065_),
    .RESET_B(net664),
    .Q(\top0.kpq[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26425_ (.CLK(clknet_leaf_57_clk_sys),
    .D(_00066_),
    .RESET_B(net644),
    .Q(\top0.kpq[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26426_ (.CLK(clknet_leaf_88_clk_sys),
    .D(_00067_),
    .RESET_B(net642),
    .Q(\top0.kpq[15] ));
 sky130_fd_sc_hd__dfrtp_1 _26427_ (.CLK(clknet_leaf_78_clk_sys),
    .D(_00068_),
    .RESET_B(net632),
    .Q(\top0.kid[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26428_ (.CLK(clknet_leaf_77_clk_sys),
    .D(_00069_),
    .RESET_B(net631),
    .Q(\top0.kid[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26429_ (.CLK(clknet_leaf_77_clk_sys),
    .D(_00070_),
    .RESET_B(net631),
    .Q(\top0.kid[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26430_ (.CLK(clknet_leaf_77_clk_sys),
    .D(_00071_),
    .RESET_B(net631),
    .Q(\top0.kid[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26431_ (.CLK(clknet_leaf_99_clk_sys),
    .D(_00072_),
    .RESET_B(net631),
    .Q(\top0.kid[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26432_ (.CLK(clknet_leaf_77_clk_sys),
    .D(_00073_),
    .RESET_B(net631),
    .Q(\top0.kid[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26433_ (.CLK(clknet_leaf_99_clk_sys),
    .D(_00074_),
    .RESET_B(net631),
    .Q(\top0.kid[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26434_ (.CLK(clknet_leaf_98_clk_sys),
    .D(_00075_),
    .RESET_B(net589),
    .Q(\top0.kid[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26435_ (.CLK(clknet_leaf_79_clk_sys),
    .D(_00076_),
    .RESET_B(net632),
    .Q(\top0.kid[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26436_ (.CLK(clknet_leaf_79_clk_sys),
    .D(_00077_),
    .RESET_B(net632),
    .Q(\top0.kid[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26437_ (.CLK(clknet_leaf_79_clk_sys),
    .D(_00078_),
    .RESET_B(net632),
    .Q(\top0.kid[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26438_ (.CLK(clknet_leaf_79_clk_sys),
    .D(_00079_),
    .RESET_B(net634),
    .Q(\top0.kid[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26439_ (.CLK(clknet_leaf_80_clk_sys),
    .D(_00080_),
    .RESET_B(net634),
    .Q(\top0.kid[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26440_ (.CLK(clknet_leaf_80_clk_sys),
    .D(_00081_),
    .RESET_B(net633),
    .Q(\top0.kid[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26441_ (.CLK(clknet_leaf_80_clk_sys),
    .D(_00082_),
    .RESET_B(net640),
    .Q(\top0.kid[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26442_ (.CLK(clknet_leaf_84_clk_sys),
    .D(_00083_),
    .RESET_B(net640),
    .Q(\top0.kid[15] ));
 sky130_fd_sc_hd__dfrtp_1 _26443_ (.CLK(clknet_leaf_87_clk_sys),
    .D(_00084_),
    .RESET_B(net644),
    .Q(\top0.kiq[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26444_ (.CLK(clknet_leaf_87_clk_sys),
    .D(_00085_),
    .RESET_B(net644),
    .Q(\top0.kiq[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26445_ (.CLK(clknet_leaf_87_clk_sys),
    .D(_00086_),
    .RESET_B(net644),
    .Q(\top0.kiq[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26446_ (.CLK(clknet_leaf_59_clk_sys),
    .D(_00087_),
    .RESET_B(net644),
    .Q(\top0.kiq[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26447_ (.CLK(clknet_leaf_59_clk_sys),
    .D(_00088_),
    .RESET_B(net644),
    .Q(\top0.kiq[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26448_ (.CLK(clknet_leaf_60_clk_sys),
    .D(_00089_),
    .RESET_B(net651),
    .Q(\top0.kiq[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26449_ (.CLK(clknet_leaf_55_clk_sys),
    .D(_00090_),
    .RESET_B(net667),
    .Q(\top0.kiq[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26450_ (.CLK(clknet_leaf_55_clk_sys),
    .D(_00091_),
    .RESET_B(net667),
    .Q(\top0.kiq[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26451_ (.CLK(clknet_leaf_55_clk_sys),
    .D(_00092_),
    .RESET_B(net668),
    .Q(\top0.kiq[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26452_ (.CLK(clknet_leaf_55_clk_sys),
    .D(_00093_),
    .RESET_B(net668),
    .Q(\top0.kiq[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26453_ (.CLK(clknet_leaf_55_clk_sys),
    .D(_00094_),
    .RESET_B(net668),
    .Q(\top0.kiq[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26454_ (.CLK(clknet_leaf_55_clk_sys),
    .D(_00095_),
    .RESET_B(net668),
    .Q(\top0.kiq[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26455_ (.CLK(clknet_leaf_57_clk_sys),
    .D(_00096_),
    .RESET_B(net642),
    .Q(\top0.kiq[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26456_ (.CLK(clknet_leaf_57_clk_sys),
    .D(_00097_),
    .RESET_B(net664),
    .Q(\top0.kiq[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26457_ (.CLK(clknet_leaf_57_clk_sys),
    .D(_00098_),
    .RESET_B(net642),
    .Q(\top0.kiq[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26458_ (.CLK(clknet_leaf_88_clk_sys),
    .D(_00099_),
    .RESET_B(net642),
    .Q(\top0.kiq[15] ));
 sky130_fd_sc_hd__dfstp_1 _26459_ (.CLK(clknet_leaf_91_clk_sys),
    .D(net692),
    .SET_B(net600),
    .Q(\spi0.cs_sync[0] ));
 sky130_fd_sc_hd__dfstp_1 _26460_ (.CLK(clknet_leaf_91_clk_sys),
    .D(net701),
    .SET_B(net600),
    .Q(\spi0.cs_sync[1] ));
 sky130_fd_sc_hd__dfstp_1 _26461_ (.CLK(clknet_leaf_91_clk_sys),
    .D(net702),
    .SET_B(net640),
    .Q(\spi0.cs_sync[2] ));
 sky130_fd_sc_hd__dfstp_1 _26462_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00014_),
    .SET_B(net601),
    .Q(\top0.matmul0.matmul_stage_inst.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26463_ (.CLK(clknet_leaf_16_clk_sys),
    .D(net560),
    .RESET_B(net611),
    .Q(\top0.matmul0.matmul_stage_inst.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26464_ (.CLK(clknet_leaf_17_clk_sys),
    .D(net567),
    .RESET_B(net612),
    .Q(\top0.matmul0.matmul_stage_inst.state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _26465_ (.CLK(clknet_leaf_14_clk_sys),
    .D(net563),
    .RESET_B(net617),
    .Q(\top0.matmul0.done_pass ));
 sky130_fd_sc_hd__dfrtp_2 _26466_ (.CLK(clknet_leaf_17_clk_sys),
    .D(_00000_),
    .RESET_B(net611),
    .Q(\top0.matmul0.matmul_stage_inst.state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26467_ (.CLK(clknet_leaf_18_clk_sys),
    .D(net575),
    .RESET_B(net612),
    .Q(\top0.matmul0.matmul_stage_inst.state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26468_ (.CLK(clknet_leaf_16_clk_sys),
    .D(net570),
    .RESET_B(net611),
    .Q(\top0.matmul0.matmul_stage_inst.state[6] ));
 sky130_fd_sc_hd__dfstp_1 _26469_ (.CLK(clknet_leaf_45_clk_sys),
    .D(_00100_),
    .SET_B(net681),
    .Q(\top0.svm0.delta[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26470_ (.CLK(clknet_leaf_12_clk_sys),
    .D(_00101_),
    .RESET_B(net618),
    .Q(\top0.periodTop[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26471_ (.CLK(clknet_leaf_12_clk_sys),
    .D(_00102_),
    .RESET_B(net603),
    .Q(\top0.periodTop[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26472_ (.CLK(clknet_leaf_12_clk_sys),
    .D(_00103_),
    .RESET_B(net603),
    .Q(\top0.periodTop[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26473_ (.CLK(clknet_leaf_12_clk_sys),
    .D(_00104_),
    .RESET_B(net603),
    .Q(\top0.periodTop[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26474_ (.CLK(clknet_leaf_12_clk_sys),
    .D(_00105_),
    .RESET_B(net604),
    .Q(\top0.periodTop[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26475_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00106_),
    .RESET_B(net604),
    .Q(\top0.periodTop[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26476_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00107_),
    .RESET_B(net603),
    .Q(\top0.periodTop[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26477_ (.CLK(clknet_leaf_89_clk_sys),
    .D(_00108_),
    .RESET_B(net603),
    .Q(\top0.periodTop[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26478_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00109_),
    .RESET_B(net604),
    .Q(\top0.periodTop[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26479_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00110_),
    .RESET_B(net604),
    .Q(\top0.periodTop[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26480_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00111_),
    .RESET_B(net601),
    .Q(\top0.periodTop[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26481_ (.CLK(clknet_leaf_89_clk_sys),
    .D(_00112_),
    .RESET_B(net603),
    .Q(\top0.periodTop[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26482_ (.CLK(clknet_leaf_89_clk_sys),
    .D(_00113_),
    .RESET_B(net604),
    .Q(\top0.periodTop[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26483_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00114_),
    .RESET_B(net604),
    .Q(\top0.periodTop[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26484_ (.CLK(clknet_leaf_89_clk_sys),
    .D(_00115_),
    .RESET_B(net604),
    .Q(\top0.periodTop[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26485_ (.CLK(clknet_leaf_89_clk_sys),
    .D(_00116_),
    .RESET_B(net603),
    .Q(\top0.periodTop[15] ));
 sky130_fd_sc_hd__dfstp_1 _26486_ (.CLK(clknet_leaf_62_clk_sys),
    .D(_00018_),
    .SET_B(net647),
    .Q(\top0.pid_q.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26487_ (.CLK(clknet_leaf_66_clk_sys),
    .D(_00007_),
    .RESET_B(net660),
    .Q(\top0.pid_q.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26488_ (.CLK(clknet_leaf_55_clk_sys),
    .D(_00008_),
    .RESET_B(net667),
    .Q(\top0.pid_q.state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _26489_ (.CLK(clknet_leaf_61_clk_sys),
    .D(_00009_),
    .RESET_B(net651),
    .Q(\top0.pid_q.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26490_ (.CLK(clknet_leaf_63_clk_sys),
    .D(_00010_),
    .RESET_B(net656),
    .Q(\top0.pid_q.state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26491_ (.CLK(clknet_leaf_67_clk_sys),
    .D(_00011_),
    .RESET_B(net659),
    .Q(\top0.pid_q.state[5] ));
 sky130_fd_sc_hd__dfstp_2 _26492_ (.CLK(clknet_leaf_85_clk_sys),
    .D(_00012_),
    .SET_B(net640),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26493_ (.CLK(clknet_leaf_86_clk_sys),
    .D(_00013_),
    .RESET_B(net640),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _26494_ (.CLK(clknet_leaf_71_clk_sys),
    .D(_00117_),
    .RESET_B(net657),
    .Q(\top0.pid_d.prev_int[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26495_ (.CLK(clknet_leaf_71_clk_sys),
    .D(_00118_),
    .RESET_B(net657),
    .Q(\top0.pid_d.prev_int[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26496_ (.CLK(clknet_leaf_73_clk_sys),
    .D(_00119_),
    .RESET_B(net655),
    .Q(\top0.pid_d.prev_int[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26497_ (.CLK(clknet_leaf_72_clk_sys),
    .D(_00120_),
    .RESET_B(net655),
    .Q(\top0.pid_d.prev_int[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26498_ (.CLK(clknet_leaf_73_clk_sys),
    .D(_00121_),
    .RESET_B(net655),
    .Q(\top0.pid_d.prev_int[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26499_ (.CLK(clknet_leaf_74_clk_sys),
    .D(_00122_),
    .RESET_B(net655),
    .Q(\top0.pid_d.prev_int[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26500_ (.CLK(clknet_leaf_74_clk_sys),
    .D(_00123_),
    .RESET_B(net637),
    .Q(\top0.pid_d.prev_int[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26501_ (.CLK(clknet_leaf_82_clk_sys),
    .D(net912),
    .RESET_B(net636),
    .Q(\top0.pid_d.prev_int[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26502_ (.CLK(clknet_leaf_81_clk_sys),
    .D(_00125_),
    .RESET_B(net636),
    .Q(\top0.pid_d.prev_int[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26503_ (.CLK(clknet_leaf_82_clk_sys),
    .D(_00126_),
    .RESET_B(net637),
    .Q(\top0.pid_d.prev_int[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26504_ (.CLK(clknet_leaf_84_clk_sys),
    .D(net829),
    .RESET_B(net633),
    .Q(\top0.pid_d.prev_int[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26505_ (.CLK(clknet_leaf_81_clk_sys),
    .D(_00128_),
    .RESET_B(net638),
    .Q(\top0.pid_d.prev_int[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26506_ (.CLK(clknet_leaf_78_clk_sys),
    .D(_00129_),
    .RESET_B(net639),
    .Q(\top0.pid_d.prev_int[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26507_ (.CLK(clknet_leaf_77_clk_sys),
    .D(_00130_),
    .RESET_B(net631),
    .Q(\top0.pid_d.prev_int[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26508_ (.CLK(clknet_leaf_77_clk_sys),
    .D(_00131_),
    .RESET_B(net631),
    .Q(\top0.pid_d.prev_int[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26509_ (.CLK(clknet_leaf_77_clk_sys),
    .D(net816),
    .RESET_B(net631),
    .Q(\top0.pid_d.prev_int[15] ));
 sky130_fd_sc_hd__dfrtp_4 _26510_ (.CLK(clknet_leaf_66_clk_sys),
    .D(_00133_),
    .RESET_B(net660),
    .Q(\top0.pid_q.out[0] ));
 sky130_fd_sc_hd__dfrtp_4 _26511_ (.CLK(clknet_leaf_64_clk_sys),
    .D(_00134_),
    .RESET_B(net656),
    .Q(\top0.pid_q.out[1] ));
 sky130_fd_sc_hd__dfrtp_4 _26512_ (.CLK(clknet_leaf_66_clk_sys),
    .D(_00135_),
    .RESET_B(net659),
    .Q(\top0.pid_q.out[2] ));
 sky130_fd_sc_hd__dfrtp_4 _26513_ (.CLK(clknet_leaf_65_clk_sys),
    .D(_00136_),
    .RESET_B(net657),
    .Q(\top0.pid_q.out[3] ));
 sky130_fd_sc_hd__dfrtp_4 _26514_ (.CLK(clknet_leaf_65_clk_sys),
    .D(_00137_),
    .RESET_B(net659),
    .Q(\top0.pid_q.out[4] ));
 sky130_fd_sc_hd__dfrtp_4 _26515_ (.CLK(clknet_leaf_66_clk_sys),
    .D(_00138_),
    .RESET_B(net659),
    .Q(\top0.pid_q.out[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26516_ (.CLK(clknet_leaf_66_clk_sys),
    .D(_00139_),
    .RESET_B(net659),
    .Q(\top0.pid_q.out[6] ));
 sky130_fd_sc_hd__dfrtp_2 _26517_ (.CLK(clknet_leaf_68_clk_sys),
    .D(_00140_),
    .RESET_B(net659),
    .Q(\top0.pid_q.out[7] ));
 sky130_fd_sc_hd__dfrtp_4 _26518_ (.CLK(clknet_leaf_67_clk_sys),
    .D(_00141_),
    .RESET_B(net659),
    .Q(\top0.pid_q.out[8] ));
 sky130_fd_sc_hd__dfrtp_4 _26519_ (.CLK(clknet_leaf_66_clk_sys),
    .D(_00142_),
    .RESET_B(net659),
    .Q(\top0.pid_q.out[9] ));
 sky130_fd_sc_hd__dfrtp_2 _26520_ (.CLK(clknet_leaf_66_clk_sys),
    .D(_00143_),
    .RESET_B(net660),
    .Q(\top0.pid_q.out[10] ));
 sky130_fd_sc_hd__dfrtp_4 _26521_ (.CLK(clknet_leaf_66_clk_sys),
    .D(_00144_),
    .RESET_B(net660),
    .Q(\top0.pid_q.out[11] ));
 sky130_fd_sc_hd__dfrtp_4 _26522_ (.CLK(clknet_leaf_66_clk_sys),
    .D(_00145_),
    .RESET_B(net660),
    .Q(\top0.pid_q.out[12] ));
 sky130_fd_sc_hd__dfrtp_4 _26523_ (.CLK(clknet_leaf_61_clk_sys),
    .D(_00146_),
    .RESET_B(net651),
    .Q(\top0.pid_q.out[13] ));
 sky130_fd_sc_hd__dfrtp_4 _26524_ (.CLK(clknet_leaf_66_clk_sys),
    .D(_00147_),
    .RESET_B(net660),
    .Q(\top0.pid_q.out[14] ));
 sky130_fd_sc_hd__dfrtp_2 _26525_ (.CLK(clknet_leaf_60_clk_sys),
    .D(_00148_),
    .RESET_B(net651),
    .Q(\top0.pid_q.out[15] ));
 sky130_fd_sc_hd__dfrtp_1 _26526_ (.CLK(clknet_leaf_63_clk_sys),
    .D(_00149_),
    .RESET_B(net647),
    .Q(\top0.pid_q.mult0.a[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26527_ (.CLK(clknet_leaf_61_clk_sys),
    .D(_00150_),
    .RESET_B(net647),
    .Q(\top0.pid_q.mult0.a[1] ));
 sky130_fd_sc_hd__dfrtp_4 _26528_ (.CLK(clknet_leaf_61_clk_sys),
    .D(_00151_),
    .RESET_B(net651),
    .Q(\top0.pid_q.mult0.a[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26529_ (.CLK(clknet_leaf_61_clk_sys),
    .D(_00152_),
    .RESET_B(net651),
    .Q(\top0.pid_q.mult0.a[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26530_ (.CLK(clknet_leaf_61_clk_sys),
    .D(_00153_),
    .RESET_B(net651),
    .Q(\top0.pid_q.mult0.a[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26531_ (.CLK(clknet_leaf_61_clk_sys),
    .D(_00154_),
    .RESET_B(net651),
    .Q(\top0.pid_q.mult0.a[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26532_ (.CLK(clknet_leaf_61_clk_sys),
    .D(_00155_),
    .RESET_B(net651),
    .Q(\top0.pid_q.mult0.a[6] ));
 sky130_fd_sc_hd__dfrtp_2 _26533_ (.CLK(clknet_leaf_61_clk_sys),
    .D(_00156_),
    .RESET_B(net651),
    .Q(\top0.pid_q.mult0.a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26534_ (.CLK(clknet_leaf_61_clk_sys),
    .D(_00157_),
    .RESET_B(net652),
    .Q(\top0.pid_q.mult0.a[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26535_ (.CLK(clknet_leaf_60_clk_sys),
    .D(_00158_),
    .RESET_B(net652),
    .Q(\top0.pid_q.mult0.a[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26536_ (.CLK(clknet_leaf_60_clk_sys),
    .D(_00159_),
    .RESET_B(net652),
    .Q(\top0.pid_q.mult0.a[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26537_ (.CLK(clknet_leaf_60_clk_sys),
    .D(_00160_),
    .RESET_B(net652),
    .Q(\top0.pid_q.mult0.a[11] ));
 sky130_fd_sc_hd__dfrtp_4 _26538_ (.CLK(clknet_leaf_60_clk_sys),
    .D(_00161_),
    .RESET_B(net653),
    .Q(\top0.pid_q.mult0.a[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26539_ (.CLK(clknet_leaf_60_clk_sys),
    .D(_00162_),
    .RESET_B(net668),
    .Q(\top0.pid_q.mult0.a[13] ));
 sky130_fd_sc_hd__dfrtp_2 _26540_ (.CLK(clknet_leaf_60_clk_sys),
    .D(_00163_),
    .RESET_B(net653),
    .Q(\top0.pid_q.mult0.a[14] ));
 sky130_fd_sc_hd__dfrtp_2 _26541_ (.CLK(clknet_leaf_60_clk_sys),
    .D(_00164_),
    .RESET_B(net653),
    .Q(\top0.pid_q.mult0.a[15] ));
 sky130_fd_sc_hd__dfrtp_1 _26542_ (.CLK(clknet_leaf_51_clk_sys),
    .D(_00165_),
    .RESET_B(net671),
    .Q(\top0.pid_q.mult0.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26543_ (.CLK(clknet_leaf_69_clk_sys),
    .D(_00166_),
    .RESET_B(net662),
    .Q(\top0.pid_q.mult0.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26544_ (.CLK(clknet_leaf_51_clk_sys),
    .D(_00167_),
    .RESET_B(net661),
    .Q(\top0.pid_q.mult0.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26545_ (.CLK(clknet_leaf_49_clk_sys),
    .D(_00168_),
    .RESET_B(net675),
    .Q(\top0.pid_q.mult0.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26546_ (.CLK(clknet_leaf_49_clk_sys),
    .D(_00169_),
    .RESET_B(net675),
    .Q(\top0.pid_q.mult0.b[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26547_ (.CLK(clknet_leaf_49_clk_sys),
    .D(_00170_),
    .RESET_B(net675),
    .Q(\top0.pid_q.mult0.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26548_ (.CLK(clknet_leaf_49_clk_sys),
    .D(_00171_),
    .RESET_B(net675),
    .Q(\top0.pid_q.mult0.b[6] ));
 sky130_fd_sc_hd__dfrtp_2 _26549_ (.CLK(clknet_leaf_50_clk_sys),
    .D(_00172_),
    .RESET_B(net675),
    .Q(\top0.pid_q.mult0.b[7] ));
 sky130_fd_sc_hd__dfrtp_2 _26550_ (.CLK(clknet_leaf_50_clk_sys),
    .D(_00173_),
    .RESET_B(net675),
    .Q(\top0.pid_q.mult0.b[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26551_ (.CLK(clknet_leaf_52_clk_sys),
    .D(_00174_),
    .RESET_B(net671),
    .Q(\top0.pid_q.mult0.b[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26552_ (.CLK(clknet_leaf_51_clk_sys),
    .D(_00175_),
    .RESET_B(net671),
    .Q(\top0.pid_q.mult0.b[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26553_ (.CLK(clknet_leaf_49_clk_sys),
    .D(_00176_),
    .RESET_B(net675),
    .Q(\top0.pid_q.mult0.b[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26554_ (.CLK(clknet_leaf_52_clk_sys),
    .D(_00177_),
    .RESET_B(net670),
    .Q(\top0.pid_q.mult0.b[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26555_ (.CLK(clknet_leaf_49_clk_sys),
    .D(_00178_),
    .RESET_B(net675),
    .Q(\top0.pid_q.mult0.b[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26556_ (.CLK(clknet_leaf_49_clk_sys),
    .D(_00179_),
    .RESET_B(net675),
    .Q(\top0.pid_q.mult0.b[14] ));
 sky130_fd_sc_hd__dfrtp_4 _26557_ (.CLK(clknet_leaf_49_clk_sys),
    .D(_00180_),
    .RESET_B(net687),
    .Q(\top0.pid_q.mult0.b[15] ));
 sky130_fd_sc_hd__dfrtp_2 _26558_ (.CLK(clknet_leaf_52_clk_sys),
    .D(_00181_),
    .RESET_B(net670),
    .Q(\top0.pid_q.curr_error[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26559_ (.CLK(clknet_leaf_51_clk_sys),
    .D(_00182_),
    .RESET_B(net670),
    .Q(\top0.pid_q.curr_error[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26560_ (.CLK(clknet_leaf_52_clk_sys),
    .D(_00183_),
    .RESET_B(net670),
    .Q(\top0.pid_q.curr_error[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26561_ (.CLK(clknet_leaf_51_clk_sys),
    .D(_00184_),
    .RESET_B(net671),
    .Q(\top0.pid_q.curr_error[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26562_ (.CLK(clknet_leaf_51_clk_sys),
    .D(_00185_),
    .RESET_B(net671),
    .Q(\top0.pid_q.curr_error[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26563_ (.CLK(clknet_leaf_50_clk_sys),
    .D(_00186_),
    .RESET_B(net671),
    .Q(\top0.pid_q.curr_error[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26564_ (.CLK(clknet_leaf_53_clk_sys),
    .D(_00187_),
    .RESET_B(net671),
    .Q(\top0.pid_q.curr_error[6] ));
 sky130_fd_sc_hd__dfrtp_2 _26565_ (.CLK(clknet_leaf_53_clk_sys),
    .D(_00188_),
    .RESET_B(net672),
    .Q(\top0.pid_q.curr_error[7] ));
 sky130_fd_sc_hd__dfrtp_2 _26566_ (.CLK(clknet_leaf_53_clk_sys),
    .D(_00189_),
    .RESET_B(net672),
    .Q(\top0.pid_q.curr_error[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26567_ (.CLK(clknet_leaf_52_clk_sys),
    .D(_00190_),
    .RESET_B(net672),
    .Q(\top0.pid_q.curr_error[9] ));
 sky130_fd_sc_hd__dfrtp_2 _26568_ (.CLK(clknet_leaf_52_clk_sys),
    .D(_00191_),
    .RESET_B(net673),
    .Q(\top0.pid_q.curr_error[10] ));
 sky130_fd_sc_hd__dfrtp_2 _26569_ (.CLK(clknet_leaf_54_clk_sys),
    .D(_00192_),
    .RESET_B(net667),
    .Q(\top0.pid_q.curr_error[11] ));
 sky130_fd_sc_hd__dfrtp_2 _26570_ (.CLK(clknet_leaf_52_clk_sys),
    .D(_00193_),
    .RESET_B(net673),
    .Q(\top0.pid_q.curr_error[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26571_ (.CLK(clknet_leaf_54_clk_sys),
    .D(_00194_),
    .RESET_B(net667),
    .Q(\top0.pid_q.curr_error[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26572_ (.CLK(clknet_leaf_54_clk_sys),
    .D(_00195_),
    .RESET_B(net667),
    .Q(\top0.pid_q.curr_error[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26573_ (.CLK(clknet_leaf_55_clk_sys),
    .D(_00196_),
    .RESET_B(net667),
    .Q(\top0.pid_q.curr_error[15] ));
 sky130_fd_sc_hd__dfrtp_2 _26574_ (.CLK(clknet_leaf_52_clk_sys),
    .D(_00197_),
    .RESET_B(net670),
    .Q(\top0.pid_q.prev_error[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26575_ (.CLK(clknet_leaf_52_clk_sys),
    .D(_00198_),
    .RESET_B(net671),
    .Q(\top0.pid_q.prev_error[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26576_ (.CLK(clknet_leaf_52_clk_sys),
    .D(_00199_),
    .RESET_B(net672),
    .Q(\top0.pid_q.prev_error[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26577_ (.CLK(clknet_leaf_50_clk_sys),
    .D(_00200_),
    .RESET_B(net671),
    .Q(\top0.pid_q.prev_error[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26578_ (.CLK(clknet_leaf_50_clk_sys),
    .D(_00201_),
    .RESET_B(net671),
    .Q(\top0.pid_q.prev_error[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26579_ (.CLK(clknet_leaf_50_clk_sys),
    .D(_00202_),
    .RESET_B(net672),
    .Q(\top0.pid_q.prev_error[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26580_ (.CLK(clknet_leaf_53_clk_sys),
    .D(_00203_),
    .RESET_B(net672),
    .Q(\top0.pid_q.prev_error[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26581_ (.CLK(clknet_leaf_53_clk_sys),
    .D(_00204_),
    .RESET_B(net674),
    .Q(\top0.pid_q.prev_error[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26582_ (.CLK(clknet_leaf_53_clk_sys),
    .D(_00205_),
    .RESET_B(net674),
    .Q(\top0.pid_q.prev_error[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26583_ (.CLK(clknet_leaf_53_clk_sys),
    .D(_00206_),
    .RESET_B(net674),
    .Q(\top0.pid_q.prev_error[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26584_ (.CLK(clknet_leaf_53_clk_sys),
    .D(_00207_),
    .RESET_B(net674),
    .Q(\top0.pid_q.prev_error[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26585_ (.CLK(clknet_leaf_54_clk_sys),
    .D(_00208_),
    .RESET_B(net673),
    .Q(\top0.pid_q.prev_error[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26586_ (.CLK(clknet_leaf_54_clk_sys),
    .D(_00209_),
    .RESET_B(net667),
    .Q(\top0.pid_q.prev_error[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26587_ (.CLK(clknet_leaf_54_clk_sys),
    .D(_00210_),
    .RESET_B(net667),
    .Q(\top0.pid_q.prev_error[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26588_ (.CLK(clknet_leaf_54_clk_sys),
    .D(_00211_),
    .RESET_B(net669),
    .Q(\top0.pid_q.prev_error[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26589_ (.CLK(clknet_leaf_54_clk_sys),
    .D(_00212_),
    .RESET_B(net669),
    .Q(\top0.pid_q.prev_error[15] ));
 sky130_fd_sc_hd__dfrtp_4 _26590_ (.CLK(clknet_leaf_65_clk_sys),
    .D(_00213_),
    .RESET_B(net660),
    .Q(\top0.pid_q.curr_int[0] ));
 sky130_fd_sc_hd__dfrtp_4 _26591_ (.CLK(clknet_leaf_65_clk_sys),
    .D(_00214_),
    .RESET_B(net657),
    .Q(\top0.pid_q.curr_int[1] ));
 sky130_fd_sc_hd__dfrtp_4 _26592_ (.CLK(clknet_leaf_65_clk_sys),
    .D(_00215_),
    .RESET_B(net657),
    .Q(\top0.pid_q.curr_int[2] ));
 sky130_fd_sc_hd__dfrtp_4 _26593_ (.CLK(clknet_leaf_70_clk_sys),
    .D(_00216_),
    .RESET_B(net662),
    .Q(\top0.pid_q.curr_int[3] ));
 sky130_fd_sc_hd__dfrtp_4 _26594_ (.CLK(clknet_leaf_68_clk_sys),
    .D(_00217_),
    .RESET_B(net662),
    .Q(\top0.pid_q.curr_int[4] ));
 sky130_fd_sc_hd__dfrtp_4 _26595_ (.CLK(clknet_leaf_68_clk_sys),
    .D(_00218_),
    .RESET_B(net662),
    .Q(\top0.pid_q.curr_int[5] ));
 sky130_fd_sc_hd__dfrtp_4 _26596_ (.CLK(clknet_leaf_68_clk_sys),
    .D(_00219_),
    .RESET_B(net659),
    .Q(\top0.pid_q.curr_int[6] ));
 sky130_fd_sc_hd__dfrtp_4 _26597_ (.CLK(clknet_leaf_68_clk_sys),
    .D(_00220_),
    .RESET_B(net662),
    .Q(\top0.pid_q.curr_int[7] ));
 sky130_fd_sc_hd__dfrtp_2 _26598_ (.CLK(clknet_leaf_67_clk_sys),
    .D(_00221_),
    .RESET_B(net661),
    .Q(\top0.pid_q.curr_int[8] ));
 sky130_fd_sc_hd__dfrtp_4 _26599_ (.CLK(clknet_leaf_68_clk_sys),
    .D(_00222_),
    .RESET_B(net662),
    .Q(\top0.pid_q.curr_int[9] ));
 sky130_fd_sc_hd__dfrtp_4 _26600_ (.CLK(clknet_leaf_67_clk_sys),
    .D(_00223_),
    .RESET_B(net661),
    .Q(\top0.pid_q.curr_int[10] ));
 sky130_fd_sc_hd__dfrtp_4 _26601_ (.CLK(clknet_leaf_68_clk_sys),
    .D(_00224_),
    .RESET_B(net659),
    .Q(\top0.pid_q.curr_int[11] ));
 sky130_fd_sc_hd__dfrtp_4 _26602_ (.CLK(clknet_leaf_51_clk_sys),
    .D(_00225_),
    .RESET_B(net670),
    .Q(\top0.pid_q.curr_int[12] ));
 sky130_fd_sc_hd__dfrtp_4 _26603_ (.CLK(clknet_leaf_54_clk_sys),
    .D(_00226_),
    .RESET_B(net670),
    .Q(\top0.pid_q.curr_int[13] ));
 sky130_fd_sc_hd__dfrtp_4 _26604_ (.CLK(clknet_leaf_51_clk_sys),
    .D(_00227_),
    .RESET_B(net670),
    .Q(\top0.pid_q.curr_int[14] ));
 sky130_fd_sc_hd__dfrtp_2 _26605_ (.CLK(clknet_leaf_67_clk_sys),
    .D(_00228_),
    .RESET_B(net660),
    .Q(\top0.pid_q.curr_int[15] ));
 sky130_fd_sc_hd__dfstp_2 _26606_ (.CLK(clknet_leaf_86_clk_sys),
    .D(_00017_),
    .SET_B(net641),
    .Q(\top0.pid_d.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26607_ (.CLK(clknet_leaf_82_clk_sys),
    .D(_00002_),
    .RESET_B(net637),
    .Q(\top0.pid_d.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26608_ (.CLK(clknet_leaf_83_clk_sys),
    .D(_00003_),
    .RESET_B(net641),
    .Q(\top0.pid_d.state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _26609_ (.CLK(clknet_leaf_86_clk_sys),
    .D(_00004_),
    .RESET_B(net641),
    .Q(\top0.pid_d.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26610_ (.CLK(clknet_leaf_80_clk_sys),
    .D(_00005_),
    .RESET_B(net633),
    .Q(\top0.pid_d.state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26611_ (.CLK(clknet_leaf_84_clk_sys),
    .D(_00006_),
    .RESET_B(net633),
    .Q(\top0.pid_d.state[5] ));
 sky130_fd_sc_hd__dfrtp_4 _26612_ (.CLK(clknet_leaf_30_clk_sys),
    .D(_00229_),
    .RESET_B(net621),
    .Q(\top0.matmul0.beta_pass[0] ));
 sky130_fd_sc_hd__dfrtp_4 _26613_ (.CLK(clknet_leaf_30_clk_sys),
    .D(_00230_),
    .RESET_B(net623),
    .Q(\top0.matmul0.beta_pass[1] ));
 sky130_fd_sc_hd__dfrtp_4 _26614_ (.CLK(clknet_leaf_30_clk_sys),
    .D(_00231_),
    .RESET_B(net623),
    .Q(\top0.matmul0.beta_pass[2] ));
 sky130_fd_sc_hd__dfrtp_4 _26615_ (.CLK(clknet_leaf_27_clk_sys),
    .D(_00232_),
    .RESET_B(net621),
    .Q(\top0.matmul0.beta_pass[3] ));
 sky130_fd_sc_hd__dfrtp_4 _26616_ (.CLK(clknet_leaf_29_clk_sys),
    .D(_00233_),
    .RESET_B(net623),
    .Q(\top0.matmul0.beta_pass[4] ));
 sky130_fd_sc_hd__dfrtp_4 _26617_ (.CLK(clknet_leaf_28_clk_sys),
    .D(_00234_),
    .RESET_B(net621),
    .Q(\top0.matmul0.beta_pass[5] ));
 sky130_fd_sc_hd__dfrtp_4 _26618_ (.CLK(clknet_leaf_29_clk_sys),
    .D(_00235_),
    .RESET_B(net623),
    .Q(\top0.matmul0.beta_pass[6] ));
 sky130_fd_sc_hd__dfrtp_4 _26619_ (.CLK(clknet_leaf_28_clk_sys),
    .D(_00236_),
    .RESET_B(net623),
    .Q(\top0.matmul0.beta_pass[7] ));
 sky130_fd_sc_hd__dfrtp_4 _26620_ (.CLK(clknet_leaf_28_clk_sys),
    .D(_00237_),
    .RESET_B(net622),
    .Q(\top0.matmul0.beta_pass[8] ));
 sky130_fd_sc_hd__dfrtp_4 _26621_ (.CLK(clknet_leaf_25_clk_sys),
    .D(_00238_),
    .RESET_B(net627),
    .Q(\top0.matmul0.beta_pass[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26622_ (.CLK(clknet_leaf_25_clk_sys),
    .D(_00239_),
    .RESET_B(net627),
    .Q(\top0.matmul0.beta_pass[10] ));
 sky130_fd_sc_hd__dfrtp_4 _26623_ (.CLK(clknet_leaf_29_clk_sys),
    .D(_00240_),
    .RESET_B(net623),
    .Q(\top0.matmul0.beta_pass[11] ));
 sky130_fd_sc_hd__dfrtp_4 _26624_ (.CLK(clknet_leaf_29_clk_sys),
    .D(_00241_),
    .RESET_B(net624),
    .Q(\top0.matmul0.beta_pass[12] ));
 sky130_fd_sc_hd__dfrtp_4 _26625_ (.CLK(clknet_leaf_31_clk_sys),
    .D(_00242_),
    .RESET_B(net619),
    .Q(\top0.matmul0.beta_pass[13] ));
 sky130_fd_sc_hd__dfrtp_2 _26626_ (.CLK(clknet_leaf_25_clk_sys),
    .D(_00243_),
    .RESET_B(net627),
    .Q(\top0.matmul0.beta_pass[14] ));
 sky130_fd_sc_hd__dfrtp_4 _26627_ (.CLK(clknet_leaf_25_clk_sys),
    .D(_00244_),
    .RESET_B(net628),
    .Q(\top0.matmul0.beta_pass[15] ));
 sky130_fd_sc_hd__dfrtp_4 _26628_ (.CLK(clknet_leaf_72_clk_sys),
    .D(_00245_),
    .RESET_B(net655),
    .Q(\top0.pid_d.out[0] ));
 sky130_fd_sc_hd__dfrtp_4 _26629_ (.CLK(clknet_leaf_64_clk_sys),
    .D(_00246_),
    .RESET_B(net656),
    .Q(\top0.pid_d.out[1] ));
 sky130_fd_sc_hd__dfrtp_4 _26630_ (.CLK(clknet_leaf_74_clk_sys),
    .D(_00247_),
    .RESET_B(net655),
    .Q(\top0.pid_d.out[2] ));
 sky130_fd_sc_hd__dfrtp_4 _26631_ (.CLK(clknet_leaf_82_clk_sys),
    .D(_00248_),
    .RESET_B(net637),
    .Q(\top0.pid_d.out[3] ));
 sky130_fd_sc_hd__dfrtp_4 _26632_ (.CLK(clknet_leaf_74_clk_sys),
    .D(_00249_),
    .RESET_B(net655),
    .Q(\top0.pid_d.out[4] ));
 sky130_fd_sc_hd__dfrtp_4 _26633_ (.CLK(clknet_leaf_82_clk_sys),
    .D(_00250_),
    .RESET_B(net638),
    .Q(\top0.pid_d.out[5] ));
 sky130_fd_sc_hd__dfrtp_4 _26634_ (.CLK(clknet_leaf_74_clk_sys),
    .D(_00251_),
    .RESET_B(net637),
    .Q(\top0.pid_d.out[6] ));
 sky130_fd_sc_hd__dfrtp_4 _26635_ (.CLK(clknet_leaf_75_clk_sys),
    .D(_00252_),
    .RESET_B(net637),
    .Q(\top0.pid_d.out[7] ));
 sky130_fd_sc_hd__dfrtp_2 _26636_ (.CLK(clknet_leaf_81_clk_sys),
    .D(_00253_),
    .RESET_B(net636),
    .Q(\top0.pid_d.out[8] ));
 sky130_fd_sc_hd__dfrtp_2 _26637_ (.CLK(clknet_leaf_82_clk_sys),
    .D(_00254_),
    .RESET_B(net638),
    .Q(\top0.pid_d.out[9] ));
 sky130_fd_sc_hd__dfrtp_2 _26638_ (.CLK(clknet_leaf_80_clk_sys),
    .D(_00255_),
    .RESET_B(net633),
    .Q(\top0.pid_d.out[10] ));
 sky130_fd_sc_hd__dfrtp_4 _26639_ (.CLK(clknet_leaf_81_clk_sys),
    .D(_00256_),
    .RESET_B(net638),
    .Q(\top0.pid_d.out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26640_ (.CLK(clknet_leaf_80_clk_sys),
    .D(_00257_),
    .RESET_B(net633),
    .Q(\top0.pid_d.out[12] ));
 sky130_fd_sc_hd__dfrtp_4 _26641_ (.CLK(clknet_leaf_80_clk_sys),
    .D(_00258_),
    .RESET_B(net634),
    .Q(\top0.pid_d.out[13] ));
 sky130_fd_sc_hd__dfrtp_4 _26642_ (.CLK(clknet_leaf_80_clk_sys),
    .D(_00259_),
    .RESET_B(net634),
    .Q(\top0.pid_d.out[14] ));
 sky130_fd_sc_hd__dfrtp_4 _26643_ (.CLK(clknet_leaf_78_clk_sys),
    .D(_00260_),
    .RESET_B(net632),
    .Q(\top0.pid_d.out[15] ));
 sky130_fd_sc_hd__dfrtp_1 _26644_ (.CLK(clknet_leaf_86_clk_sys),
    .D(_00261_),
    .RESET_B(net640),
    .Q(\top0.pid_d.out_valid ));
 sky130_fd_sc_hd__dfrtp_4 _26645_ (.CLK(clknet_leaf_75_clk_sys),
    .D(_00262_),
    .RESET_B(net639),
    .Q(\top0.pid_d.mult0.a[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26646_ (.CLK(clknet_leaf_75_clk_sys),
    .D(_00263_),
    .RESET_B(net637),
    .Q(\top0.pid_d.mult0.a[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26647_ (.CLK(clknet_leaf_76_clk_sys),
    .D(_00264_),
    .RESET_B(net639),
    .Q(\top0.pid_d.mult0.a[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26648_ (.CLK(clknet_leaf_75_clk_sys),
    .D(_00265_),
    .RESET_B(net639),
    .Q(\top0.pid_d.mult0.a[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26649_ (.CLK(clknet_leaf_75_clk_sys),
    .D(_00266_),
    .RESET_B(net639),
    .Q(\top0.pid_d.mult0.a[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26650_ (.CLK(clknet_leaf_76_clk_sys),
    .D(_00267_),
    .RESET_B(net639),
    .Q(\top0.pid_d.mult0.a[5] ));
 sky130_fd_sc_hd__dfrtp_4 _26651_ (.CLK(clknet_leaf_75_clk_sys),
    .D(_00268_),
    .RESET_B(net639),
    .Q(\top0.pid_d.mult0.a[6] ));
 sky130_fd_sc_hd__dfrtp_2 _26652_ (.CLK(clknet_leaf_75_clk_sys),
    .D(_00269_),
    .RESET_B(net639),
    .Q(\top0.pid_d.mult0.a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26653_ (.CLK(clknet_leaf_75_clk_sys),
    .D(_00270_),
    .RESET_B(net636),
    .Q(\top0.pid_d.mult0.a[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26654_ (.CLK(clknet_leaf_76_clk_sys),
    .D(_00271_),
    .RESET_B(net639),
    .Q(\top0.pid_d.mult0.a[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26655_ (.CLK(clknet_leaf_81_clk_sys),
    .D(_00272_),
    .RESET_B(net633),
    .Q(\top0.pid_d.mult0.a[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26656_ (.CLK(clknet_leaf_79_clk_sys),
    .D(_00273_),
    .RESET_B(net632),
    .Q(\top0.pid_d.mult0.a[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26657_ (.CLK(clknet_leaf_78_clk_sys),
    .D(_00274_),
    .RESET_B(net631),
    .Q(\top0.pid_d.mult0.a[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26658_ (.CLK(clknet_leaf_77_clk_sys),
    .D(_00275_),
    .RESET_B(net635),
    .Q(\top0.pid_d.mult0.a[13] ));
 sky130_fd_sc_hd__dfrtp_4 _26659_ (.CLK(clknet_leaf_77_clk_sys),
    .D(_00276_),
    .RESET_B(net635),
    .Q(\top0.pid_d.mult0.a[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26660_ (.CLK(clknet_leaf_77_clk_sys),
    .D(_00277_),
    .RESET_B(net635),
    .Q(\top0.pid_d.mult0.a[15] ));
 sky130_fd_sc_hd__dfrtp_1 _26661_ (.CLK(clknet_leaf_75_clk_sys),
    .D(_00278_),
    .RESET_B(net637),
    .Q(\top0.pid_d.mult0.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26662_ (.CLK(clknet_leaf_75_clk_sys),
    .D(_00279_),
    .RESET_B(net637),
    .Q(\top0.pid_d.mult0.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26663_ (.CLK(clknet_leaf_63_clk_sys),
    .D(_00280_),
    .RESET_B(net656),
    .Q(\top0.pid_d.mult0.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26664_ (.CLK(clknet_leaf_63_clk_sys),
    .D(_00281_),
    .RESET_B(net656),
    .Q(\top0.pid_d.mult0.b[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26665_ (.CLK(clknet_leaf_75_clk_sys),
    .D(_00282_),
    .RESET_B(net637),
    .Q(\top0.pid_d.mult0.b[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26666_ (.CLK(clknet_leaf_82_clk_sys),
    .D(_00283_),
    .RESET_B(net647),
    .Q(\top0.pid_d.mult0.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26667_ (.CLK(clknet_leaf_82_clk_sys),
    .D(_00284_),
    .RESET_B(net647),
    .Q(\top0.pid_d.mult0.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26668_ (.CLK(clknet_leaf_82_clk_sys),
    .D(_00285_),
    .RESET_B(net647),
    .Q(\top0.pid_d.mult0.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26669_ (.CLK(clknet_leaf_82_clk_sys),
    .D(_00286_),
    .RESET_B(net646),
    .Q(\top0.pid_d.mult0.b[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26670_ (.CLK(clknet_leaf_82_clk_sys),
    .D(_00287_),
    .RESET_B(net647),
    .Q(\top0.pid_d.mult0.b[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26671_ (.CLK(clknet_leaf_82_clk_sys),
    .D(_00288_),
    .RESET_B(net646),
    .Q(\top0.pid_d.mult0.b[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26672_ (.CLK(clknet_leaf_82_clk_sys),
    .D(_00289_),
    .RESET_B(net646),
    .Q(\top0.pid_d.mult0.b[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26673_ (.CLK(clknet_leaf_81_clk_sys),
    .D(_00290_),
    .RESET_B(net636),
    .Q(\top0.pid_d.mult0.b[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26674_ (.CLK(clknet_leaf_81_clk_sys),
    .D(_00291_),
    .RESET_B(net636),
    .Q(\top0.pid_d.mult0.b[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26675_ (.CLK(clknet_leaf_81_clk_sys),
    .D(_00292_),
    .RESET_B(net636),
    .Q(\top0.pid_d.mult0.b[14] ));
 sky130_fd_sc_hd__dfrtp_2 _26676_ (.CLK(clknet_leaf_81_clk_sys),
    .D(_00293_),
    .RESET_B(net636),
    .Q(\top0.pid_d.mult0.b[15] ));
 sky130_fd_sc_hd__dfrtp_2 _26677_ (.CLK(clknet_leaf_64_clk_sys),
    .D(_00294_),
    .RESET_B(net656),
    .Q(\top0.pid_d.curr_error[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26678_ (.CLK(clknet_leaf_64_clk_sys),
    .D(_00295_),
    .RESET_B(net656),
    .Q(\top0.pid_d.curr_error[1] ));
 sky130_fd_sc_hd__dfrtp_2 _26679_ (.CLK(clknet_leaf_64_clk_sys),
    .D(_00296_),
    .RESET_B(net656),
    .Q(\top0.pid_d.curr_error[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26680_ (.CLK(clknet_leaf_64_clk_sys),
    .D(_00297_),
    .RESET_B(net656),
    .Q(\top0.pid_d.curr_error[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26681_ (.CLK(clknet_leaf_63_clk_sys),
    .D(_00298_),
    .RESET_B(net647),
    .Q(\top0.pid_d.curr_error[4] ));
 sky130_fd_sc_hd__dfrtp_2 _26682_ (.CLK(clknet_leaf_62_clk_sys),
    .D(_00299_),
    .RESET_B(net648),
    .Q(\top0.pid_d.curr_error[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26683_ (.CLK(clknet_leaf_62_clk_sys),
    .D(_00300_),
    .RESET_B(net648),
    .Q(\top0.pid_d.curr_error[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26684_ (.CLK(clknet_leaf_62_clk_sys),
    .D(_00301_),
    .RESET_B(net646),
    .Q(\top0.pid_d.curr_error[7] ));
 sky130_fd_sc_hd__dfrtp_2 _26685_ (.CLK(clknet_leaf_62_clk_sys),
    .D(_00302_),
    .RESET_B(net646),
    .Q(\top0.pid_d.curr_error[8] ));
 sky130_fd_sc_hd__dfrtp_2 _26686_ (.CLK(clknet_leaf_83_clk_sys),
    .D(_00303_),
    .RESET_B(net647),
    .Q(\top0.pid_d.curr_error[9] ));
 sky130_fd_sc_hd__dfrtp_2 _26687_ (.CLK(clknet_leaf_83_clk_sys),
    .D(_00304_),
    .RESET_B(net646),
    .Q(\top0.pid_d.curr_error[10] ));
 sky130_fd_sc_hd__dfrtp_2 _26688_ (.CLK(clknet_leaf_83_clk_sys),
    .D(_00305_),
    .RESET_B(net649),
    .Q(\top0.pid_d.curr_error[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26689_ (.CLK(clknet_leaf_84_clk_sys),
    .D(_00306_),
    .RESET_B(net641),
    .Q(\top0.pid_d.curr_error[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26690_ (.CLK(clknet_leaf_84_clk_sys),
    .D(_00307_),
    .RESET_B(net641),
    .Q(\top0.pid_d.curr_error[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26691_ (.CLK(clknet_leaf_83_clk_sys),
    .D(_00308_),
    .RESET_B(net641),
    .Q(\top0.pid_d.curr_error[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26692_ (.CLK(clknet_leaf_83_clk_sys),
    .D(_00309_),
    .RESET_B(net641),
    .Q(\top0.pid_d.curr_error[15] ));
 sky130_fd_sc_hd__dfrtp_2 _26693_ (.CLK(clknet_leaf_64_clk_sys),
    .D(_00310_),
    .RESET_B(net658),
    .Q(\top0.pid_d.prev_error[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26694_ (.CLK(clknet_leaf_71_clk_sys),
    .D(_00311_),
    .RESET_B(net657),
    .Q(\top0.pid_d.prev_error[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26695_ (.CLK(clknet_leaf_71_clk_sys),
    .D(net893),
    .RESET_B(net657),
    .Q(\top0.pid_d.prev_error[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26696_ (.CLK(clknet_leaf_64_clk_sys),
    .D(_00313_),
    .RESET_B(net656),
    .Q(\top0.pid_d.prev_error[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26697_ (.CLK(clknet_leaf_63_clk_sys),
    .D(_00314_),
    .RESET_B(net647),
    .Q(\top0.pid_d.prev_error[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26698_ (.CLK(clknet_leaf_64_clk_sys),
    .D(_00315_),
    .RESET_B(net648),
    .Q(\top0.pid_d.prev_error[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26699_ (.CLK(clknet_leaf_63_clk_sys),
    .D(_00316_),
    .RESET_B(net648),
    .Q(\top0.pid_d.prev_error[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26700_ (.CLK(clknet_leaf_62_clk_sys),
    .D(net881),
    .RESET_B(net648),
    .Q(\top0.pid_d.prev_error[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26701_ (.CLK(clknet_leaf_83_clk_sys),
    .D(net877),
    .RESET_B(net649),
    .Q(\top0.pid_d.prev_error[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26702_ (.CLK(clknet_leaf_82_clk_sys),
    .D(net890),
    .RESET_B(net646),
    .Q(\top0.pid_d.prev_error[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26703_ (.CLK(clknet_leaf_83_clk_sys),
    .D(net875),
    .RESET_B(net646),
    .Q(\top0.pid_d.prev_error[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26704_ (.CLK(clknet_leaf_84_clk_sys),
    .D(_00321_),
    .RESET_B(net646),
    .Q(\top0.pid_d.prev_error[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26705_ (.CLK(clknet_leaf_84_clk_sys),
    .D(net904),
    .RESET_B(net641),
    .Q(\top0.pid_d.prev_error[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26706_ (.CLK(clknet_leaf_84_clk_sys),
    .D(_00323_),
    .RESET_B(net641),
    .Q(\top0.pid_d.prev_error[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26707_ (.CLK(clknet_leaf_85_clk_sys),
    .D(net766),
    .RESET_B(net641),
    .Q(\top0.pid_d.prev_error[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26708_ (.CLK(clknet_leaf_84_clk_sys),
    .D(net723),
    .RESET_B(net645),
    .Q(\top0.pid_d.prev_error[15] ));
 sky130_fd_sc_hd__dfrtp_4 _26709_ (.CLK(clknet_leaf_71_clk_sys),
    .D(_00326_),
    .RESET_B(net657),
    .Q(\top0.pid_d.curr_int[0] ));
 sky130_fd_sc_hd__dfrtp_4 _26710_ (.CLK(clknet_leaf_71_clk_sys),
    .D(_00327_),
    .RESET_B(net657),
    .Q(\top0.pid_d.curr_int[1] ));
 sky130_fd_sc_hd__dfrtp_4 _26711_ (.CLK(clknet_leaf_72_clk_sys),
    .D(_00328_),
    .RESET_B(net655),
    .Q(\top0.pid_d.curr_int[2] ));
 sky130_fd_sc_hd__dfrtp_4 _26712_ (.CLK(clknet_leaf_72_clk_sys),
    .D(_00329_),
    .RESET_B(net655),
    .Q(\top0.pid_d.curr_int[3] ));
 sky130_fd_sc_hd__dfrtp_4 _26713_ (.CLK(clknet_leaf_72_clk_sys),
    .D(_00330_),
    .RESET_B(net663),
    .Q(\top0.pid_d.curr_int[4] ));
 sky130_fd_sc_hd__dfrtp_4 _26714_ (.CLK(clknet_leaf_73_clk_sys),
    .D(_00331_),
    .RESET_B(net655),
    .Q(\top0.pid_d.curr_int[5] ));
 sky130_fd_sc_hd__dfrtp_4 _26715_ (.CLK(clknet_leaf_74_clk_sys),
    .D(_00332_),
    .RESET_B(net638),
    .Q(\top0.pid_d.curr_int[6] ));
 sky130_fd_sc_hd__dfrtp_4 _26716_ (.CLK(clknet_leaf_74_clk_sys),
    .D(_00333_),
    .RESET_B(net638),
    .Q(\top0.pid_d.curr_int[7] ));
 sky130_fd_sc_hd__dfrtp_4 _26717_ (.CLK(clknet_leaf_75_clk_sys),
    .D(_00334_),
    .RESET_B(net636),
    .Q(\top0.pid_d.curr_int[8] ));
 sky130_fd_sc_hd__dfrtp_2 _26718_ (.CLK(clknet_leaf_82_clk_sys),
    .D(_00335_),
    .RESET_B(net638),
    .Q(\top0.pid_d.curr_int[9] ));
 sky130_fd_sc_hd__dfrtp_2 _26719_ (.CLK(clknet_leaf_81_clk_sys),
    .D(_00336_),
    .RESET_B(net634),
    .Q(\top0.pid_d.curr_int[10] ));
 sky130_fd_sc_hd__dfrtp_4 _26720_ (.CLK(clknet_leaf_82_clk_sys),
    .D(_00337_),
    .RESET_B(net638),
    .Q(\top0.pid_d.curr_int[11] ));
 sky130_fd_sc_hd__dfrtp_4 _26721_ (.CLK(clknet_leaf_81_clk_sys),
    .D(_00338_),
    .RESET_B(net636),
    .Q(\top0.pid_d.curr_int[12] ));
 sky130_fd_sc_hd__dfrtp_4 _26722_ (.CLK(clknet_leaf_78_clk_sys),
    .D(_00339_),
    .RESET_B(net633),
    .Q(\top0.pid_d.curr_int[13] ));
 sky130_fd_sc_hd__dfrtp_4 _26723_ (.CLK(clknet_leaf_78_clk_sys),
    .D(_00340_),
    .RESET_B(net633),
    .Q(\top0.pid_d.curr_int[14] ));
 sky130_fd_sc_hd__dfrtp_2 _26724_ (.CLK(clknet_leaf_78_clk_sys),
    .D(_00341_),
    .RESET_B(net633),
    .Q(\top0.pid_d.curr_int[15] ));
 sky130_fd_sc_hd__dfstp_1 _26725_ (.CLK(clknet_leaf_103_clk_sys),
    .D(_00342_),
    .SET_B(net576),
    .Q(\top0.cordic0.vec[0][0] ));
 sky130_fd_sc_hd__dfstp_1 _26726_ (.CLK(clknet_leaf_104_clk_sys),
    .D(_00343_),
    .SET_B(net576),
    .Q(\top0.cordic0.vec[0][1] ));
 sky130_fd_sc_hd__dfstp_1 _26727_ (.CLK(clknet_leaf_104_clk_sys),
    .D(_00344_),
    .SET_B(net576),
    .Q(\top0.cordic0.vec[0][2] ));
 sky130_fd_sc_hd__dfstp_1 _26728_ (.CLK(clknet_leaf_104_clk_sys),
    .D(_00345_),
    .SET_B(net576),
    .Q(\top0.cordic0.vec[0][3] ));
 sky130_fd_sc_hd__dfstp_1 _26729_ (.CLK(clknet_leaf_104_clk_sys),
    .D(_00346_),
    .SET_B(net576),
    .Q(\top0.cordic0.vec[0][4] ));
 sky130_fd_sc_hd__dfstp_1 _26730_ (.CLK(clknet_leaf_100_clk_sys),
    .D(_00347_),
    .SET_B(net576),
    .Q(\top0.cordic0.vec[0][5] ));
 sky130_fd_sc_hd__dfstp_1 _26731_ (.CLK(clknet_leaf_103_clk_sys),
    .D(_00348_),
    .SET_B(net576),
    .Q(\top0.cordic0.vec[0][6] ));
 sky130_fd_sc_hd__dfstp_1 _26732_ (.CLK(clknet_leaf_103_clk_sys),
    .D(_00349_),
    .SET_B(net576),
    .Q(\top0.cordic0.vec[0][7] ));
 sky130_fd_sc_hd__dfstp_1 _26733_ (.CLK(clknet_leaf_100_clk_sys),
    .D(_00350_),
    .SET_B(net587),
    .Q(\top0.cordic0.vec[0][8] ));
 sky130_fd_sc_hd__dfstp_1 _26734_ (.CLK(clknet_leaf_100_clk_sys),
    .D(_00351_),
    .SET_B(net587),
    .Q(\top0.cordic0.vec[0][9] ));
 sky130_fd_sc_hd__dfstp_2 _26735_ (.CLK(clknet_leaf_100_clk_sys),
    .D(_00352_),
    .SET_B(net587),
    .Q(\top0.cordic0.vec[0][10] ));
 sky130_fd_sc_hd__dfstp_1 _26736_ (.CLK(clknet_leaf_101_clk_sys),
    .D(_00353_),
    .SET_B(net587),
    .Q(\top0.cordic0.vec[0][11] ));
 sky130_fd_sc_hd__dfstp_1 _26737_ (.CLK(clknet_leaf_101_clk_sys),
    .D(_00354_),
    .SET_B(net587),
    .Q(\top0.cordic0.vec[0][12] ));
 sky130_fd_sc_hd__dfstp_1 _26738_ (.CLK(clknet_leaf_101_clk_sys),
    .D(_00355_),
    .SET_B(net587),
    .Q(\top0.cordic0.vec[0][13] ));
 sky130_fd_sc_hd__dfstp_1 _26739_ (.CLK(clknet_leaf_96_clk_sys),
    .D(_00356_),
    .SET_B(net587),
    .Q(\top0.cordic0.vec[0][14] ));
 sky130_fd_sc_hd__dfstp_1 _26740_ (.CLK(clknet_leaf_101_clk_sys),
    .D(_00357_),
    .SET_B(net587),
    .Q(\top0.cordic0.vec[0][15] ));
 sky130_fd_sc_hd__dfrtp_1 _26741_ (.CLK(clknet_leaf_96_clk_sys),
    .D(_00358_),
    .RESET_B(net587),
    .Q(\top0.cordic0.vec[0][16] ));
 sky130_fd_sc_hd__dfrtp_1 _26742_ (.CLK(clknet_leaf_96_clk_sys),
    .D(_00359_),
    .RESET_B(net587),
    .Q(\top0.cordic0.vec[0][17] ));
 sky130_fd_sc_hd__dfrtp_1 _26743_ (.CLK(clknet_leaf_96_clk_sys),
    .D(_00360_),
    .RESET_B(net588),
    .Q(\top0.cordic0.slte0.opA[0] ));
 sky130_fd_sc_hd__dfrtp_4 _26744_ (.CLK(clknet_leaf_96_clk_sys),
    .D(_00361_),
    .RESET_B(net588),
    .Q(\top0.cordic0.slte0.opA[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26745_ (.CLK(clknet_leaf_96_clk_sys),
    .D(_00362_),
    .RESET_B(net588),
    .Q(\top0.cordic0.slte0.opA[2] ));
 sky130_fd_sc_hd__dfrtp_4 _26746_ (.CLK(clknet_leaf_97_clk_sys),
    .D(_00363_),
    .RESET_B(net588),
    .Q(\top0.cordic0.slte0.opA[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26747_ (.CLK(clknet_leaf_92_clk_sys),
    .D(_00364_),
    .RESET_B(net599),
    .Q(\top0.cordic0.slte0.opA[4] ));
 sky130_fd_sc_hd__dfrtp_4 _26748_ (.CLK(clknet_leaf_97_clk_sys),
    .D(_00365_),
    .RESET_B(net588),
    .Q(\top0.cordic0.slte0.opA[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26749_ (.CLK(clknet_leaf_92_clk_sys),
    .D(_00366_),
    .RESET_B(net599),
    .Q(\top0.cordic0.slte0.opA[6] ));
 sky130_fd_sc_hd__dfrtp_4 _26750_ (.CLK(clknet_leaf_92_clk_sys),
    .D(_00367_),
    .RESET_B(net599),
    .Q(\top0.cordic0.slte0.opA[7] ));
 sky130_fd_sc_hd__dfrtp_4 _26751_ (.CLK(clknet_leaf_94_clk_sys),
    .D(_00368_),
    .RESET_B(net591),
    .Q(\top0.cordic0.slte0.opA[8] ));
 sky130_fd_sc_hd__dfrtp_4 _26752_ (.CLK(clknet_leaf_94_clk_sys),
    .D(_00369_),
    .RESET_B(net591),
    .Q(\top0.cordic0.slte0.opA[9] ));
 sky130_fd_sc_hd__dfrtp_2 _26753_ (.CLK(clknet_leaf_93_clk_sys),
    .D(_00370_),
    .RESET_B(net591),
    .Q(\top0.cordic0.slte0.opA[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26754_ (.CLK(clknet_leaf_6_clk_sys),
    .D(_00371_),
    .RESET_B(net591),
    .Q(\top0.cordic0.slte0.opA[11] ));
 sky130_fd_sc_hd__dfrtp_2 _26755_ (.CLK(clknet_leaf_5_clk_sys),
    .D(_00372_),
    .RESET_B(net590),
    .Q(\top0.cordic0.slte0.opA[12] ));
 sky130_fd_sc_hd__dfrtp_4 _26756_ (.CLK(clknet_leaf_5_clk_sys),
    .D(_00373_),
    .RESET_B(net590),
    .Q(\top0.cordic0.slte0.opA[13] ));
 sky130_fd_sc_hd__dfrtp_4 _26757_ (.CLK(clknet_leaf_94_clk_sys),
    .D(_00374_),
    .RESET_B(net591),
    .Q(\top0.cordic0.slte0.opA[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26758_ (.CLK(clknet_leaf_5_clk_sys),
    .D(_00375_),
    .RESET_B(net590),
    .Q(\top0.cordic0.slte0.opA[15] ));
 sky130_fd_sc_hd__dfrtp_1 _26759_ (.CLK(clknet_leaf_94_clk_sys),
    .D(_00376_),
    .RESET_B(net590),
    .Q(\top0.cordic0.slte0.opA[16] ));
 sky130_fd_sc_hd__dfrtp_2 _26760_ (.CLK(clknet_3_0__leaf_clk_sys),
    .D(_00377_),
    .RESET_B(net589),
    .Q(\top0.cordic0.slte0.opA[17] ));
 sky130_fd_sc_hd__dfrtp_1 _26761_ (.CLK(clknet_leaf_7_clk_sys),
    .D(_00378_),
    .RESET_B(net593),
    .Q(\top0.cordic0.domain[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26762_ (.CLK(clknet_leaf_93_clk_sys),
    .D(_00379_),
    .RESET_B(net599),
    .Q(\top0.cordic0.domain[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26763_ (.CLK(clknet_leaf_87_clk_sys),
    .D(_00380_),
    .RESET_B(net645),
    .Q(\top0.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26764_ (.CLK(clknet_leaf_87_clk_sys),
    .D(_00381_),
    .RESET_B(net642),
    .Q(\top0.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26765_ (.CLK(clknet_leaf_87_clk_sys),
    .D(_00382_),
    .RESET_B(net642),
    .Q(\top0.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26766_ (.CLK(clknet_leaf_4_clk_sys),
    .D(_00383_),
    .RESET_B(net580),
    .Q(\top0.cordic0.cos[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26767_ (.CLK(clknet_leaf_4_clk_sys),
    .D(_00384_),
    .RESET_B(net580),
    .Q(\top0.cordic0.cos[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26768_ (.CLK(clknet_leaf_4_clk_sys),
    .D(_00385_),
    .RESET_B(net580),
    .Q(\top0.cordic0.cos[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26769_ (.CLK(clknet_leaf_5_clk_sys),
    .D(_00386_),
    .RESET_B(net590),
    .Q(\top0.cordic0.cos[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26770_ (.CLK(clknet_leaf_4_clk_sys),
    .D(_00387_),
    .RESET_B(net580),
    .Q(\top0.cordic0.cos[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26771_ (.CLK(clknet_leaf_6_clk_sys),
    .D(_00388_),
    .RESET_B(net590),
    .Q(\top0.cordic0.cos[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26772_ (.CLK(clknet_leaf_7_clk_sys),
    .D(_00389_),
    .RESET_B(net593),
    .Q(\top0.cordic0.cos[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26773_ (.CLK(clknet_leaf_6_clk_sys),
    .D(_00390_),
    .RESET_B(net590),
    .Q(\top0.cordic0.cos[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26774_ (.CLK(clknet_leaf_4_clk_sys),
    .D(_00391_),
    .RESET_B(net580),
    .Q(\top0.cordic0.cos[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26775_ (.CLK(clknet_leaf_7_clk_sys),
    .D(_00392_),
    .RESET_B(net593),
    .Q(\top0.cordic0.cos[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26776_ (.CLK(clknet_leaf_5_clk_sys),
    .D(_00393_),
    .RESET_B(net590),
    .Q(\top0.cordic0.cos[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26777_ (.CLK(clknet_leaf_7_clk_sys),
    .D(_00394_),
    .RESET_B(net593),
    .Q(\top0.cordic0.cos[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26778_ (.CLK(clknet_leaf_6_clk_sys),
    .D(_00395_),
    .RESET_B(net591),
    .Q(\top0.cordic0.cos[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26779_ (.CLK(clknet_leaf_6_clk_sys),
    .D(_00396_),
    .RESET_B(net590),
    .Q(\top0.cordic0.cos[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26780_ (.CLK(clknet_leaf_109_clk_sys),
    .D(_00397_),
    .RESET_B(net579),
    .Q(\top0.cordic0.sin[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26781_ (.CLK(clknet_leaf_109_clk_sys),
    .D(_00398_),
    .RESET_B(net579),
    .Q(\top0.cordic0.sin[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26782_ (.CLK(clknet_leaf_110_clk_sys),
    .D(_00399_),
    .RESET_B(net579),
    .Q(\top0.cordic0.sin[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26783_ (.CLK(clknet_leaf_109_clk_sys),
    .D(_00400_),
    .RESET_B(net579),
    .Q(\top0.cordic0.sin[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26784_ (.CLK(clknet_leaf_109_clk_sys),
    .D(_00401_),
    .RESET_B(net578),
    .Q(\top0.cordic0.sin[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26785_ (.CLK(clknet_leaf_3_clk_sys),
    .D(_00402_),
    .RESET_B(net582),
    .Q(\top0.cordic0.sin[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26786_ (.CLK(clknet_leaf_1_clk_sys),
    .D(_00403_),
    .RESET_B(net582),
    .Q(\top0.cordic0.sin[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26787_ (.CLK(clknet_leaf_3_clk_sys),
    .D(_00404_),
    .RESET_B(net583),
    .Q(\top0.cordic0.sin[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26788_ (.CLK(clknet_leaf_3_clk_sys),
    .D(_00405_),
    .RESET_B(net583),
    .Q(\top0.cordic0.sin[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26789_ (.CLK(clknet_leaf_3_clk_sys),
    .D(_00406_),
    .RESET_B(net583),
    .Q(\top0.cordic0.sin[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26790_ (.CLK(clknet_leaf_1_clk_sys),
    .D(_00407_),
    .RESET_B(net582),
    .Q(\top0.cordic0.sin[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26791_ (.CLK(clknet_leaf_1_clk_sys),
    .D(_00408_),
    .RESET_B(net578),
    .Q(\top0.cordic0.sin[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26792_ (.CLK(clknet_leaf_0_clk_sys),
    .D(_00409_),
    .RESET_B(net578),
    .Q(\top0.cordic0.sin[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26793_ (.CLK(clknet_leaf_109_clk_sys),
    .D(_00410_),
    .RESET_B(net578),
    .Q(\top0.cordic0.sin[13] ));
 sky130_fd_sc_hd__dfrtp_2 _26794_ (.CLK(clknet_leaf_92_clk_sys),
    .D(_00411_),
    .RESET_B(net599),
    .Q(\top0.cordic0.out_valid ));
 sky130_fd_sc_hd__dfrtp_4 _26795_ (.CLK(clknet_leaf_88_clk_sys),
    .D(_00412_),
    .RESET_B(net642),
    .Q(\top0.start_svm ));
 sky130_fd_sc_hd__dfrtp_1 _26796_ (.CLK(clknet_leaf_104_clk_sys),
    .D(_00413_),
    .RESET_B(net576),
    .Q(\top0.cordic0.gm0.iter[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26797_ (.CLK(clknet_leaf_105_clk_sys),
    .D(_00414_),
    .RESET_B(net576),
    .Q(\top0.cordic0.gm0.iter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26798_ (.CLK(clknet_leaf_102_clk_sys),
    .D(_00415_),
    .RESET_B(net589),
    .Q(\top0.cordic0.gm0.iter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26799_ (.CLK(clknet_leaf_102_clk_sys),
    .D(_00416_),
    .RESET_B(net589),
    .Q(\top0.cordic0.gm0.iter[3] ));
 sky130_fd_sc_hd__dfrtp_2 _26800_ (.CLK(clknet_leaf_108_clk_sys),
    .D(_00417_),
    .RESET_B(net606),
    .Q(\top0.cordic0.gm0.iter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26801_ (.CLK(clknet_leaf_6_clk_sys),
    .D(_00418_),
    .RESET_B(net591),
    .Q(\top0.cordic0.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26802_ (.CLK(clknet_leaf_64_clk_sys),
    .D(_00419_),
    .RESET_B(net658),
    .Q(\top0.pid_q.prev_int[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26803_ (.CLK(clknet_leaf_65_clk_sys),
    .D(_00420_),
    .RESET_B(net657),
    .Q(\top0.pid_q.prev_int[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26804_ (.CLK(clknet_leaf_71_clk_sys),
    .D(_00421_),
    .RESET_B(net658),
    .Q(\top0.pid_q.prev_int[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26805_ (.CLK(clknet_leaf_70_clk_sys),
    .D(_00422_),
    .RESET_B(net658),
    .Q(\top0.pid_q.prev_int[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26806_ (.CLK(clknet_leaf_70_clk_sys),
    .D(_00423_),
    .RESET_B(net662),
    .Q(\top0.pid_q.prev_int[4] ));
 sky130_fd_sc_hd__dfrtp_4 _26807_ (.CLK(clknet_leaf_69_clk_sys),
    .D(_00424_),
    .RESET_B(net662),
    .Q(\top0.pid_q.prev_int[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26808_ (.CLK(clknet_leaf_68_clk_sys),
    .D(_00425_),
    .RESET_B(net662),
    .Q(\top0.pid_q.prev_int[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26809_ (.CLK(clknet_leaf_68_clk_sys),
    .D(_00426_),
    .RESET_B(net662),
    .Q(\top0.pid_q.prev_int[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26810_ (.CLK(clknet_leaf_68_clk_sys),
    .D(_00427_),
    .RESET_B(net663),
    .Q(\top0.pid_q.prev_int[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26811_ (.CLK(clknet_leaf_69_clk_sys),
    .D(_00428_),
    .RESET_B(net663),
    .Q(\top0.pid_q.prev_int[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26812_ (.CLK(clknet_leaf_51_clk_sys),
    .D(_00429_),
    .RESET_B(net670),
    .Q(\top0.pid_q.prev_int[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26813_ (.CLK(clknet_leaf_67_clk_sys),
    .D(_00430_),
    .RESET_B(net660),
    .Q(\top0.pid_q.prev_int[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26814_ (.CLK(clknet_leaf_51_clk_sys),
    .D(_00431_),
    .RESET_B(net670),
    .Q(\top0.pid_q.prev_int[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26815_ (.CLK(clknet_leaf_55_clk_sys),
    .D(_00432_),
    .RESET_B(net667),
    .Q(\top0.pid_q.prev_int[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26816_ (.CLK(clknet_leaf_60_clk_sys),
    .D(_00433_),
    .RESET_B(net652),
    .Q(\top0.pid_q.prev_int[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26817_ (.CLK(clknet_leaf_60_clk_sys),
    .D(net773),
    .RESET_B(net652),
    .Q(\top0.pid_q.prev_int[15] ));
 sky130_fd_sc_hd__dfrtp_4 _26818_ (.CLK(clknet_leaf_47_clk_sys),
    .D(_00435_),
    .RESET_B(net676),
    .Q(\top0.svm0.out_valid ));
 sky130_fd_sc_hd__dfrtp_4 _26819_ (.CLK(clknet_leaf_48_clk_sys),
    .D(_00436_),
    .RESET_B(net676),
    .Q(\top0.svm0.state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _26820_ (.CLK(clknet_leaf_48_clk_sys),
    .D(_00437_),
    .RESET_B(net676),
    .Q(\top0.svm0.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26821_ (.CLK(clknet_leaf_36_clk_sys),
    .D(_00438_),
    .RESET_B(net676),
    .Q(\top0.svm0.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26822_ (.CLK(clknet_leaf_38_clk_sys),
    .D(net705),
    .RESET_B(net677),
    .Q(net4));
 sky130_fd_sc_hd__dfrtp_1 _26823_ (.CLK(clknet_leaf_37_clk_sys),
    .D(net709),
    .RESET_B(net679),
    .Q(net5));
 sky130_fd_sc_hd__dfrtp_1 _26824_ (.CLK(clknet_leaf_37_clk_sys),
    .D(net707),
    .RESET_B(net679),
    .Q(net6));
 sky130_fd_sc_hd__dfrtp_2 _26825_ (.CLK(clknet_leaf_46_clk_sys),
    .D(_00442_),
    .RESET_B(net680),
    .Q(\top0.svm0.counter[0] ));
 sky130_fd_sc_hd__dfrtp_4 _26826_ (.CLK(clknet_leaf_46_clk_sys),
    .D(_00443_),
    .RESET_B(net680),
    .Q(\top0.svm0.counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26827_ (.CLK(clknet_leaf_46_clk_sys),
    .D(_00444_),
    .RESET_B(net680),
    .Q(\top0.svm0.counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26828_ (.CLK(clknet_leaf_46_clk_sys),
    .D(_00445_),
    .RESET_B(net680),
    .Q(\top0.svm0.counter[3] ));
 sky130_fd_sc_hd__dfrtp_4 _26829_ (.CLK(clknet_leaf_46_clk_sys),
    .D(_00446_),
    .RESET_B(net680),
    .Q(\top0.svm0.counter[4] ));
 sky130_fd_sc_hd__dfrtp_4 _26830_ (.CLK(clknet_leaf_43_clk_sys),
    .D(_00447_),
    .RESET_B(net680),
    .Q(\top0.svm0.counter[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26831_ (.CLK(clknet_leaf_46_clk_sys),
    .D(_00448_),
    .RESET_B(net680),
    .Q(\top0.svm0.counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26832_ (.CLK(clknet_leaf_42_clk_sys),
    .D(_00449_),
    .RESET_B(net684),
    .Q(\top0.svm0.counter[7] ));
 sky130_fd_sc_hd__dfrtp_4 _26833_ (.CLK(clknet_leaf_42_clk_sys),
    .D(_00450_),
    .RESET_B(net684),
    .Q(\top0.svm0.counter[8] ));
 sky130_fd_sc_hd__dfrtp_4 _26834_ (.CLK(clknet_leaf_43_clk_sys),
    .D(_00451_),
    .RESET_B(net682),
    .Q(\top0.svm0.counter[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26835_ (.CLK(clknet_leaf_40_clk_sys),
    .D(_00452_),
    .RESET_B(net682),
    .Q(\top0.svm0.counter[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26836_ (.CLK(clknet_leaf_36_clk_sys),
    .D(_00453_),
    .RESET_B(net678),
    .Q(\top0.svm0.counter[11] ));
 sky130_fd_sc_hd__dfrtp_4 _26837_ (.CLK(clknet_leaf_36_clk_sys),
    .D(_00454_),
    .RESET_B(net676),
    .Q(\top0.svm0.counter[12] ));
 sky130_fd_sc_hd__dfrtp_4 _26838_ (.CLK(clknet_leaf_36_clk_sys),
    .D(_00455_),
    .RESET_B(net676),
    .Q(\top0.svm0.counter[13] ));
 sky130_fd_sc_hd__dfrtp_2 _26839_ (.CLK(clknet_leaf_47_clk_sys),
    .D(_00456_),
    .RESET_B(net680),
    .Q(\top0.svm0.counter[14] ));
 sky130_fd_sc_hd__dfrtp_4 _26840_ (.CLK(clknet_leaf_46_clk_sys),
    .D(_00457_),
    .RESET_B(net676),
    .Q(\top0.svm0.counter[15] ));
 sky130_fd_sc_hd__dfrtp_4 _26841_ (.CLK(clknet_leaf_45_clk_sys),
    .D(_00458_),
    .RESET_B(net681),
    .Q(\top0.svm0.delta[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26842_ (.CLK(clknet_leaf_44_clk_sys),
    .D(_00459_),
    .RESET_B(net681),
    .Q(\top0.svm0.delta[2] ));
 sky130_fd_sc_hd__dfrtp_4 _26843_ (.CLK(clknet_leaf_45_clk_sys),
    .D(_00460_),
    .RESET_B(net681),
    .Q(\top0.svm0.delta[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26844_ (.CLK(clknet_leaf_44_clk_sys),
    .D(_00461_),
    .RESET_B(net681),
    .Q(\top0.svm0.delta[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26845_ (.CLK(clknet_leaf_44_clk_sys),
    .D(_00462_),
    .RESET_B(net681),
    .Q(\top0.svm0.delta[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26846_ (.CLK(clknet_leaf_44_clk_sys),
    .D(_00463_),
    .RESET_B(net681),
    .Q(\top0.svm0.delta[6] ));
 sky130_fd_sc_hd__dfrtp_4 _26847_ (.CLK(clknet_leaf_43_clk_sys),
    .D(_00464_),
    .RESET_B(net681),
    .Q(\top0.svm0.delta[7] ));
 sky130_fd_sc_hd__dfrtp_4 _26848_ (.CLK(clknet_leaf_44_clk_sys),
    .D(_00465_),
    .RESET_B(net686),
    .Q(\top0.svm0.delta[8] ));
 sky130_fd_sc_hd__dfrtp_2 _26849_ (.CLK(clknet_leaf_44_clk_sys),
    .D(_00466_),
    .RESET_B(net686),
    .Q(\top0.svm0.delta[9] ));
 sky130_fd_sc_hd__dfrtp_4 _26850_ (.CLK(clknet_leaf_46_clk_sys),
    .D(_00467_),
    .RESET_B(net681),
    .Q(\top0.svm0.delta[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26851_ (.CLK(clknet_leaf_47_clk_sys),
    .D(_00468_),
    .RESET_B(net676),
    .Q(\top0.svm0.delta[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26852_ (.CLK(clknet_leaf_47_clk_sys),
    .D(_00469_),
    .RESET_B(net676),
    .Q(\top0.svm0.delta[12] ));
 sky130_fd_sc_hd__dfrtp_2 _26853_ (.CLK(clknet_leaf_47_clk_sys),
    .D(_00470_),
    .RESET_B(net676),
    .Q(\top0.svm0.delta[13] ));
 sky130_fd_sc_hd__dfrtp_4 _26854_ (.CLK(clknet_leaf_46_clk_sys),
    .D(_00471_),
    .RESET_B(net680),
    .Q(\top0.svm0.delta[14] ));
 sky130_fd_sc_hd__dfrtp_2 _26855_ (.CLK(clknet_leaf_46_clk_sys),
    .D(_00472_),
    .RESET_B(net680),
    .Q(\top0.svm0.delta[15] ));
 sky130_fd_sc_hd__dfstp_1 _26856_ (.CLK(clknet_leaf_36_clk_sys),
    .D(_00473_),
    .SET_B(net686),
    .Q(\top0.svm0.rising ));
 sky130_fd_sc_hd__dfrtp_1 _26857_ (.CLK(clknet_leaf_38_clk_sys),
    .D(_00474_),
    .RESET_B(net677),
    .Q(\top0.svm0.calc_ready ));
 sky130_fd_sc_hd__dfrtp_1 _26858_ (.CLK(clknet_leaf_40_clk_sys),
    .D(_00475_),
    .RESET_B(net678),
    .Q(\top0.svm0.tA[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26859_ (.CLK(clknet_leaf_36_clk_sys),
    .D(_00476_),
    .RESET_B(net678),
    .Q(\top0.svm0.tA[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26860_ (.CLK(clknet_leaf_36_clk_sys),
    .D(_00477_),
    .RESET_B(net678),
    .Q(\top0.svm0.tA[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26861_ (.CLK(clknet_leaf_40_clk_sys),
    .D(_00478_),
    .RESET_B(net682),
    .Q(\top0.svm0.tA[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26862_ (.CLK(clknet_leaf_40_clk_sys),
    .D(_00479_),
    .RESET_B(net682),
    .Q(\top0.svm0.tA[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26863_ (.CLK(clknet_leaf_41_clk_sys),
    .D(_00480_),
    .RESET_B(net683),
    .Q(\top0.svm0.tA[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26864_ (.CLK(clknet_leaf_41_clk_sys),
    .D(_00481_),
    .RESET_B(net683),
    .Q(\top0.svm0.tA[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26865_ (.CLK(clknet_leaf_41_clk_sys),
    .D(_00482_),
    .RESET_B(net683),
    .Q(\top0.svm0.tA[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26866_ (.CLK(clknet_leaf_41_clk_sys),
    .D(_00483_),
    .RESET_B(net683),
    .Q(\top0.svm0.tA[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26867_ (.CLK(clknet_leaf_39_clk_sys),
    .D(_00484_),
    .RESET_B(net683),
    .Q(\top0.svm0.tA[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26868_ (.CLK(clknet_leaf_40_clk_sys),
    .D(_00485_),
    .RESET_B(net677),
    .Q(\top0.svm0.tA[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26869_ (.CLK(clknet_leaf_40_clk_sys),
    .D(_00486_),
    .RESET_B(net678),
    .Q(\top0.svm0.tA[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26870_ (.CLK(clknet_leaf_36_clk_sys),
    .D(_00487_),
    .RESET_B(net678),
    .Q(\top0.svm0.tA[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26871_ (.CLK(clknet_leaf_37_clk_sys),
    .D(_00488_),
    .RESET_B(net678),
    .Q(\top0.svm0.tA[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26872_ (.CLK(clknet_leaf_37_clk_sys),
    .D(_00489_),
    .RESET_B(net679),
    .Q(\top0.svm0.tA[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26873_ (.CLK(clknet_leaf_37_clk_sys),
    .D(_00490_),
    .RESET_B(net679),
    .Q(\top0.svm0.tA[15] ));
 sky130_fd_sc_hd__dfrtp_1 _26874_ (.CLK(clknet_leaf_40_clk_sys),
    .D(_00491_),
    .RESET_B(net682),
    .Q(\top0.svm0.tB[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26875_ (.CLK(clknet_leaf_40_clk_sys),
    .D(_00492_),
    .RESET_B(net682),
    .Q(\top0.svm0.tB[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26876_ (.CLK(clknet_leaf_42_clk_sys),
    .D(_00493_),
    .RESET_B(net684),
    .Q(\top0.svm0.tB[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26877_ (.CLK(clknet_leaf_42_clk_sys),
    .D(_00494_),
    .RESET_B(net684),
    .Q(\top0.svm0.tB[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26878_ (.CLK(clknet_leaf_42_clk_sys),
    .D(_00495_),
    .RESET_B(net684),
    .Q(\top0.svm0.tB[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26879_ (.CLK(clknet_leaf_42_clk_sys),
    .D(_00496_),
    .RESET_B(net685),
    .Q(\top0.svm0.tB[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26880_ (.CLK(clknet_leaf_41_clk_sys),
    .D(_00497_),
    .RESET_B(net685),
    .Q(\top0.svm0.tB[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26881_ (.CLK(clknet_leaf_41_clk_sys),
    .D(_00498_),
    .RESET_B(net685),
    .Q(\top0.svm0.tB[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26882_ (.CLK(clknet_leaf_41_clk_sys),
    .D(_00499_),
    .RESET_B(net683),
    .Q(\top0.svm0.tB[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26883_ (.CLK(clknet_leaf_39_clk_sys),
    .D(_00500_),
    .RESET_B(net683),
    .Q(\top0.svm0.tB[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26884_ (.CLK(clknet_leaf_38_clk_sys),
    .D(_00501_),
    .RESET_B(net677),
    .Q(\top0.svm0.tB[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26885_ (.CLK(clknet_leaf_38_clk_sys),
    .D(_00502_),
    .RESET_B(net678),
    .Q(\top0.svm0.tB[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26886_ (.CLK(clknet_leaf_38_clk_sys),
    .D(_00503_),
    .RESET_B(net677),
    .Q(\top0.svm0.tB[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26887_ (.CLK(clknet_leaf_38_clk_sys),
    .D(_00504_),
    .RESET_B(net677),
    .Q(\top0.svm0.tB[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26888_ (.CLK(clknet_leaf_37_clk_sys),
    .D(_00505_),
    .RESET_B(net679),
    .Q(\top0.svm0.tB[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26889_ (.CLK(clknet_leaf_37_clk_sys),
    .D(_00506_),
    .RESET_B(net679),
    .Q(\top0.svm0.tB[15] ));
 sky130_fd_sc_hd__dfrtp_1 _26890_ (.CLK(clknet_leaf_105_clk_sys),
    .D(_00507_),
    .RESET_B(net577),
    .Q(\top0.cordic0.vec[1][0] ));
 sky130_fd_sc_hd__dfrtp_1 _26891_ (.CLK(clknet_leaf_105_clk_sys),
    .D(_00508_),
    .RESET_B(net577),
    .Q(\top0.cordic0.vec[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _26892_ (.CLK(clknet_leaf_105_clk_sys),
    .D(_00509_),
    .RESET_B(net577),
    .Q(\top0.cordic0.vec[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _26893_ (.CLK(clknet_leaf_107_clk_sys),
    .D(_00510_),
    .RESET_B(net577),
    .Q(\top0.cordic0.vec[1][3] ));
 sky130_fd_sc_hd__dfrtp_2 _26894_ (.CLK(clknet_leaf_106_clk_sys),
    .D(_00511_),
    .RESET_B(net577),
    .Q(\top0.cordic0.vec[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _26895_ (.CLK(clknet_leaf_106_clk_sys),
    .D(_00512_),
    .RESET_B(net577),
    .Q(\top0.cordic0.vec[1][5] ));
 sky130_fd_sc_hd__dfrtp_1 _26896_ (.CLK(clknet_leaf_106_clk_sys),
    .D(_00513_),
    .RESET_B(net577),
    .Q(\top0.cordic0.vec[1][6] ));
 sky130_fd_sc_hd__dfrtp_1 _26897_ (.CLK(clknet_leaf_107_clk_sys),
    .D(_00514_),
    .RESET_B(net577),
    .Q(\top0.cordic0.vec[1][7] ));
 sky130_fd_sc_hd__dfrtp_1 _26898_ (.CLK(clknet_leaf_107_clk_sys),
    .D(_00515_),
    .RESET_B(net577),
    .Q(\top0.cordic0.vec[1][8] ));
 sky130_fd_sc_hd__dfrtp_1 _26899_ (.CLK(clknet_leaf_108_clk_sys),
    .D(_00516_),
    .RESET_B(net581),
    .Q(\top0.cordic0.vec[1][9] ));
 sky130_fd_sc_hd__dfrtp_1 _26900_ (.CLK(clknet_leaf_108_clk_sys),
    .D(_00517_),
    .RESET_B(net585),
    .Q(\top0.cordic0.vec[1][10] ));
 sky130_fd_sc_hd__dfrtp_1 _26901_ (.CLK(clknet_leaf_108_clk_sys),
    .D(_00518_),
    .RESET_B(net585),
    .Q(\top0.cordic0.vec[1][11] ));
 sky130_fd_sc_hd__dfrtp_1 _26902_ (.CLK(clknet_leaf_4_clk_sys),
    .D(_00519_),
    .RESET_B(net585),
    .Q(\top0.cordic0.vec[1][12] ));
 sky130_fd_sc_hd__dfrtp_1 _26903_ (.CLK(clknet_leaf_4_clk_sys),
    .D(_00520_),
    .RESET_B(net580),
    .Q(\top0.cordic0.vec[1][13] ));
 sky130_fd_sc_hd__dfrtp_2 _26904_ (.CLK(clknet_leaf_4_clk_sys),
    .D(_00521_),
    .RESET_B(net580),
    .Q(\top0.cordic0.vec[1][14] ));
 sky130_fd_sc_hd__dfrtp_1 _26905_ (.CLK(clknet_leaf_4_clk_sys),
    .D(_00522_),
    .RESET_B(net580),
    .Q(\top0.cordic0.vec[1][15] ));
 sky130_fd_sc_hd__dfrtp_1 _26906_ (.CLK(clknet_leaf_5_clk_sys),
    .D(_00523_),
    .RESET_B(net581),
    .Q(\top0.cordic0.vec[1][16] ));
 sky130_fd_sc_hd__dfrtp_1 _26907_ (.CLK(clknet_leaf_5_clk_sys),
    .D(_00524_),
    .RESET_B(net590),
    .Q(\top0.cordic0.vec[1][17] ));
 sky130_fd_sc_hd__dfrtp_4 _26908_ (.CLK(clknet_leaf_109_clk_sys),
    .D(_00525_),
    .RESET_B(net579),
    .Q(\top0.matmul0.sin[0] ));
 sky130_fd_sc_hd__dfrtp_4 _26909_ (.CLK(clknet_leaf_110_clk_sys),
    .D(_00526_),
    .RESET_B(net579),
    .Q(\top0.matmul0.sin[1] ));
 sky130_fd_sc_hd__dfrtp_4 _26910_ (.CLK(clknet_leaf_110_clk_sys),
    .D(_00527_),
    .RESET_B(net579),
    .Q(\top0.matmul0.sin[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26911_ (.CLK(clknet_leaf_109_clk_sys),
    .D(_00528_),
    .RESET_B(net579),
    .Q(\top0.matmul0.sin[3] ));
 sky130_fd_sc_hd__dfrtp_4 _26912_ (.CLK(clknet_leaf_0_clk_sys),
    .D(_00529_),
    .RESET_B(net578),
    .Q(\top0.matmul0.sin[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26913_ (.CLK(clknet_leaf_2_clk_sys),
    .D(_00530_),
    .RESET_B(net582),
    .Q(\top0.matmul0.sin[5] ));
 sky130_fd_sc_hd__dfrtp_2 _26914_ (.CLK(clknet_leaf_1_clk_sys),
    .D(_00531_),
    .RESET_B(net582),
    .Q(\top0.matmul0.sin[6] ));
 sky130_fd_sc_hd__dfrtp_4 _26915_ (.CLK(clknet_leaf_7_clk_sys),
    .D(_00532_),
    .RESET_B(net583),
    .Q(\top0.matmul0.sin[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26916_ (.CLK(clknet_leaf_2_clk_sys),
    .D(_00533_),
    .RESET_B(net583),
    .Q(\top0.matmul0.sin[8] ));
 sky130_fd_sc_hd__dfrtp_2 _26917_ (.CLK(clknet_leaf_3_clk_sys),
    .D(_00534_),
    .RESET_B(net583),
    .Q(\top0.matmul0.sin[9] ));
 sky130_fd_sc_hd__dfrtp_4 _26918_ (.CLK(clknet_leaf_1_clk_sys),
    .D(_00535_),
    .RESET_B(net582),
    .Q(\top0.matmul0.sin[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26919_ (.CLK(clknet_leaf_1_clk_sys),
    .D(_00536_),
    .RESET_B(net582),
    .Q(\top0.matmul0.sin[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26920_ (.CLK(clknet_leaf_0_clk_sys),
    .D(_00537_),
    .RESET_B(net578),
    .Q(\top0.matmul0.sin[12] ));
 sky130_fd_sc_hd__dfrtp_4 _26921_ (.CLK(clknet_leaf_0_clk_sys),
    .D(_00538_),
    .RESET_B(net578),
    .Q(\top0.matmul0.sin[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26922_ (.CLK(clknet_leaf_3_clk_sys),
    .D(_00539_),
    .RESET_B(net581),
    .Q(\top0.matmul0.cos[0] ));
 sky130_fd_sc_hd__dfrtp_2 _26923_ (.CLK(clknet_leaf_4_clk_sys),
    .D(_00540_),
    .RESET_B(net581),
    .Q(\top0.matmul0.cos[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26924_ (.CLK(clknet_leaf_4_clk_sys),
    .D(_00541_),
    .RESET_B(net580),
    .Q(\top0.matmul0.cos[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26925_ (.CLK(clknet_leaf_5_clk_sys),
    .D(_00542_),
    .RESET_B(net598),
    .Q(\top0.matmul0.cos[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26926_ (.CLK(clknet_leaf_4_clk_sys),
    .D(_00543_),
    .RESET_B(net580),
    .Q(\top0.matmul0.cos[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26927_ (.CLK(clknet_leaf_7_clk_sys),
    .D(_00544_),
    .RESET_B(net593),
    .Q(\top0.matmul0.cos[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26928_ (.CLK(clknet_leaf_7_clk_sys),
    .D(_00545_),
    .RESET_B(net592),
    .Q(\top0.matmul0.cos[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26929_ (.CLK(clknet_leaf_7_clk_sys),
    .D(_00546_),
    .RESET_B(net593),
    .Q(\top0.matmul0.cos[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26930_ (.CLK(clknet_leaf_3_clk_sys),
    .D(_00547_),
    .RESET_B(net583),
    .Q(\top0.matmul0.cos[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26931_ (.CLK(clknet_leaf_7_clk_sys),
    .D(_00548_),
    .RESET_B(net592),
    .Q(\top0.matmul0.cos[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26932_ (.CLK(clknet_leaf_7_clk_sys),
    .D(_00549_),
    .RESET_B(net593),
    .Q(\top0.matmul0.cos[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26933_ (.CLK(clknet_leaf_3_clk_sys),
    .D(_00550_),
    .RESET_B(net583),
    .Q(\top0.matmul0.cos[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26934_ (.CLK(clknet_leaf_7_clk_sys),
    .D(_00551_),
    .RESET_B(net593),
    .Q(\top0.matmul0.cos[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26935_ (.CLK(clknet_leaf_3_clk_sys),
    .D(_00552_),
    .RESET_B(net583),
    .Q(\top0.matmul0.cos[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26936_ (.CLK(clknet_leaf_8_clk_sys),
    .D(_00553_),
    .RESET_B(net595),
    .Q(\top0.matmul0.a[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26937_ (.CLK(clknet_leaf_9_clk_sys),
    .D(_00554_),
    .RESET_B(net595),
    .Q(\top0.matmul0.a[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26938_ (.CLK(clknet_leaf_9_clk_sys),
    .D(_00555_),
    .RESET_B(net595),
    .Q(\top0.matmul0.a[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26939_ (.CLK(clknet_leaf_8_clk_sys),
    .D(_00556_),
    .RESET_B(net595),
    .Q(\top0.matmul0.a[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26940_ (.CLK(clknet_leaf_9_clk_sys),
    .D(_00557_),
    .RESET_B(net594),
    .Q(\top0.matmul0.a[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26941_ (.CLK(clknet_leaf_9_clk_sys),
    .D(_00558_),
    .RESET_B(net594),
    .Q(\top0.matmul0.a[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26942_ (.CLK(clknet_leaf_6_clk_sys),
    .D(_00559_),
    .RESET_B(net594),
    .Q(\top0.matmul0.a[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26943_ (.CLK(clknet_leaf_9_clk_sys),
    .D(_00560_),
    .RESET_B(net594),
    .Q(\top0.matmul0.a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26944_ (.CLK(clknet_leaf_6_clk_sys),
    .D(_00561_),
    .RESET_B(net594),
    .Q(\top0.matmul0.a[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26945_ (.CLK(clknet_leaf_8_clk_sys),
    .D(_00562_),
    .RESET_B(net595),
    .Q(\top0.matmul0.a[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26946_ (.CLK(clknet_leaf_9_clk_sys),
    .D(_00563_),
    .RESET_B(net595),
    .Q(\top0.matmul0.a[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26947_ (.CLK(clknet_leaf_13_clk_sys),
    .D(_00564_),
    .RESET_B(net595),
    .Q(\top0.matmul0.a[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26948_ (.CLK(clknet_leaf_9_clk_sys),
    .D(_00565_),
    .RESET_B(net595),
    .Q(\top0.matmul0.a[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26949_ (.CLK(clknet_leaf_9_clk_sys),
    .D(_00566_),
    .RESET_B(net596),
    .Q(\top0.matmul0.a[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26950_ (.CLK(clknet_leaf_13_clk_sys),
    .D(_00567_),
    .RESET_B(net616),
    .Q(\top0.matmul0.a[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26951_ (.CLK(clknet_leaf_9_clk_sys),
    .D(_00568_),
    .RESET_B(net596),
    .Q(\top0.matmul0.a[15] ));
 sky130_fd_sc_hd__dfrtp_1 _26952_ (.CLK(clknet_leaf_16_clk_sys),
    .D(_00569_),
    .RESET_B(net613),
    .Q(\top0.matmul0.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26953_ (.CLK(clknet_leaf_16_clk_sys),
    .D(_00570_),
    .RESET_B(net613),
    .Q(\top0.matmul0.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _26954_ (.CLK(clknet_leaf_16_clk_sys),
    .D(_00571_),
    .RESET_B(net613),
    .Q(\top0.matmul0.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _26955_ (.CLK(clknet_leaf_13_clk_sys),
    .D(_00572_),
    .RESET_B(net613),
    .Q(\top0.matmul0.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26956_ (.CLK(clknet_leaf_13_clk_sys),
    .D(_00573_),
    .RESET_B(net616),
    .Q(\top0.matmul0.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26957_ (.CLK(clknet_leaf_13_clk_sys),
    .D(_00574_),
    .RESET_B(net616),
    .Q(\top0.matmul0.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26958_ (.CLK(clknet_leaf_13_clk_sys),
    .D(_00575_),
    .RESET_B(net616),
    .Q(\top0.matmul0.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26959_ (.CLK(clknet_leaf_15_clk_sys),
    .D(_00576_),
    .RESET_B(net613),
    .Q(\top0.matmul0.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26960_ (.CLK(clknet_leaf_14_clk_sys),
    .D(_00577_),
    .RESET_B(net617),
    .Q(\top0.matmul0.b[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26961_ (.CLK(clknet_leaf_31_clk_sys),
    .D(_00578_),
    .RESET_B(net617),
    .Q(\top0.matmul0.b[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26962_ (.CLK(clknet_leaf_14_clk_sys),
    .D(_00579_),
    .RESET_B(net617),
    .Q(\top0.matmul0.b[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26963_ (.CLK(clknet_leaf_14_clk_sys),
    .D(_00580_),
    .RESET_B(net617),
    .Q(\top0.matmul0.b[11] ));
 sky130_fd_sc_hd__dfrtp_1 _26964_ (.CLK(clknet_leaf_31_clk_sys),
    .D(_00581_),
    .RESET_B(net617),
    .Q(\top0.matmul0.b[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26965_ (.CLK(clknet_leaf_31_clk_sys),
    .D(_00582_),
    .RESET_B(net621),
    .Q(\top0.matmul0.b[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26966_ (.CLK(clknet_leaf_30_clk_sys),
    .D(_00583_),
    .RESET_B(net621),
    .Q(\top0.matmul0.b[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26967_ (.CLK(clknet_leaf_15_clk_sys),
    .D(_00584_),
    .RESET_B(net613),
    .Q(\top0.matmul0.b[15] ));
 sky130_fd_sc_hd__dfrtp_4 _26968_ (.CLK(clknet_leaf_30_clk_sys),
    .D(_00585_),
    .RESET_B(net623),
    .Q(\top0.matmul0.alpha_pass[0] ));
 sky130_fd_sc_hd__dfrtp_4 _26969_ (.CLK(clknet_leaf_30_clk_sys),
    .D(_00586_),
    .RESET_B(net623),
    .Q(\top0.matmul0.alpha_pass[1] ));
 sky130_fd_sc_hd__dfrtp_4 _26970_ (.CLK(clknet_leaf_29_clk_sys),
    .D(_00587_),
    .RESET_B(net623),
    .Q(\top0.matmul0.alpha_pass[2] ));
 sky130_fd_sc_hd__dfrtp_4 _26971_ (.CLK(clknet_leaf_27_clk_sys),
    .D(_00588_),
    .RESET_B(net621),
    .Q(\top0.matmul0.alpha_pass[3] ));
 sky130_fd_sc_hd__dfrtp_4 _26972_ (.CLK(clknet_leaf_29_clk_sys),
    .D(_00589_),
    .RESET_B(net624),
    .Q(\top0.matmul0.alpha_pass[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26973_ (.CLK(clknet_leaf_28_clk_sys),
    .D(_00590_),
    .RESET_B(net622),
    .Q(\top0.matmul0.alpha_pass[5] ));
 sky130_fd_sc_hd__dfrtp_4 _26974_ (.CLK(clknet_leaf_28_clk_sys),
    .D(_00591_),
    .RESET_B(net624),
    .Q(\top0.matmul0.alpha_pass[6] ));
 sky130_fd_sc_hd__dfrtp_4 _26975_ (.CLK(clknet_leaf_28_clk_sys),
    .D(_00592_),
    .RESET_B(net622),
    .Q(\top0.matmul0.alpha_pass[7] ));
 sky130_fd_sc_hd__dfrtp_4 _26976_ (.CLK(clknet_leaf_28_clk_sys),
    .D(_00593_),
    .RESET_B(net622),
    .Q(\top0.matmul0.alpha_pass[8] ));
 sky130_fd_sc_hd__dfrtp_4 _26977_ (.CLK(clknet_leaf_25_clk_sys),
    .D(_00594_),
    .RESET_B(net627),
    .Q(\top0.matmul0.alpha_pass[9] ));
 sky130_fd_sc_hd__dfrtp_4 _26978_ (.CLK(clknet_leaf_25_clk_sys),
    .D(_00595_),
    .RESET_B(net628),
    .Q(\top0.matmul0.alpha_pass[10] ));
 sky130_fd_sc_hd__dfrtp_4 _26979_ (.CLK(clknet_leaf_29_clk_sys),
    .D(_00596_),
    .RESET_B(net624),
    .Q(\top0.matmul0.alpha_pass[11] ));
 sky130_fd_sc_hd__dfrtp_4 _26980_ (.CLK(clknet_leaf_25_clk_sys),
    .D(_00597_),
    .RESET_B(net628),
    .Q(\top0.matmul0.alpha_pass[12] ));
 sky130_fd_sc_hd__dfrtp_4 _26981_ (.CLK(clknet_leaf_31_clk_sys),
    .D(_00598_),
    .RESET_B(net619),
    .Q(\top0.matmul0.alpha_pass[13] ));
 sky130_fd_sc_hd__dfrtp_4 _26982_ (.CLK(clknet_leaf_25_clk_sys),
    .D(_00599_),
    .RESET_B(net627),
    .Q(\top0.matmul0.alpha_pass[14] ));
 sky130_fd_sc_hd__dfrtp_4 _26983_ (.CLK(clknet_leaf_25_clk_sys),
    .D(_00600_),
    .RESET_B(net628),
    .Q(\top0.matmul0.alpha_pass[15] ));
 sky130_fd_sc_hd__dfrtp_2 _26984_ (.CLK(clknet_leaf_30_clk_sys),
    .D(_00601_),
    .RESET_B(net621),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _26985_ (.CLK(clknet_leaf_27_clk_sys),
    .D(_00602_),
    .RESET_B(net621),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[1] ));
 sky130_fd_sc_hd__dfrtp_2 _26986_ (.CLK(clknet_leaf_27_clk_sys),
    .D(_00603_),
    .RESET_B(net621),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[2] ));
 sky130_fd_sc_hd__dfrtp_2 _26987_ (.CLK(clknet_leaf_27_clk_sys),
    .D(_00604_),
    .RESET_B(net615),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _26988_ (.CLK(clknet_leaf_28_clk_sys),
    .D(_00605_),
    .RESET_B(net622),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _26989_ (.CLK(clknet_leaf_28_clk_sys),
    .D(_00606_),
    .RESET_B(net622),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _26990_ (.CLK(clknet_leaf_25_clk_sys),
    .D(_00607_),
    .RESET_B(net627),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _26991_ (.CLK(clknet_leaf_26_clk_sys),
    .D(_00608_),
    .RESET_B(net625),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _26992_ (.CLK(clknet_leaf_26_clk_sys),
    .D(_00609_),
    .RESET_B(net627),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _26993_ (.CLK(clknet_leaf_26_clk_sys),
    .D(_00610_),
    .RESET_B(net625),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _26994_ (.CLK(clknet_leaf_23_clk_sys),
    .D(_00611_),
    .RESET_B(net625),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _26995_ (.CLK(clknet_leaf_23_clk_sys),
    .D(_00612_),
    .RESET_B(net625),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[11] ));
 sky130_fd_sc_hd__dfrtp_2 _26996_ (.CLK(clknet_leaf_24_clk_sys),
    .D(_00613_),
    .RESET_B(net625),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[12] ));
 sky130_fd_sc_hd__dfrtp_1 _26997_ (.CLK(clknet_leaf_24_clk_sys),
    .D(_00614_),
    .RESET_B(net625),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _26998_ (.CLK(clknet_leaf_23_clk_sys),
    .D(_00615_),
    .RESET_B(net625),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _26999_ (.CLK(clknet_leaf_24_clk_sys),
    .D(_00616_),
    .RESET_B(net626),
    .Q(\top0.matmul0.matmul_stage_inst.mult2[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27000_ (.CLK(clknet_leaf_27_clk_sys),
    .D(_00617_),
    .RESET_B(net615),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _27001_ (.CLK(clknet_leaf_27_clk_sys),
    .D(_00618_),
    .RESET_B(net615),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _27002_ (.CLK(clknet_leaf_27_clk_sys),
    .D(_00619_),
    .RESET_B(net615),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _27003_ (.CLK(clknet_leaf_28_clk_sys),
    .D(_00620_),
    .RESET_B(net622),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _27004_ (.CLK(clknet_leaf_28_clk_sys),
    .D(_00621_),
    .RESET_B(net622),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _27005_ (.CLK(clknet_leaf_25_clk_sys),
    .D(_00622_),
    .RESET_B(net627),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _27006_ (.CLK(clknet_leaf_25_clk_sys),
    .D(_00623_),
    .RESET_B(net627),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _27007_ (.CLK(clknet_leaf_26_clk_sys),
    .D(_00624_),
    .RESET_B(net627),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _27008_ (.CLK(clknet_leaf_26_clk_sys),
    .D(_00625_),
    .RESET_B(net625),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _27009_ (.CLK(clknet_leaf_23_clk_sys),
    .D(_00626_),
    .RESET_B(net625),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _27010_ (.CLK(clknet_leaf_23_clk_sys),
    .D(_00627_),
    .RESET_B(net625),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _27011_ (.CLK(clknet_leaf_23_clk_sys),
    .D(_00628_),
    .RESET_B(net626),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _27012_ (.CLK(clknet_leaf_23_clk_sys),
    .D(_00629_),
    .RESET_B(net626),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _27013_ (.CLK(clknet_leaf_24_clk_sys),
    .D(_00630_),
    .RESET_B(net626),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _27014_ (.CLK(clknet_leaf_24_clk_sys),
    .D(_00631_),
    .RESET_B(net626),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _27015_ (.CLK(clknet_leaf_24_clk_sys),
    .D(_00632_),
    .RESET_B(net626),
    .Q(\top0.matmul0.matmul_stage_inst.mult1[15] ));
 sky130_fd_sc_hd__dfrtp_2 _27016_ (.CLK(clknet_leaf_16_clk_sys),
    .D(_00633_),
    .RESET_B(net613),
    .Q(\top0.matmul0.matmul_stage_inst.f[0] ));
 sky130_fd_sc_hd__dfrtp_1 _27017_ (.CLK(clknet_leaf_16_clk_sys),
    .D(_00634_),
    .RESET_B(net611),
    .Q(\top0.matmul0.matmul_stage_inst.f[1] ));
 sky130_fd_sc_hd__dfrtp_4 _27018_ (.CLK(clknet_leaf_16_clk_sys),
    .D(_00635_),
    .RESET_B(net613),
    .Q(\top0.matmul0.matmul_stage_inst.f[2] ));
 sky130_fd_sc_hd__dfrtp_1 _27019_ (.CLK(clknet_leaf_17_clk_sys),
    .D(_00636_),
    .RESET_B(net611),
    .Q(\top0.matmul0.matmul_stage_inst.f[3] ));
 sky130_fd_sc_hd__dfrtp_1 _27020_ (.CLK(clknet_leaf_16_clk_sys),
    .D(_00637_),
    .RESET_B(net612),
    .Q(\top0.matmul0.matmul_stage_inst.f[4] ));
 sky130_fd_sc_hd__dfrtp_1 _27021_ (.CLK(clknet_leaf_18_clk_sys),
    .D(_00638_),
    .RESET_B(net614),
    .Q(\top0.matmul0.matmul_stage_inst.f[5] ));
 sky130_fd_sc_hd__dfrtp_1 _27022_ (.CLK(clknet_leaf_16_clk_sys),
    .D(_00639_),
    .RESET_B(net612),
    .Q(\top0.matmul0.matmul_stage_inst.f[6] ));
 sky130_fd_sc_hd__dfrtp_1 _27023_ (.CLK(clknet_leaf_15_clk_sys),
    .D(_00640_),
    .RESET_B(net614),
    .Q(\top0.matmul0.matmul_stage_inst.f[7] ));
 sky130_fd_sc_hd__dfrtp_1 _27024_ (.CLK(clknet_leaf_18_clk_sys),
    .D(_00641_),
    .RESET_B(net612),
    .Q(\top0.matmul0.matmul_stage_inst.f[8] ));
 sky130_fd_sc_hd__dfrtp_1 _27025_ (.CLK(clknet_leaf_15_clk_sys),
    .D(_00642_),
    .RESET_B(net617),
    .Q(\top0.matmul0.matmul_stage_inst.f[9] ));
 sky130_fd_sc_hd__dfrtp_1 _27026_ (.CLK(clknet_leaf_15_clk_sys),
    .D(_00643_),
    .RESET_B(net617),
    .Q(\top0.matmul0.matmul_stage_inst.f[10] ));
 sky130_fd_sc_hd__dfrtp_1 _27027_ (.CLK(clknet_leaf_15_clk_sys),
    .D(_00644_),
    .RESET_B(net614),
    .Q(\top0.matmul0.matmul_stage_inst.f[11] ));
 sky130_fd_sc_hd__dfrtp_1 _27028_ (.CLK(clknet_leaf_18_clk_sys),
    .D(_00645_),
    .RESET_B(net614),
    .Q(\top0.matmul0.matmul_stage_inst.f[12] ));
 sky130_fd_sc_hd__dfrtp_1 _27029_ (.CLK(clknet_3_3__leaf_clk_sys),
    .D(_00646_),
    .RESET_B(net615),
    .Q(\top0.matmul0.matmul_stage_inst.f[13] ));
 sky130_fd_sc_hd__dfrtp_1 _27030_ (.CLK(clknet_leaf_27_clk_sys),
    .D(_00647_),
    .RESET_B(net621),
    .Q(\top0.matmul0.matmul_stage_inst.f[14] ));
 sky130_fd_sc_hd__dfrtp_1 _27031_ (.CLK(clknet_leaf_15_clk_sys),
    .D(_00648_),
    .RESET_B(net614),
    .Q(\top0.matmul0.matmul_stage_inst.f[15] ));
 sky130_fd_sc_hd__dfrtp_4 _27032_ (.CLK(clknet_leaf_15_clk_sys),
    .D(_00649_),
    .RESET_B(net613),
    .Q(\top0.matmul0.matmul_stage_inst.e[0] ));
 sky130_fd_sc_hd__dfrtp_1 _27033_ (.CLK(clknet_leaf_18_clk_sys),
    .D(_00650_),
    .RESET_B(net614),
    .Q(\top0.matmul0.matmul_stage_inst.e[1] ));
 sky130_fd_sc_hd__dfrtp_4 _27034_ (.CLK(clknet_leaf_15_clk_sys),
    .D(_00651_),
    .RESET_B(net614),
    .Q(\top0.matmul0.matmul_stage_inst.e[2] ));
 sky130_fd_sc_hd__dfrtp_1 _27035_ (.CLK(clknet_leaf_8_clk_sys),
    .D(_00652_),
    .RESET_B(net595),
    .Q(\top0.matmul0.matmul_stage_inst.e[3] ));
 sky130_fd_sc_hd__dfrtp_2 _27036_ (.CLK(clknet_leaf_9_clk_sys),
    .D(_00653_),
    .RESET_B(net594),
    .Q(\top0.matmul0.matmul_stage_inst.e[4] ));
 sky130_fd_sc_hd__dfrtp_2 _27037_ (.CLK(clknet_leaf_8_clk_sys),
    .D(_00654_),
    .RESET_B(net592),
    .Q(\top0.matmul0.matmul_stage_inst.e[5] ));
 sky130_fd_sc_hd__dfrtp_2 _27038_ (.CLK(clknet_leaf_7_clk_sys),
    .D(_00655_),
    .RESET_B(net593),
    .Q(\top0.matmul0.matmul_stage_inst.e[6] ));
 sky130_fd_sc_hd__dfrtp_1 _27039_ (.CLK(clknet_leaf_7_clk_sys),
    .D(_00656_),
    .RESET_B(net592),
    .Q(\top0.matmul0.matmul_stage_inst.e[7] ));
 sky130_fd_sc_hd__dfrtp_1 _27040_ (.CLK(clknet_leaf_7_clk_sys),
    .D(_00657_),
    .RESET_B(net593),
    .Q(\top0.matmul0.matmul_stage_inst.e[8] ));
 sky130_fd_sc_hd__dfrtp_1 _27041_ (.CLK(clknet_leaf_8_clk_sys),
    .D(_00658_),
    .RESET_B(net597),
    .Q(\top0.matmul0.matmul_stage_inst.e[9] ));
 sky130_fd_sc_hd__dfrtp_1 _27042_ (.CLK(clknet_leaf_8_clk_sys),
    .D(_00659_),
    .RESET_B(net597),
    .Q(\top0.matmul0.matmul_stage_inst.e[10] ));
 sky130_fd_sc_hd__dfrtp_1 _27043_ (.CLK(clknet_leaf_16_clk_sys),
    .D(_00660_),
    .RESET_B(net612),
    .Q(\top0.matmul0.matmul_stage_inst.e[11] ));
 sky130_fd_sc_hd__dfrtp_1 _27044_ (.CLK(clknet_leaf_16_clk_sys),
    .D(_00661_),
    .RESET_B(net613),
    .Q(\top0.matmul0.matmul_stage_inst.e[12] ));
 sky130_fd_sc_hd__dfrtp_1 _27045_ (.CLK(clknet_leaf_8_clk_sys),
    .D(_00662_),
    .RESET_B(net592),
    .Q(\top0.matmul0.matmul_stage_inst.e[13] ));
 sky130_fd_sc_hd__dfrtp_1 _27046_ (.CLK(clknet_leaf_16_clk_sys),
    .D(_00663_),
    .RESET_B(net612),
    .Q(\top0.matmul0.matmul_stage_inst.e[14] ));
 sky130_fd_sc_hd__dfrtp_1 _27047_ (.CLK(clknet_leaf_8_clk_sys),
    .D(_00664_),
    .RESET_B(net592),
    .Q(\top0.matmul0.matmul_stage_inst.e[15] ));
 sky130_fd_sc_hd__dfrtp_1 _27048_ (.CLK(clknet_leaf_17_clk_sys),
    .D(_00665_),
    .RESET_B(net611),
    .Q(\top0.matmul0.matmul_stage_inst.d[0] ));
 sky130_fd_sc_hd__dfrtp_1 _27049_ (.CLK(clknet_leaf_22_clk_sys),
    .D(_00666_),
    .RESET_B(net607),
    .Q(\top0.matmul0.matmul_stage_inst.d[1] ));
 sky130_fd_sc_hd__dfrtp_1 _27050_ (.CLK(clknet_leaf_22_clk_sys),
    .D(_00667_),
    .RESET_B(net607),
    .Q(\top0.matmul0.matmul_stage_inst.d[2] ));
 sky130_fd_sc_hd__dfrtp_1 _27051_ (.CLK(clknet_leaf_22_clk_sys),
    .D(_00668_),
    .RESET_B(net607),
    .Q(\top0.matmul0.matmul_stage_inst.d[4] ));
 sky130_fd_sc_hd__dfrtp_1 _27052_ (.CLK(clknet_leaf_20_clk_sys),
    .D(_00669_),
    .RESET_B(net611),
    .Q(\top0.matmul0.matmul_stage_inst.d[5] ));
 sky130_fd_sc_hd__dfrtp_1 _27053_ (.CLK(clknet_leaf_20_clk_sys),
    .D(_00670_),
    .RESET_B(net609),
    .Q(\top0.matmul0.matmul_stage_inst.d[6] ));
 sky130_fd_sc_hd__dfrtp_1 _27054_ (.CLK(clknet_leaf_17_clk_sys),
    .D(_00671_),
    .RESET_B(net609),
    .Q(\top0.matmul0.matmul_stage_inst.d[7] ));
 sky130_fd_sc_hd__dfrtp_1 _27055_ (.CLK(clknet_leaf_20_clk_sys),
    .D(_00672_),
    .RESET_B(net609),
    .Q(\top0.matmul0.matmul_stage_inst.d[8] ));
 sky130_fd_sc_hd__dfrtp_1 _27056_ (.CLK(clknet_leaf_20_clk_sys),
    .D(_00673_),
    .RESET_B(net609),
    .Q(\top0.matmul0.matmul_stage_inst.d[9] ));
 sky130_fd_sc_hd__dfrtp_1 _27057_ (.CLK(clknet_leaf_20_clk_sys),
    .D(_00674_),
    .RESET_B(net609),
    .Q(\top0.matmul0.matmul_stage_inst.d[10] ));
 sky130_fd_sc_hd__dfrtp_1 _27058_ (.CLK(clknet_leaf_20_clk_sys),
    .D(_00675_),
    .RESET_B(net610),
    .Q(\top0.matmul0.matmul_stage_inst.d[11] ));
 sky130_fd_sc_hd__dfrtp_1 _27059_ (.CLK(clknet_leaf_21_clk_sys),
    .D(_00676_),
    .RESET_B(net610),
    .Q(\top0.matmul0.matmul_stage_inst.d[12] ));
 sky130_fd_sc_hd__dfrtp_1 _27060_ (.CLK(clknet_leaf_21_clk_sys),
    .D(_00677_),
    .RESET_B(net610),
    .Q(\top0.matmul0.matmul_stage_inst.d[13] ));
 sky130_fd_sc_hd__dfrtp_1 _27061_ (.CLK(clknet_leaf_21_clk_sys),
    .D(_00678_),
    .RESET_B(net610),
    .Q(\top0.matmul0.matmul_stage_inst.a[14] ));
 sky130_fd_sc_hd__dfrtp_1 _27062_ (.CLK(clknet_leaf_110_clk_sys),
    .D(_00679_),
    .RESET_B(net578),
    .Q(\top0.matmul0.matmul_stage_inst.c[1] ));
 sky130_fd_sc_hd__dfrtp_1 _27063_ (.CLK(clknet_leaf_110_clk_sys),
    .D(_00680_),
    .RESET_B(net578),
    .Q(\top0.matmul0.matmul_stage_inst.c[2] ));
 sky130_fd_sc_hd__dfrtp_1 _27064_ (.CLK(clknet_leaf_110_clk_sys),
    .D(_00681_),
    .RESET_B(net578),
    .Q(\top0.matmul0.matmul_stage_inst.c[3] ));
 sky130_fd_sc_hd__dfrtp_1 _27065_ (.CLK(clknet_leaf_0_clk_sys),
    .D(_00682_),
    .RESET_B(net586),
    .Q(\top0.matmul0.matmul_stage_inst.c[4] ));
 sky130_fd_sc_hd__dfrtp_1 _27066_ (.CLK(clknet_leaf_8_clk_sys),
    .D(_00683_),
    .RESET_B(net592),
    .Q(\top0.matmul0.matmul_stage_inst.c[5] ));
 sky130_fd_sc_hd__dfrtp_1 _27067_ (.CLK(clknet_leaf_2_clk_sys),
    .D(_00684_),
    .RESET_B(net582),
    .Q(\top0.matmul0.matmul_stage_inst.c[6] ));
 sky130_fd_sc_hd__dfrtp_1 _27068_ (.CLK(clknet_leaf_2_clk_sys),
    .D(_00685_),
    .RESET_B(net583),
    .Q(\top0.matmul0.matmul_stage_inst.c[7] ));
 sky130_fd_sc_hd__dfrtp_1 _27069_ (.CLK(clknet_leaf_2_clk_sys),
    .D(_00686_),
    .RESET_B(net584),
    .Q(\top0.matmul0.matmul_stage_inst.c[8] ));
 sky130_fd_sc_hd__dfrtp_1 _27070_ (.CLK(clknet_leaf_2_clk_sys),
    .D(_00687_),
    .RESET_B(net584),
    .Q(\top0.matmul0.matmul_stage_inst.c[9] ));
 sky130_fd_sc_hd__dfrtp_1 _27071_ (.CLK(clknet_leaf_2_clk_sys),
    .D(_00688_),
    .RESET_B(net582),
    .Q(\top0.matmul0.matmul_stage_inst.c[10] ));
 sky130_fd_sc_hd__dfrtp_1 _27072_ (.CLK(clknet_leaf_2_clk_sys),
    .D(_00689_),
    .RESET_B(net582),
    .Q(\top0.matmul0.matmul_stage_inst.c[11] ));
 sky130_fd_sc_hd__dfrtp_1 _27073_ (.CLK(clknet_leaf_21_clk_sys),
    .D(_00690_),
    .RESET_B(net610),
    .Q(\top0.matmul0.matmul_stage_inst.c[12] ));
 sky130_fd_sc_hd__dfrtp_1 _27074_ (.CLK(clknet_leaf_21_clk_sys),
    .D(_00691_),
    .RESET_B(net607),
    .Q(\top0.matmul0.matmul_stage_inst.c[13] ));
 sky130_fd_sc_hd__dfrtp_1 _27075_ (.CLK(clknet_leaf_22_clk_sys),
    .D(_00692_),
    .RESET_B(net607),
    .Q(\top0.matmul0.matmul_stage_inst.c[14] ));
 sky130_fd_sc_hd__dfrtp_1 _27076_ (.CLK(clknet_leaf_22_clk_sys),
    .D(_00693_),
    .RESET_B(net607),
    .Q(\top0.matmul0.matmul_stage_inst.c[15] ));
 sky130_fd_sc_hd__dfrtp_1 _27077_ (.CLK(clknet_leaf_22_clk_sys),
    .D(_00694_),
    .RESET_B(net607),
    .Q(\top0.matmul0.matmul_stage_inst.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _27078_ (.CLK(clknet_leaf_110_clk_sys),
    .D(_00695_),
    .RESET_B(net579),
    .Q(\top0.matmul0.matmul_stage_inst.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _27079_ (.CLK(clknet_leaf_22_clk_sys),
    .D(_00696_),
    .RESET_B(net607),
    .Q(\top0.matmul0.matmul_stage_inst.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _27080_ (.CLK(clknet_leaf_22_clk_sys),
    .D(_00697_),
    .RESET_B(net607),
    .Q(\top0.matmul0.matmul_stage_inst.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _27081_ (.CLK(clknet_leaf_0_clk_sys),
    .D(_00698_),
    .RESET_B(net586),
    .Q(\top0.matmul0.matmul_stage_inst.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _27082_ (.CLK(clknet_leaf_20_clk_sys),
    .D(_00699_),
    .RESET_B(net609),
    .Q(\top0.matmul0.matmul_stage_inst.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _27083_ (.CLK(clknet_leaf_20_clk_sys),
    .D(_00700_),
    .RESET_B(net609),
    .Q(\top0.matmul0.matmul_stage_inst.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _27084_ (.CLK(clknet_leaf_8_clk_sys),
    .D(_00701_),
    .RESET_B(net592),
    .Q(\top0.matmul0.matmul_stage_inst.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _27085_ (.CLK(clknet_leaf_8_clk_sys),
    .D(_00702_),
    .RESET_B(net592),
    .Q(\top0.matmul0.matmul_stage_inst.b[8] ));
 sky130_fd_sc_hd__dfrtp_1 _27086_ (.CLK(clknet_leaf_8_clk_sys),
    .D(_00703_),
    .RESET_B(net584),
    .Q(\top0.matmul0.matmul_stage_inst.b[9] ));
 sky130_fd_sc_hd__dfrtp_1 _27087_ (.CLK(clknet_leaf_2_clk_sys),
    .D(_00704_),
    .RESET_B(net610),
    .Q(\top0.matmul0.matmul_stage_inst.b[10] ));
 sky130_fd_sc_hd__dfrtp_1 _27088_ (.CLK(clknet_leaf_1_clk_sys),
    .D(_00705_),
    .RESET_B(net584),
    .Q(\top0.matmul0.matmul_stage_inst.b[11] ));
 sky130_fd_sc_hd__dfrtp_1 _27089_ (.CLK(clknet_leaf_1_clk_sys),
    .D(_00706_),
    .RESET_B(net584),
    .Q(\top0.matmul0.matmul_stage_inst.b[12] ));
 sky130_fd_sc_hd__dfrtp_1 _27090_ (.CLK(clknet_leaf_1_clk_sys),
    .D(_00707_),
    .RESET_B(net584),
    .Q(\top0.matmul0.matmul_stage_inst.b[13] ));
 sky130_fd_sc_hd__dfrtp_1 _27091_ (.CLK(clknet_leaf_22_clk_sys),
    .D(_00708_),
    .RESET_B(net607),
    .Q(\top0.matmul0.matmul_stage_inst.b[14] ));
 sky130_fd_sc_hd__dfrtp_1 _27092_ (.CLK(clknet_leaf_22_clk_sys),
    .D(_00709_),
    .RESET_B(net608),
    .Q(\top0.matmul0.matmul_stage_inst.b[15] ));
 sky130_fd_sc_hd__dfrtp_1 _27093_ (.CLK(clknet_leaf_17_clk_sys),
    .D(_00710_),
    .RESET_B(net611),
    .Q(\top0.matmul0.matmul_stage_inst.a[0] ));
 sky130_fd_sc_hd__dfrtp_1 _27094_ (.CLK(clknet_leaf_22_clk_sys),
    .D(_00711_),
    .RESET_B(net608),
    .Q(\top0.matmul0.matmul_stage_inst.a[1] ));
 sky130_fd_sc_hd__dfrtp_1 _27095_ (.CLK(clknet_leaf_22_clk_sys),
    .D(_00712_),
    .RESET_B(net608),
    .Q(\top0.matmul0.matmul_stage_inst.a[2] ));
 sky130_fd_sc_hd__dfrtp_1 _27096_ (.CLK(clknet_leaf_17_clk_sys),
    .D(_00713_),
    .RESET_B(net611),
    .Q(\top0.matmul0.matmul_stage_inst.a[3] ));
 sky130_fd_sc_hd__dfrtp_1 _27097_ (.CLK(clknet_leaf_0_clk_sys),
    .D(_00714_),
    .RESET_B(net586),
    .Q(\top0.matmul0.matmul_stage_inst.a[4] ));
 sky130_fd_sc_hd__dfrtp_1 _27098_ (.CLK(clknet_leaf_20_clk_sys),
    .D(_00715_),
    .RESET_B(net609),
    .Q(\top0.matmul0.matmul_stage_inst.a[5] ));
 sky130_fd_sc_hd__dfrtp_1 _27099_ (.CLK(clknet_leaf_20_clk_sys),
    .D(_00716_),
    .RESET_B(net610),
    .Q(\top0.matmul0.matmul_stage_inst.a[6] ));
 sky130_fd_sc_hd__dfrtp_1 _27100_ (.CLK(clknet_leaf_16_clk_sys),
    .D(_00717_),
    .RESET_B(net611),
    .Q(\top0.matmul0.matmul_stage_inst.a[7] ));
 sky130_fd_sc_hd__dfrtp_1 _27101_ (.CLK(clknet_leaf_20_clk_sys),
    .D(_00718_),
    .RESET_B(net609),
    .Q(\top0.matmul0.matmul_stage_inst.a[8] ));
 sky130_fd_sc_hd__dfrtp_1 _27102_ (.CLK(clknet_leaf_20_clk_sys),
    .D(_00719_),
    .RESET_B(net610),
    .Q(\top0.matmul0.matmul_stage_inst.a[9] ));
 sky130_fd_sc_hd__dfrtp_1 _27103_ (.CLK(clknet_leaf_20_clk_sys),
    .D(_00720_),
    .RESET_B(net609),
    .Q(\top0.matmul0.matmul_stage_inst.a[10] ));
 sky130_fd_sc_hd__dfrtp_1 _27104_ (.CLK(clknet_leaf_21_clk_sys),
    .D(_00721_),
    .RESET_B(net610),
    .Q(\top0.matmul0.matmul_stage_inst.a[11] ));
 sky130_fd_sc_hd__dfrtp_1 _27105_ (.CLK(clknet_leaf_22_clk_sys),
    .D(_00722_),
    .RESET_B(net608),
    .Q(\top0.matmul0.matmul_stage_inst.a[12] ));
 sky130_fd_sc_hd__dfrtp_1 _27106_ (.CLK(clknet_leaf_21_clk_sys),
    .D(_00723_),
    .RESET_B(net610),
    .Q(\top0.matmul0.matmul_stage_inst.a[13] ));
 sky130_fd_sc_hd__dfrtp_1 _27107_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00724_),
    .RESET_B(net601),
    .Q(\top0.matmul0.op[0] ));
 sky130_fd_sc_hd__dfrtp_1 _27108_ (.CLK(clknet_leaf_8_clk_sys),
    .D(_00725_),
    .RESET_B(net592),
    .Q(\top0.matmul0.op[1] ));
 sky130_fd_sc_hd__dfstp_1 _27109_ (.CLK(clknet_leaf_89_clk_sys),
    .D(_00015_),
    .SET_B(net603),
    .Q(\top0.matmul0.state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _27110_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00016_),
    .RESET_B(net601),
    .Q(\top0.matmul0.state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27111_ (.CLK(clknet_leaf_9_clk_sys),
    .D(_00001_),
    .RESET_B(net595),
    .Q(\top0.matmul0.matmul_stage_inst.start ));
 sky130_fd_sc_hd__dfrtp_1 _27112_ (.CLK(clknet_leaf_87_clk_sys),
    .D(_00726_),
    .RESET_B(net644),
    .Q(\top0.pid_d.iterate_enable ));
 sky130_fd_sc_hd__dfrtp_2 _27113_ (.CLK(clknet_leaf_89_clk_sys),
    .D(_00727_),
    .RESET_B(net603),
    .Q(\top0.matmul0.start ));
 sky130_fd_sc_hd__dfrtp_4 _27114_ (.CLK(clknet_leaf_86_clk_sys),
    .D(_00728_),
    .RESET_B(net600),
    .Q(\top0.cordic0.in_valid ));
 sky130_fd_sc_hd__dfrtp_1 _27115_ (.CLK(clknet_leaf_89_clk_sys),
    .D(_00729_),
    .RESET_B(net603),
    .Q(\top0.clarke_done ));
 sky130_fd_sc_hd__dfrtp_1 _27116_ (.CLK(clknet_leaf_90_clk_sys),
    .D(_00730_),
    .RESET_B(net600),
    .Q(\top0.cordic_done ));
 sky130_fd_sc_hd__dfrtp_1 _27117_ (.CLK(clknet_leaf_33_clk_sys),
    .D(_00731_),
    .RESET_B(net665),
    .Q(\top0.c_out_calc[0] ));
 sky130_fd_sc_hd__dfrtp_1 _27118_ (.CLK(clknet_leaf_33_clk_sys),
    .D(_00732_),
    .RESET_B(net665),
    .Q(\top0.c_out_calc[1] ));
 sky130_fd_sc_hd__dfrtp_1 _27119_ (.CLK(clknet_leaf_33_clk_sys),
    .D(_00733_),
    .RESET_B(net665),
    .Q(\top0.c_out_calc[2] ));
 sky130_fd_sc_hd__dfrtp_1 _27120_ (.CLK(clknet_leaf_33_clk_sys),
    .D(_00734_),
    .RESET_B(net665),
    .Q(\top0.c_out_calc[3] ));
 sky130_fd_sc_hd__dfrtp_1 _27121_ (.CLK(clknet_3_6__leaf_clk_sys),
    .D(_00735_),
    .RESET_B(net665),
    .Q(\top0.c_out_calc[4] ));
 sky130_fd_sc_hd__dfrtp_1 _27122_ (.CLK(clknet_leaf_33_clk_sys),
    .D(_00736_),
    .RESET_B(net665),
    .Q(\top0.c_out_calc[5] ));
 sky130_fd_sc_hd__dfrtp_1 _27123_ (.CLK(clknet_leaf_30_clk_sys),
    .D(_00737_),
    .RESET_B(net623),
    .Q(\top0.c_out_calc[6] ));
 sky130_fd_sc_hd__dfrtp_1 _27124_ (.CLK(clknet_leaf_33_clk_sys),
    .D(_00738_),
    .RESET_B(net665),
    .Q(\top0.c_out_calc[7] ));
 sky130_fd_sc_hd__dfrtp_1 _27125_ (.CLK(clknet_leaf_33_clk_sys),
    .D(_00739_),
    .RESET_B(net665),
    .Q(\top0.c_out_calc[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27126_ (.CLK(clknet_3_6__leaf_clk_sys),
    .D(_00740_),
    .RESET_B(net665),
    .Q(\top0.c_out_calc[9] ));
 sky130_fd_sc_hd__dfrtp_1 _27127_ (.CLK(clknet_leaf_33_clk_sys),
    .D(_00741_),
    .RESET_B(net666),
    .Q(\top0.c_out_calc[10] ));
 sky130_fd_sc_hd__dfrtp_1 _27128_ (.CLK(clknet_leaf_33_clk_sys),
    .D(_00742_),
    .RESET_B(net666),
    .Q(\top0.c_out_calc[11] ));
 sky130_fd_sc_hd__dfrtp_1 _27129_ (.CLK(clknet_leaf_33_clk_sys),
    .D(_00743_),
    .RESET_B(net664),
    .Q(\top0.c_out_calc[12] ));
 sky130_fd_sc_hd__dfrtp_1 _27130_ (.CLK(clknet_leaf_33_clk_sys),
    .D(_00744_),
    .RESET_B(net665),
    .Q(\top0.c_out_calc[13] ));
 sky130_fd_sc_hd__dfrtp_1 _27131_ (.CLK(clknet_leaf_33_clk_sys),
    .D(_00745_),
    .RESET_B(net664),
    .Q(\top0.c_out_calc[14] ));
 sky130_fd_sc_hd__dfrtp_1 _27132_ (.CLK(clknet_leaf_32_clk_sys),
    .D(_00746_),
    .RESET_B(net664),
    .Q(\top0.c_out_calc[15] ));
 sky130_fd_sc_hd__dfrtp_1 _27133_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00747_),
    .RESET_B(net601),
    .Q(\top0.matmul0.op_in[0] ));
 sky130_fd_sc_hd__dfrtp_1 _27134_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00748_),
    .RESET_B(net601),
    .Q(\top0.matmul0.op_in[1] ));
 sky130_fd_sc_hd__dfrtp_1 _27135_ (.CLK(clknet_leaf_12_clk_sys),
    .D(_00749_),
    .RESET_B(net616),
    .Q(\top0.b_in_matmul[0] ));
 sky130_fd_sc_hd__dfrtp_1 _27136_ (.CLK(clknet_leaf_13_clk_sys),
    .D(_00750_),
    .RESET_B(net616),
    .Q(\top0.b_in_matmul[1] ));
 sky130_fd_sc_hd__dfrtp_1 _27137_ (.CLK(clknet_leaf_12_clk_sys),
    .D(_00751_),
    .RESET_B(net616),
    .Q(\top0.b_in_matmul[2] ));
 sky130_fd_sc_hd__dfrtp_1 _27138_ (.CLK(clknet_leaf_12_clk_sys),
    .D(_00752_),
    .RESET_B(net616),
    .Q(\top0.b_in_matmul[3] ));
 sky130_fd_sc_hd__dfrtp_1 _27139_ (.CLK(clknet_leaf_13_clk_sys),
    .D(_00753_),
    .RESET_B(net616),
    .Q(\top0.b_in_matmul[4] ));
 sky130_fd_sc_hd__dfrtp_1 _27140_ (.CLK(clknet_leaf_14_clk_sys),
    .D(_00754_),
    .RESET_B(net618),
    .Q(\top0.b_in_matmul[5] ));
 sky130_fd_sc_hd__dfrtp_1 _27141_ (.CLK(clknet_leaf_13_clk_sys),
    .D(_00755_),
    .RESET_B(net616),
    .Q(\top0.b_in_matmul[6] ));
 sky130_fd_sc_hd__dfrtp_1 _27142_ (.CLK(clknet_leaf_14_clk_sys),
    .D(_00756_),
    .RESET_B(net620),
    .Q(\top0.b_in_matmul[7] ));
 sky130_fd_sc_hd__dfrtp_1 _27143_ (.CLK(clknet_leaf_31_clk_sys),
    .D(_00757_),
    .RESET_B(net619),
    .Q(\top0.b_in_matmul[8] ));
 sky130_fd_sc_hd__dfrtp_1 _27144_ (.CLK(clknet_leaf_31_clk_sys),
    .D(_00758_),
    .RESET_B(net617),
    .Q(\top0.b_in_matmul[9] ));
 sky130_fd_sc_hd__dfrtp_1 _27145_ (.CLK(clknet_leaf_31_clk_sys),
    .D(_00759_),
    .RESET_B(net619),
    .Q(\top0.b_in_matmul[10] ));
 sky130_fd_sc_hd__dfrtp_1 _27146_ (.CLK(clknet_leaf_14_clk_sys),
    .D(_00760_),
    .RESET_B(net617),
    .Q(\top0.b_in_matmul[11] ));
 sky130_fd_sc_hd__dfrtp_1 _27147_ (.CLK(clknet_leaf_31_clk_sys),
    .D(_00761_),
    .RESET_B(net619),
    .Q(\top0.b_in_matmul[12] ));
 sky130_fd_sc_hd__dfrtp_1 _27148_ (.CLK(clknet_leaf_30_clk_sys),
    .D(_00762_),
    .RESET_B(net619),
    .Q(\top0.b_in_matmul[13] ));
 sky130_fd_sc_hd__dfrtp_1 _27149_ (.CLK(clknet_leaf_31_clk_sys),
    .D(_00763_),
    .RESET_B(net620),
    .Q(\top0.b_in_matmul[14] ));
 sky130_fd_sc_hd__dfrtp_1 _27150_ (.CLK(clknet_leaf_12_clk_sys),
    .D(_00764_),
    .RESET_B(net618),
    .Q(\top0.b_in_matmul[15] ));
 sky130_fd_sc_hd__dfrtp_1 _27151_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00765_),
    .RESET_B(net601),
    .Q(\top0.a_in_matmul[0] ));
 sky130_fd_sc_hd__dfrtp_1 _27152_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00766_),
    .RESET_B(net601),
    .Q(\top0.a_in_matmul[1] ));
 sky130_fd_sc_hd__dfrtp_1 _27153_ (.CLK(clknet_leaf_9_clk_sys),
    .D(_00767_),
    .RESET_B(net594),
    .Q(\top0.a_in_matmul[2] ));
 sky130_fd_sc_hd__dfrtp_1 _27154_ (.CLK(clknet_leaf_10_clk_sys),
    .D(_00768_),
    .RESET_B(net602),
    .Q(\top0.a_in_matmul[3] ));
 sky130_fd_sc_hd__dfrtp_1 _27155_ (.CLK(clknet_leaf_6_clk_sys),
    .D(_00769_),
    .RESET_B(net594),
    .Q(\top0.a_in_matmul[4] ));
 sky130_fd_sc_hd__dfrtp_1 _27156_ (.CLK(clknet_leaf_10_clk_sys),
    .D(_00770_),
    .RESET_B(net594),
    .Q(\top0.a_in_matmul[5] ));
 sky130_fd_sc_hd__dfrtp_1 _27157_ (.CLK(clknet_leaf_6_clk_sys),
    .D(_00771_),
    .RESET_B(net596),
    .Q(\top0.a_in_matmul[6] ));
 sky130_fd_sc_hd__dfrtp_1 _27158_ (.CLK(clknet_leaf_9_clk_sys),
    .D(_00772_),
    .RESET_B(net596),
    .Q(\top0.a_in_matmul[7] ));
 sky130_fd_sc_hd__dfrtp_1 _27159_ (.CLK(clknet_leaf_6_clk_sys),
    .D(_00773_),
    .RESET_B(net594),
    .Q(\top0.a_in_matmul[8] ));
 sky130_fd_sc_hd__dfrtp_1 _27160_ (.CLK(clknet_leaf_90_clk_sys),
    .D(_00774_),
    .RESET_B(net602),
    .Q(\top0.a_in_matmul[9] ));
 sky130_fd_sc_hd__dfrtp_1 _27161_ (.CLK(clknet_leaf_9_clk_sys),
    .D(_00775_),
    .RESET_B(net596),
    .Q(\top0.a_in_matmul[10] ));
 sky130_fd_sc_hd__dfrtp_1 _27162_ (.CLK(clknet_leaf_10_clk_sys),
    .D(_00776_),
    .RESET_B(net602),
    .Q(\top0.a_in_matmul[11] ));
 sky130_fd_sc_hd__dfrtp_1 _27163_ (.CLK(clknet_leaf_10_clk_sys),
    .D(_00777_),
    .RESET_B(net602),
    .Q(\top0.a_in_matmul[12] ));
 sky130_fd_sc_hd__dfrtp_1 _27164_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00778_),
    .RESET_B(net602),
    .Q(\top0.a_in_matmul[13] ));
 sky130_fd_sc_hd__dfrtp_1 _27165_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00779_),
    .RESET_B(net601),
    .Q(\top0.a_in_matmul[14] ));
 sky130_fd_sc_hd__dfrtp_1 _27166_ (.CLK(clknet_leaf_11_clk_sys),
    .D(_00780_),
    .RESET_B(net601),
    .Q(\top0.a_in_matmul[15] ));
 sky130_fd_sc_hd__dfrtp_4 _27167_ (.CLK(clknet_leaf_32_clk_sys),
    .D(_00781_),
    .RESET_B(net618),
    .Q(\top0.periodTop_r[0] ));
 sky130_fd_sc_hd__dfrtp_4 _27168_ (.CLK(clknet_leaf_32_clk_sys),
    .D(_00782_),
    .RESET_B(net664),
    .Q(\top0.periodTop_r[1] ));
 sky130_fd_sc_hd__dfrtp_4 _27169_ (.CLK(clknet_leaf_32_clk_sys),
    .D(_00783_),
    .RESET_B(net664),
    .Q(\top0.periodTop_r[2] ));
 sky130_fd_sc_hd__dfrtp_1 _27170_ (.CLK(clknet_leaf_12_clk_sys),
    .D(_00784_),
    .RESET_B(net618),
    .Q(\top0.periodTop_r[3] ));
 sky130_fd_sc_hd__dfrtp_4 _27171_ (.CLK(clknet_leaf_12_clk_sys),
    .D(_00785_),
    .RESET_B(net618),
    .Q(\top0.periodTop_r[4] ));
 sky130_fd_sc_hd__dfrtp_1 _27172_ (.CLK(clknet_leaf_12_clk_sys),
    .D(_00786_),
    .RESET_B(net618),
    .Q(\top0.periodTop_r[5] ));
 sky130_fd_sc_hd__dfrtp_1 _27173_ (.CLK(clknet_leaf_32_clk_sys),
    .D(_00787_),
    .RESET_B(net618),
    .Q(\top0.periodTop_r[6] ));
 sky130_fd_sc_hd__dfrtp_2 _27174_ (.CLK(clknet_leaf_32_clk_sys),
    .D(_00788_),
    .RESET_B(net618),
    .Q(\top0.periodTop_r[7] ));
 sky130_fd_sc_hd__dfrtp_2 _27175_ (.CLK(clknet_leaf_32_clk_sys),
    .D(_00789_),
    .RESET_B(net618),
    .Q(\top0.periodTop_r[8] ));
 sky130_fd_sc_hd__dfrtp_4 _27176_ (.CLK(clknet_leaf_32_clk_sys),
    .D(_00790_),
    .RESET_B(net619),
    .Q(\top0.periodTop_r[9] ));
 sky130_fd_sc_hd__dfrtp_1 _27177_ (.CLK(clknet_leaf_88_clk_sys),
    .D(_00791_),
    .RESET_B(net643),
    .Q(\top0.periodTop_r[10] ));
 sky130_fd_sc_hd__dfrtp_1 _27178_ (.CLK(clknet_leaf_88_clk_sys),
    .D(_00792_),
    .RESET_B(net642),
    .Q(\top0.periodTop_r[11] ));
 sky130_fd_sc_hd__dfrtp_1 _27179_ (.CLK(clknet_leaf_57_clk_sys),
    .D(_00793_),
    .RESET_B(net643),
    .Q(\top0.periodTop_r[12] ));
 sky130_fd_sc_hd__dfrtp_1 _27180_ (.CLK(clknet_leaf_88_clk_sys),
    .D(_00794_),
    .RESET_B(net643),
    .Q(\top0.periodTop_r[13] ));
 sky130_fd_sc_hd__dfrtp_1 _27181_ (.CLK(clknet_leaf_88_clk_sys),
    .D(_00795_),
    .RESET_B(net643),
    .Q(\top0.periodTop_r[14] ));
 sky130_fd_sc_hd__dfrtp_1 _27182_ (.CLK(clknet_leaf_88_clk_sys),
    .D(_00796_),
    .RESET_B(net642),
    .Q(\top0.periodTop_r[15] ));
 sky130_fd_sc_hd__dfrtp_1 _27183_ (.CLK(clknet_leaf_58_clk_sys),
    .D(_00797_),
    .RESET_B(net643),
    .Q(\top0.currT_r[0] ));
 sky130_fd_sc_hd__dfrtp_2 _27184_ (.CLK(clknet_leaf_59_clk_sys),
    .D(_00798_),
    .RESET_B(net644),
    .Q(\top0.currT_r[1] ));
 sky130_fd_sc_hd__dfrtp_2 _27185_ (.CLK(clknet_leaf_58_clk_sys),
    .D(_00799_),
    .RESET_B(net644),
    .Q(\top0.currT_r[2] ));
 sky130_fd_sc_hd__dfrtp_2 _27186_ (.CLK(clknet_leaf_57_clk_sys),
    .D(_00800_),
    .RESET_B(net645),
    .Q(\top0.currT_r[3] ));
 sky130_fd_sc_hd__dfrtp_2 _27187_ (.CLK(clknet_leaf_56_clk_sys),
    .D(_00801_),
    .RESET_B(net666),
    .Q(\top0.currT_r[4] ));
 sky130_fd_sc_hd__dfrtp_2 _27188_ (.CLK(clknet_leaf_56_clk_sys),
    .D(_00802_),
    .RESET_B(net666),
    .Q(\top0.currT_r[5] ));
 sky130_fd_sc_hd__dfrtp_1 _27189_ (.CLK(clknet_leaf_54_clk_sys),
    .D(_00803_),
    .RESET_B(net668),
    .Q(\top0.currT_r[6] ));
 sky130_fd_sc_hd__dfrtp_1 _27190_ (.CLK(clknet_leaf_55_clk_sys),
    .D(_00804_),
    .RESET_B(net668),
    .Q(\top0.currT_r[7] ));
 sky130_fd_sc_hd__dfrtp_1 _27191_ (.CLK(clknet_leaf_56_clk_sys),
    .D(_00805_),
    .RESET_B(net668),
    .Q(\top0.currT_r[8] ));
 sky130_fd_sc_hd__dfrtp_2 _27192_ (.CLK(clknet_leaf_56_clk_sys),
    .D(_00806_),
    .RESET_B(net668),
    .Q(\top0.currT_r[9] ));
 sky130_fd_sc_hd__dfrtp_2 _27193_ (.CLK(clknet_leaf_56_clk_sys),
    .D(_00807_),
    .RESET_B(net668),
    .Q(\top0.currT_r[10] ));
 sky130_fd_sc_hd__dfrtp_1 _27194_ (.CLK(clknet_leaf_56_clk_sys),
    .D(_00808_),
    .RESET_B(net666),
    .Q(\top0.currT_r[11] ));
 sky130_fd_sc_hd__dfrtp_1 _27195_ (.CLK(clknet_leaf_56_clk_sys),
    .D(_00809_),
    .RESET_B(net666),
    .Q(\top0.currT_r[12] ));
 sky130_fd_sc_hd__dfrtp_4 _27196_ (.CLK(clknet_leaf_57_clk_sys),
    .D(_00810_),
    .RESET_B(net664),
    .Q(\top0.currT_r[13] ));
 sky130_fd_sc_hd__dfrtp_4 _27197_ (.CLK(clknet_leaf_57_clk_sys),
    .D(_00811_),
    .RESET_B(net664),
    .Q(\top0.currT_r[14] ));
 sky130_fd_sc_hd__dfrtp_1 _27198_ (.CLK(clknet_leaf_32_clk_sys),
    .D(_00812_),
    .RESET_B(net664),
    .Q(\top0.currT_r[15] ));
 sky130_fd_sc_hd__dfrtp_1 _27199_ (.CLK(clknet_leaf_91_clk_sys),
    .D(_00813_),
    .RESET_B(net599),
    .Q(\top0.cordic0.slte0.opB[2] ));
 sky130_fd_sc_hd__dfrtp_1 _27200_ (.CLK(clknet_leaf_91_clk_sys),
    .D(_00814_),
    .RESET_B(net600),
    .Q(\top0.cordic0.slte0.opB[3] ));
 sky130_fd_sc_hd__dfrtp_1 _27201_ (.CLK(clknet_leaf_91_clk_sys),
    .D(_00815_),
    .RESET_B(net600),
    .Q(\top0.cordic0.slte0.opB[4] ));
 sky130_fd_sc_hd__dfrtp_1 _27202_ (.CLK(clknet_leaf_92_clk_sys),
    .D(_00816_),
    .RESET_B(net599),
    .Q(\top0.cordic0.slte0.opB[5] ));
 sky130_fd_sc_hd__dfrtp_1 _27203_ (.CLK(clknet_leaf_91_clk_sys),
    .D(_00817_),
    .RESET_B(net599),
    .Q(\top0.cordic0.slte0.opB[6] ));
 sky130_fd_sc_hd__dfrtp_1 _27204_ (.CLK(clknet_leaf_92_clk_sys),
    .D(_00818_),
    .RESET_B(net599),
    .Q(\top0.cordic0.slte0.opB[7] ));
 sky130_fd_sc_hd__dfrtp_1 _27205_ (.CLK(clknet_leaf_92_clk_sys),
    .D(_00819_),
    .RESET_B(net599),
    .Q(\top0.cordic0.slte0.opB[8] ));
 sky130_fd_sc_hd__dfrtp_1 _27206_ (.CLK(clknet_leaf_92_clk_sys),
    .D(_00820_),
    .RESET_B(net600),
    .Q(\top0.cordic0.slte0.opB[9] ));
 sky130_fd_sc_hd__dfrtp_1 _27207_ (.CLK(clknet_leaf_93_clk_sys),
    .D(_00821_),
    .RESET_B(net600),
    .Q(\top0.cordic0.slte0.opB[10] ));
 sky130_fd_sc_hd__dfrtp_1 _27208_ (.CLK(clknet_leaf_93_clk_sys),
    .D(_00822_),
    .RESET_B(net600),
    .Q(\top0.cordic0.slte0.opB[11] ));
 sky130_fd_sc_hd__dfrtp_1 _27209_ (.CLK(clknet_leaf_6_clk_sys),
    .D(_00823_),
    .RESET_B(net591),
    .Q(\top0.cordic0.slte0.opB[12] ));
 sky130_fd_sc_hd__dfrtp_1 _27210_ (.CLK(clknet_leaf_93_clk_sys),
    .D(_00824_),
    .RESET_B(net591),
    .Q(\top0.cordic0.slte0.opB[13] ));
 sky130_fd_sc_hd__dfrtp_1 _27211_ (.CLK(clknet_leaf_6_clk_sys),
    .D(_00825_),
    .RESET_B(net591),
    .Q(\top0.cordic0.slte0.opB[14] ));
 sky130_fd_sc_hd__dfrtp_1 _27212_ (.CLK(clknet_leaf_6_clk_sys),
    .D(_00826_),
    .RESET_B(net598),
    .Q(\top0.cordic0.slte0.opB[15] ));
 sky130_fd_sc_hd__dfstp_1 _27213_ (.CLK(clknet_leaf_87_clk_sys),
    .D(_00827_),
    .SET_B(net642),
    .Q(\top0.ready ));
 sky130_fd_sc_hd__dfxtp_2 _27214_ (.CLK(clknet_3_4__leaf_clk_mosi),
    .D(_00828_),
    .Q(\spi0.data_packed[0] ));
 sky130_fd_sc_hd__dfxtp_2 _27215_ (.CLK(clknet_3_1__leaf_clk_mosi),
    .D(_00829_),
    .Q(\spi0.data_packed[1] ));
 sky130_fd_sc_hd__dfxtp_1 _27216_ (.CLK(clknet_3_1__leaf_clk_mosi),
    .D(_00830_),
    .Q(\spi0.data_packed[2] ));
 sky130_fd_sc_hd__dfxtp_2 _27217_ (.CLK(clknet_3_1__leaf_clk_mosi),
    .D(_00831_),
    .Q(\spi0.data_packed[3] ));
 sky130_fd_sc_hd__dfxtp_1 _27218_ (.CLK(clknet_3_1__leaf_clk_mosi),
    .D(_00832_),
    .Q(\spi0.data_packed[4] ));
 sky130_fd_sc_hd__dfxtp_2 _27219_ (.CLK(clknet_3_1__leaf_clk_mosi),
    .D(_00833_),
    .Q(\spi0.data_packed[5] ));
 sky130_fd_sc_hd__dfxtp_2 _27220_ (.CLK(clknet_3_5__leaf_clk_mosi),
    .D(_00834_),
    .Q(\spi0.data_packed[6] ));
 sky130_fd_sc_hd__dfxtp_1 _27221_ (.CLK(clknet_3_5__leaf_clk_mosi),
    .D(_00835_),
    .Q(\spi0.data_packed[7] ));
 sky130_fd_sc_hd__dfxtp_2 _27222_ (.CLK(clknet_3_4__leaf_clk_mosi),
    .D(_00836_),
    .Q(\spi0.data_packed[8] ));
 sky130_fd_sc_hd__dfxtp_1 _27223_ (.CLK(clknet_3_5__leaf_clk_mosi),
    .D(_00837_),
    .Q(\spi0.data_packed[9] ));
 sky130_fd_sc_hd__dfxtp_1 _27224_ (.CLK(clknet_3_4__leaf_clk_mosi),
    .D(_00838_),
    .Q(\spi0.data_packed[10] ));
 sky130_fd_sc_hd__dfxtp_2 _27225_ (.CLK(clknet_3_5__leaf_clk_mosi),
    .D(_00839_),
    .Q(\spi0.data_packed[11] ));
 sky130_fd_sc_hd__dfxtp_1 _27226_ (.CLK(clknet_3_4__leaf_clk_mosi),
    .D(_00840_),
    .Q(\spi0.data_packed[12] ));
 sky130_fd_sc_hd__dfxtp_1 _27227_ (.CLK(clknet_3_4__leaf_clk_mosi),
    .D(_00841_),
    .Q(\spi0.data_packed[13] ));
 sky130_fd_sc_hd__dfxtp_1 _27228_ (.CLK(clknet_3_4__leaf_clk_mosi),
    .D(_00842_),
    .Q(\spi0.data_packed[14] ));
 sky130_fd_sc_hd__dfxtp_2 _27229_ (.CLK(clknet_3_1__leaf_clk_mosi),
    .D(_00843_),
    .Q(\spi0.data_packed[15] ));
 sky130_fd_sc_hd__dfxtp_1 _27230_ (.CLK(clknet_3_1__leaf_clk_mosi),
    .D(_00844_),
    .Q(\spi0.data_packed[16] ));
 sky130_fd_sc_hd__dfxtp_1 _27231_ (.CLK(clknet_3_5__leaf_clk_mosi),
    .D(_00845_),
    .Q(\spi0.data_packed[17] ));
 sky130_fd_sc_hd__dfxtp_1 _27232_ (.CLK(clknet_3_4__leaf_clk_mosi),
    .D(_00846_),
    .Q(\spi0.data_packed[18] ));
 sky130_fd_sc_hd__dfxtp_1 _27233_ (.CLK(clknet_3_6__leaf_clk_mosi),
    .D(_00847_),
    .Q(\spi0.data_packed[19] ));
 sky130_fd_sc_hd__dfxtp_1 _27234_ (.CLK(clknet_3_6__leaf_clk_mosi),
    .D(_00848_),
    .Q(\spi0.data_packed[20] ));
 sky130_fd_sc_hd__dfxtp_1 _27235_ (.CLK(clknet_3_7__leaf_clk_mosi),
    .D(_00849_),
    .Q(\spi0.data_packed[21] ));
 sky130_fd_sc_hd__dfxtp_1 _27236_ (.CLK(clknet_3_7__leaf_clk_mosi),
    .D(_00850_),
    .Q(\spi0.data_packed[22] ));
 sky130_fd_sc_hd__dfxtp_1 _27237_ (.CLK(clknet_3_7__leaf_clk_mosi),
    .D(_00851_),
    .Q(\spi0.data_packed[23] ));
 sky130_fd_sc_hd__dfxtp_1 _27238_ (.CLK(clknet_3_7__leaf_clk_mosi),
    .D(_00852_),
    .Q(\spi0.data_packed[24] ));
 sky130_fd_sc_hd__dfxtp_1 _27239_ (.CLK(clknet_3_7__leaf_clk_mosi),
    .D(_00853_),
    .Q(\spi0.data_packed[25] ));
 sky130_fd_sc_hd__dfxtp_1 _27240_ (.CLK(clknet_3_7__leaf_clk_mosi),
    .D(_00854_),
    .Q(\spi0.data_packed[26] ));
 sky130_fd_sc_hd__dfxtp_1 _27241_ (.CLK(clknet_3_7__leaf_clk_mosi),
    .D(_00855_),
    .Q(\spi0.data_packed[27] ));
 sky130_fd_sc_hd__dfxtp_1 _27242_ (.CLK(clknet_3_7__leaf_clk_mosi),
    .D(_00856_),
    .Q(\spi0.data_packed[28] ));
 sky130_fd_sc_hd__dfxtp_1 _27243_ (.CLK(clknet_3_7__leaf_clk_mosi),
    .D(_00857_),
    .Q(\spi0.data_packed[29] ));
 sky130_fd_sc_hd__dfxtp_1 _27244_ (.CLK(clknet_3_5__leaf_clk_mosi),
    .D(_00858_),
    .Q(\spi0.data_packed[30] ));
 sky130_fd_sc_hd__dfxtp_1 _27245_ (.CLK(clknet_3_5__leaf_clk_mosi),
    .D(_00859_),
    .Q(\spi0.data_packed[31] ));
 sky130_fd_sc_hd__dfxtp_1 _27246_ (.CLK(clknet_3_0__leaf_clk_mosi),
    .D(_00860_),
    .Q(\spi0.data_packed[32] ));
 sky130_fd_sc_hd__dfxtp_1 _27247_ (.CLK(clknet_3_2__leaf_clk_mosi),
    .D(_00861_),
    .Q(\spi0.data_packed[33] ));
 sky130_fd_sc_hd__dfxtp_1 _27248_ (.CLK(clknet_3_2__leaf_clk_mosi),
    .D(_00862_),
    .Q(\spi0.data_packed[34] ));
 sky130_fd_sc_hd__dfxtp_1 _27249_ (.CLK(clknet_3_2__leaf_clk_mosi),
    .D(_00863_),
    .Q(\spi0.data_packed[35] ));
 sky130_fd_sc_hd__dfxtp_1 _27250_ (.CLK(clknet_3_2__leaf_clk_mosi),
    .D(_00864_),
    .Q(\spi0.data_packed[36] ));
 sky130_fd_sc_hd__dfxtp_1 _27251_ (.CLK(clknet_3_2__leaf_clk_mosi),
    .D(_00865_),
    .Q(\spi0.data_packed[37] ));
 sky130_fd_sc_hd__dfxtp_1 _27252_ (.CLK(clknet_3_2__leaf_clk_mosi),
    .D(_00866_),
    .Q(\spi0.data_packed[38] ));
 sky130_fd_sc_hd__dfxtp_1 _27253_ (.CLK(clknet_3_2__leaf_clk_mosi),
    .D(_00867_),
    .Q(\spi0.data_packed[39] ));
 sky130_fd_sc_hd__dfxtp_1 _27254_ (.CLK(clknet_3_2__leaf_clk_mosi),
    .D(_00868_),
    .Q(\spi0.data_packed[40] ));
 sky130_fd_sc_hd__dfxtp_1 _27255_ (.CLK(clknet_3_2__leaf_clk_mosi),
    .D(_00869_),
    .Q(\spi0.data_packed[41] ));
 sky130_fd_sc_hd__dfxtp_1 _27256_ (.CLK(clknet_3_2__leaf_clk_mosi),
    .D(_00870_),
    .Q(\spi0.data_packed[42] ));
 sky130_fd_sc_hd__dfxtp_1 _27257_ (.CLK(clknet_3_3__leaf_clk_mosi),
    .D(_00871_),
    .Q(\spi0.data_packed[43] ));
 sky130_fd_sc_hd__dfxtp_1 _27258_ (.CLK(clknet_3_3__leaf_clk_mosi),
    .D(_00872_),
    .Q(\spi0.data_packed[44] ));
 sky130_fd_sc_hd__dfxtp_1 _27259_ (.CLK(clknet_3_3__leaf_clk_mosi),
    .D(_00873_),
    .Q(\spi0.data_packed[45] ));
 sky130_fd_sc_hd__dfxtp_1 _27260_ (.CLK(clknet_3_3__leaf_clk_mosi),
    .D(_00874_),
    .Q(\spi0.data_packed[46] ));
 sky130_fd_sc_hd__dfxtp_1 _27261_ (.CLK(clknet_3_0__leaf_clk_mosi),
    .D(_00875_),
    .Q(\spi0.data_packed[47] ));
 sky130_fd_sc_hd__dfxtp_1 _27262_ (.CLK(clknet_3_4__leaf_clk_mosi),
    .D(_00876_),
    .Q(\spi0.data_packed[48] ));
 sky130_fd_sc_hd__dfxtp_1 _27263_ (.CLK(clknet_3_6__leaf_clk_mosi),
    .D(_00877_),
    .Q(\spi0.data_packed[49] ));
 sky130_fd_sc_hd__dfxtp_1 _27264_ (.CLK(clknet_3_6__leaf_clk_mosi),
    .D(_00878_),
    .Q(\spi0.data_packed[50] ));
 sky130_fd_sc_hd__dfxtp_1 _27265_ (.CLK(clknet_3_6__leaf_clk_mosi),
    .D(_00879_),
    .Q(\spi0.data_packed[51] ));
 sky130_fd_sc_hd__dfxtp_1 _27266_ (.CLK(clknet_3_6__leaf_clk_mosi),
    .D(_00880_),
    .Q(\spi0.data_packed[52] ));
 sky130_fd_sc_hd__dfxtp_1 _27267_ (.CLK(clknet_3_6__leaf_clk_mosi),
    .D(_00881_),
    .Q(\spi0.data_packed[53] ));
 sky130_fd_sc_hd__dfxtp_1 _27268_ (.CLK(clknet_3_6__leaf_clk_mosi),
    .D(_00882_),
    .Q(\spi0.data_packed[54] ));
 sky130_fd_sc_hd__dfxtp_1 _27269_ (.CLK(clknet_3_6__leaf_clk_mosi),
    .D(_00883_),
    .Q(\spi0.data_packed[55] ));
 sky130_fd_sc_hd__dfxtp_1 _27270_ (.CLK(clknet_3_6__leaf_clk_mosi),
    .D(_00884_),
    .Q(\spi0.data_packed[56] ));
 sky130_fd_sc_hd__dfxtp_1 _27271_ (.CLK(clknet_3_7__leaf_clk_mosi),
    .D(_00885_),
    .Q(\spi0.data_packed[57] ));
 sky130_fd_sc_hd__dfxtp_1 _27272_ (.CLK(clknet_3_7__leaf_clk_mosi),
    .D(_00886_),
    .Q(\spi0.data_packed[58] ));
 sky130_fd_sc_hd__dfxtp_1 _27273_ (.CLK(clknet_3_7__leaf_clk_mosi),
    .D(_00887_),
    .Q(\spi0.data_packed[59] ));
 sky130_fd_sc_hd__dfxtp_1 _27274_ (.CLK(clknet_3_7__leaf_clk_mosi),
    .D(_00888_),
    .Q(\spi0.data_packed[60] ));
 sky130_fd_sc_hd__dfxtp_1 _27275_ (.CLK(clknet_3_7__leaf_clk_mosi),
    .D(_00889_),
    .Q(\spi0.data_packed[61] ));
 sky130_fd_sc_hd__dfxtp_1 _27276_ (.CLK(clknet_3_7__leaf_clk_mosi),
    .D(_00890_),
    .Q(\spi0.data_packed[62] ));
 sky130_fd_sc_hd__dfxtp_1 _27277_ (.CLK(clknet_3_5__leaf_clk_mosi),
    .D(_00891_),
    .Q(\spi0.data_packed[63] ));
 sky130_fd_sc_hd__dfxtp_1 _27278_ (.CLK(clknet_3_4__leaf_clk_mosi),
    .D(_00892_),
    .Q(\spi0.data_packed[64] ));
 sky130_fd_sc_hd__dfxtp_1 _27279_ (.CLK(clknet_3_4__leaf_clk_mosi),
    .D(_00893_),
    .Q(\spi0.data_packed[65] ));
 sky130_fd_sc_hd__dfxtp_1 _27280_ (.CLK(clknet_3_1__leaf_clk_mosi),
    .D(_00894_),
    .Q(\spi0.data_packed[66] ));
 sky130_fd_sc_hd__dfxtp_1 _27281_ (.CLK(clknet_3_0__leaf_clk_mosi),
    .D(_00895_),
    .Q(\spi0.data_packed[67] ));
 sky130_fd_sc_hd__dfxtp_1 _27282_ (.CLK(clknet_3_3__leaf_clk_mosi),
    .D(_00896_),
    .Q(\spi0.data_packed[68] ));
 sky130_fd_sc_hd__dfxtp_1 _27283_ (.CLK(clknet_3_0__leaf_clk_mosi),
    .D(_00897_),
    .Q(\spi0.data_packed[69] ));
 sky130_fd_sc_hd__dfxtp_1 _27284_ (.CLK(clknet_3_2__leaf_clk_mosi),
    .D(_00898_),
    .Q(\spi0.data_packed[70] ));
 sky130_fd_sc_hd__dfxtp_1 _27285_ (.CLK(clknet_3_2__leaf_clk_mosi),
    .D(_00899_),
    .Q(\spi0.data_packed[71] ));
 sky130_fd_sc_hd__dfxtp_1 _27286_ (.CLK(clknet_3_2__leaf_clk_mosi),
    .D(_00900_),
    .Q(\spi0.data_packed[72] ));
 sky130_fd_sc_hd__dfxtp_1 _27287_ (.CLK(clknet_3_3__leaf_clk_mosi),
    .D(_00901_),
    .Q(\spi0.data_packed[73] ));
 sky130_fd_sc_hd__dfxtp_1 _27288_ (.CLK(clknet_3_0__leaf_clk_mosi),
    .D(_00902_),
    .Q(\spi0.data_packed[74] ));
 sky130_fd_sc_hd__dfxtp_1 _27289_ (.CLK(clknet_3_3__leaf_clk_mosi),
    .D(_00903_),
    .Q(\spi0.data_packed[75] ));
 sky130_fd_sc_hd__dfxtp_1 _27290_ (.CLK(clknet_3_3__leaf_clk_mosi),
    .D(_00904_),
    .Q(\spi0.data_packed[76] ));
 sky130_fd_sc_hd__dfxtp_1 _27291_ (.CLK(clknet_3_3__leaf_clk_mosi),
    .D(_00905_),
    .Q(\spi0.data_packed[77] ));
 sky130_fd_sc_hd__dfxtp_1 _27292_ (.CLK(clknet_3_0__leaf_clk_mosi),
    .D(_00906_),
    .Q(\spi0.data_packed[78] ));
 sky130_fd_sc_hd__dfxtp_1 _27293_ (.CLK(clknet_3_0__leaf_clk_mosi),
    .D(_00907_),
    .Q(\spi0.data_packed[79] ));
 sky130_fd_sc_hd__dfxtp_1 _27294_ (.CLK(clknet_3_0__leaf_clk_mosi),
    .D(_00908_),
    .Q(\spi0.opcode[0] ));
 sky130_fd_sc_hd__dfxtp_1 _27295_ (.CLK(clknet_3_0__leaf_clk_mosi),
    .D(_00909_),
    .Q(\spi0.opcode[1] ));
 sky130_fd_sc_hd__dfxtp_1 _27296_ (.CLK(clknet_3_0__leaf_clk_mosi),
    .D(_00910_),
    .Q(\spi0.opcode[2] ));
 sky130_fd_sc_hd__dfxtp_1 _27297_ (.CLK(clknet_3_1__leaf_clk_mosi),
    .D(_00911_),
    .Q(\spi0.opcode[3] ));
 sky130_fd_sc_hd__dfxtp_1 _27298_ (.CLK(clknet_3_1__leaf_clk_mosi),
    .D(_00912_),
    .Q(\spi0.opcode[4] ));
 sky130_fd_sc_hd__dfxtp_1 _27299_ (.CLK(clknet_3_1__leaf_clk_mosi),
    .D(_00913_),
    .Q(\spi0.opcode[5] ));
 sky130_fd_sc_hd__dfxtp_1 _27300_ (.CLK(clknet_3_1__leaf_clk_mosi),
    .D(_00914_),
    .Q(\spi0.opcode[6] ));
 sky130_fd_sc_hd__dfxtp_1 _27301_ (.CLK(clknet_3_1__leaf_clk_mosi),
    .D(_00915_),
    .Q(\spi0.opcode[7] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Right_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Right_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Right_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Right_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Right_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Right_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Right_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Right_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Right_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Right_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Right_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Right_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Right_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Right_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Right_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Right_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Right_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Right_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Right_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Right_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Right_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Right_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Right_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Right_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Right_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Right_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Right_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Right_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Right_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Left_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Left_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Left_365 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Left_366 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Left_367 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Left_368 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Left_369 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Left_370 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Left_371 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Left_372 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Left_373 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Left_374 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Left_375 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Left_376 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Left_377 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Left_378 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Left_379 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Left_380 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Left_381 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Left_382 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Left_383 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Left_384 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Left_385 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Left_386 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Left_387 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Left_388 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Left_389 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Left_390 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Left_391 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Left_392 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Left_393 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Left_394 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Left_395 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Left_396 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Left_397 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Left_398 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Left_399 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Left_400 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Left_401 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Left_402 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Left_403 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Left_404 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Left_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4710 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(cs),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(rstb),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(spi_mosi),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 output4 (.A(net4),
    .X(pwmA));
 sky130_fd_sc_hd__clkbuf_4 output5 (.A(net5),
    .X(pwmB));
 sky130_fd_sc_hd__clkbuf_4 output6 (.A(net6),
    .X(pwmC));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(ready));
 sky130_fd_sc_hd__clkbuf_2 max_cap8 (.A(_03432_),
    .X(net8));
 sky130_fd_sc_hd__buf_1 wire9 (.A(_02593_),
    .X(net9));
 sky130_fd_sc_hd__buf_1 max_cap10 (.A(net1012),
    .X(net10));
 sky130_fd_sc_hd__buf_1 max_cap11 (.A(net12),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 max_cap12 (.A(_05066_),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 max_cap13 (.A(_07699_),
    .X(net13));
 sky130_fd_sc_hd__buf_2 max_cap14 (.A(_07141_),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 max_cap15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 wire16 (.A(net17),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 max_cap17 (.A(_05430_),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(net19),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 fanout19 (.A(\spi0.data_packed[14] ),
    .X(net19));
 sky130_fd_sc_hd__buf_2 fanout20 (.A(net22),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout21 (.A(net22),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 fanout22 (.A(net23),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 fanout23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__buf_2 fanout24 (.A(\top0.periodTop_r[15] ),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 fanout25 (.A(net27),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 fanout26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 fanout28 (.A(net1030),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 fanout29 (.A(\top0.periodTop_r[14] ),
    .X(net29));
 sky130_fd_sc_hd__buf_4 fanout30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__buf_4 fanout31 (.A(net32),
    .X(net31));
 sky130_fd_sc_hd__buf_4 fanout32 (.A(\top0.periodTop_r[13] ),
    .X(net32));
 sky130_fd_sc_hd__buf_4 fanout33 (.A(net35),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(\top0.periodTop_r[12] ),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(\top0.periodTop_r[11] ),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__buf_4 fanout40 (.A(\top0.periodTop_r[10] ),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 fanout41 (.A(\top0.periodTop_r[9] ),
    .X(net41));
 sky130_fd_sc_hd__buf_4 fanout42 (.A(\top0.periodTop_r[9] ),
    .X(net42));
 sky130_fd_sc_hd__buf_4 fanout43 (.A(\top0.periodTop_r[8] ),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 fanout44 (.A(\top0.periodTop_r[8] ),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(\top0.periodTop_r[7] ),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 fanout46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__buf_4 fanout47 (.A(\top0.periodTop_r[7] ),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__buf_4 fanout49 (.A(\top0.periodTop_r[6] ),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(\top0.periodTop_r[6] ),
    .X(net50));
 sky130_fd_sc_hd__buf_4 fanout51 (.A(net1027),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 fanout52 (.A(net1027),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 fanout53 (.A(\top0.periodTop_r[5] ),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(\top0.periodTop_r[4] ),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 fanout55 (.A(\top0.periodTop_r[4] ),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 fanout56 (.A(net58),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 fanout57 (.A(net58),
    .X(net57));
 sky130_fd_sc_hd__buf_4 fanout58 (.A(\top0.periodTop_r[3] ),
    .X(net58));
 sky130_fd_sc_hd__buf_4 fanout59 (.A(\top0.periodTop_r[2] ),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(\top0.periodTop_r[2] ),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 fanout61 (.A(\top0.periodTop_r[2] ),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(\top0.periodTop_r[1] ),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net64),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 fanout64 (.A(\top0.periodTop_r[1] ),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 fanout65 (.A(net67),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 fanout66 (.A(net67),
    .X(net66));
 sky130_fd_sc_hd__buf_2 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__buf_4 fanout68 (.A(\top0.periodTop_r[0] ),
    .X(net68));
 sky130_fd_sc_hd__buf_2 fanout69 (.A(\top0.matmul0.op[1] ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__buf_2 fanout71 (.A(\top0.matmul0.op[1] ),
    .X(net71));
 sky130_fd_sc_hd__buf_2 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__buf_2 fanout73 (.A(net74),
    .X(net73));
 sky130_fd_sc_hd__buf_2 fanout74 (.A(\top0.matmul0.op[0] ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 fanout75 (.A(\top0.matmul0.alpha_pass[8] ),
    .X(net75));
 sky130_fd_sc_hd__buf_4 fanout76 (.A(\top0.matmul0.alpha_pass[5] ),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_4 fanout77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_4 fanout78 (.A(net81),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_4 fanout79 (.A(net80),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 fanout80 (.A(net81),
    .X(net80));
 sky130_fd_sc_hd__buf_2 fanout81 (.A(\top0.cordic0.vec[1][17] ),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 fanout82 (.A(net84),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 fanout83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__buf_2 fanout84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 fanout85 (.A(\top0.cordic0.vec[1][17] ),
    .X(net85));
 sky130_fd_sc_hd__buf_4 fanout86 (.A(net89),
    .X(net86));
 sky130_fd_sc_hd__buf_2 fanout87 (.A(net89),
    .X(net87));
 sky130_fd_sc_hd__buf_4 fanout88 (.A(net89),
    .X(net88));
 sky130_fd_sc_hd__buf_4 fanout89 (.A(\top0.cordic0.vec[1][16] ),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 fanout90 (.A(net93),
    .X(net90));
 sky130_fd_sc_hd__buf_2 fanout91 (.A(net92),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 fanout92 (.A(net93),
    .X(net92));
 sky130_fd_sc_hd__buf_2 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__buf_4 fanout94 (.A(\top0.cordic0.vec[1][15] ),
    .X(net94));
 sky130_fd_sc_hd__buf_2 fanout95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__buf_2 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__buf_4 fanout97 (.A(\top0.cordic0.vec[1][14] ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 fanout98 (.A(\top0.cordic0.vec[1][14] ),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_4 fanout99 (.A(net101),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_4 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 fanout101 (.A(net102),
    .X(net101));
 sky130_fd_sc_hd__buf_4 fanout102 (.A(\top0.cordic0.vec[1][13] ),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 fanout103 (.A(\top0.cordic0.vec[1][13] ),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_8 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_4 fanout106 (.A(\top0.cordic0.vec[1][12] ),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 fanout107 (.A(net108),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 fanout108 (.A(\top0.cordic0.vec[1][12] ),
    .X(net108));
 sky130_fd_sc_hd__buf_4 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__buf_2 fanout110 (.A(net112),
    .X(net110));
 sky130_fd_sc_hd__buf_4 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(\top0.cordic0.vec[1][11] ),
    .X(net113));
 sky130_fd_sc_hd__buf_4 fanout114 (.A(net116),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 fanout115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 fanout116 (.A(net1031),
    .X(net116));
 sky130_fd_sc_hd__buf_1 fanout117 (.A(\top0.cordic0.vec[1][10] ),
    .X(net117));
 sky130_fd_sc_hd__buf_4 fanout118 (.A(net120),
    .X(net118));
 sky130_fd_sc_hd__buf_4 fanout119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_4 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__buf_4 fanout121 (.A(\top0.cordic0.vec[1][9] ),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_8 fanout122 (.A(net125),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_4 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_4 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__buf_2 fanout125 (.A(\top0.cordic0.vec[1][8] ),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_4 fanout126 (.A(net128),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 fanout127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__buf_4 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__buf_4 fanout129 (.A(\top0.cordic0.vec[1][7] ),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(\top0.cordic0.vec[1][6] ),
    .X(net130));
 sky130_fd_sc_hd__buf_4 fanout131 (.A(net134),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 fanout132 (.A(net134),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_8 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__buf_2 fanout134 (.A(\top0.cordic0.vec[1][6] ),
    .X(net134));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(net137),
    .X(net135));
 sky130_fd_sc_hd__buf_2 fanout136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__buf_2 fanout137 (.A(\top0.cordic0.vec[1][5] ),
    .X(net137));
 sky130_fd_sc_hd__buf_2 fanout138 (.A(net140),
    .X(net138));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(\top0.cordic0.vec[1][5] ),
    .X(net139));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout140 (.A(\top0.cordic0.vec[1][5] ),
    .X(net140));
 sky130_fd_sc_hd__buf_2 fanout141 (.A(net143),
    .X(net141));
 sky130_fd_sc_hd__buf_2 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_4 fanout143 (.A(\top0.cordic0.vec[1][4] ),
    .X(net143));
 sky130_fd_sc_hd__buf_2 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_4 fanout145 (.A(\top0.cordic0.vec[1][4] ),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_4 fanout146 (.A(net148),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_4 fanout147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_4 fanout149 (.A(\top0.cordic0.vec[1][3] ),
    .X(net149));
 sky130_fd_sc_hd__buf_4 fanout150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_4 fanout151 (.A(\top0.cordic0.vec[1][3] ),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 fanout152 (.A(net154),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 fanout153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 fanout154 (.A(net157),
    .X(net154));
 sky130_fd_sc_hd__buf_2 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 fanout157 (.A(\top0.cordic0.vec[1][2] ),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 fanout158 (.A(\top0.cordic0.vec[1][1] ),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 fanout159 (.A(\top0.cordic0.vec[1][1] ),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_4 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__buf_2 fanout161 (.A(\top0.cordic0.vec[1][1] ),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 fanout162 (.A(net167),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 fanout163 (.A(net167),
    .X(net163));
 sky130_fd_sc_hd__buf_2 fanout164 (.A(net167),
    .X(net164));
 sky130_fd_sc_hd__buf_2 fanout165 (.A(net167),
    .X(net165));
 sky130_fd_sc_hd__buf_2 fanout166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__buf_2 fanout167 (.A(\top0.cordic0.vec[1][0] ),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 fanout168 (.A(\top0.svm0.counter[14] ),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_4 fanout169 (.A(\top0.svm0.counter[10] ),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 fanout170 (.A(\top0.svm0.counter[7] ),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_4 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__buf_2 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(\top0.svm0.state[2] ),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_4 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_4 fanout175 (.A(\top0.cordic0.state[0] ),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_4 fanout176 (.A(net178),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_4 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__buf_2 fanout178 (.A(\top0.cordic0.state[0] ),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_4 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 fanout180 (.A(\top0.cordic0.gm0.iter[4] ),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 fanout181 (.A(\top0.cordic0.gm0.iter[4] ),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 fanout182 (.A(net186),
    .X(net182));
 sky130_fd_sc_hd__buf_2 fanout183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 fanout185 (.A(net186),
    .X(net185));
 sky130_fd_sc_hd__buf_2 fanout186 (.A(\top0.cordic0.gm0.iter[3] ),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_4 fanout188 (.A(\top0.cordic0.gm0.iter[2] ),
    .X(net188));
 sky130_fd_sc_hd__buf_2 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 fanout190 (.A(\top0.cordic0.gm0.iter[2] ),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_4 fanout191 (.A(net193),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_4 fanout193 (.A(\top0.cordic0.gm0.iter[1] ),
    .X(net193));
 sky130_fd_sc_hd__buf_2 fanout194 (.A(net196),
    .X(net194));
 sky130_fd_sc_hd__buf_2 fanout195 (.A(net196),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_4 fanout196 (.A(\top0.cordic0.gm0.iter[1] ),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 fanout197 (.A(net198),
    .X(net197));
 sky130_fd_sc_hd__buf_4 fanout198 (.A(net200),
    .X(net198));
 sky130_fd_sc_hd__buf_4 fanout199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__buf_2 fanout200 (.A(\top0.cordic0.gm0.iter[0] ),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_4 fanout201 (.A(net203),
    .X(net201));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_4 fanout203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_4 fanout204 (.A(\top0.cordic0.gm0.iter[0] ),
    .X(net204));
 sky130_fd_sc_hd__buf_2 fanout205 (.A(\top0.state[2] ),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_2 fanout206 (.A(\top0.state[2] ),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_4 fanout207 (.A(\top0.state[1] ),
    .X(net207));
 sky130_fd_sc_hd__buf_2 fanout208 (.A(\top0.state[0] ),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 fanout209 (.A(\top0.state[0] ),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_4 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__buf_2 fanout211 (.A(\top0.cordic0.domain[1] ),
    .X(net211));
 sky130_fd_sc_hd__buf_2 fanout212 (.A(\top0.cordic0.slte0.opA[15] ),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__buf_4 fanout214 (.A(\top0.cordic0.vec[0][17] ),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_4 fanout215 (.A(net217),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 fanout216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout217 (.A(net220),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_4 fanout218 (.A(net220),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 fanout219 (.A(net220),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 fanout220 (.A(\top0.cordic0.vec[0][17] ),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_8 fanout221 (.A(net224),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 fanout222 (.A(net224),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_4 fanout223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__buf_2 fanout224 (.A(\top0.cordic0.vec[0][16] ),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_4 fanout225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__buf_2 fanout226 (.A(\top0.cordic0.vec[0][15] ),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_4 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__buf_2 fanout228 (.A(\top0.cordic0.vec[0][15] ),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_8 fanout229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_4 fanout230 (.A(\top0.cordic0.vec[0][14] ),
    .X(net230));
 sky130_fd_sc_hd__buf_2 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_2 fanout233 (.A(\top0.cordic0.vec[0][14] ),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_8 fanout234 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_4 fanout235 (.A(net236),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_4 fanout236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_4 fanout237 (.A(\top0.cordic0.vec[0][13] ),
    .X(net237));
 sky130_fd_sc_hd__buf_4 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_2 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_8 fanout240 (.A(\top0.cordic0.vec[0][12] ),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_4 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__buf_2 fanout242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_2 fanout243 (.A(\top0.cordic0.vec[0][12] ),
    .X(net243));
 sky130_fd_sc_hd__buf_4 fanout244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__buf_4 fanout245 (.A(\top0.cordic0.vec[0][11] ),
    .X(net245));
 sky130_fd_sc_hd__buf_2 fanout246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 fanout247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__buf_4 fanout248 (.A(\top0.cordic0.vec[0][11] ),
    .X(net248));
 sky130_fd_sc_hd__buf_4 fanout249 (.A(\top0.cordic0.vec[0][10] ),
    .X(net249));
 sky130_fd_sc_hd__buf_2 fanout250 (.A(\top0.cordic0.vec[0][10] ),
    .X(net250));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(net252),
    .X(net251));
 sky130_fd_sc_hd__buf_6 fanout252 (.A(\top0.cordic0.vec[0][10] ),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_4 fanout253 (.A(net256),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_4 fanout254 (.A(net256),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_2 fanout255 (.A(net256),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_4 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_4 fanout257 (.A(\top0.cordic0.vec[0][9] ),
    .X(net257));
 sky130_fd_sc_hd__buf_4 fanout258 (.A(net261),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_4 fanout259 (.A(net261),
    .X(net259));
 sky130_fd_sc_hd__buf_1 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_4 fanout261 (.A(net262),
    .X(net261));
 sky130_fd_sc_hd__buf_4 fanout262 (.A(\top0.cordic0.vec[0][8] ),
    .X(net262));
 sky130_fd_sc_hd__buf_4 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__buf_4 fanout264 (.A(net268),
    .X(net264));
 sky130_fd_sc_hd__buf_4 fanout265 (.A(net268),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_2 fanout266 (.A(net268),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_4 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__buf_2 fanout268 (.A(\top0.cordic0.vec[0][7] ),
    .X(net268));
 sky130_fd_sc_hd__buf_4 fanout269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_4 fanout270 (.A(\top0.cordic0.vec[0][6] ),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_4 fanout271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__buf_2 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__buf_4 fanout273 (.A(\top0.cordic0.vec[0][6] ),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_4 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__buf_4 fanout275 (.A(net279),
    .X(net275));
 sky130_fd_sc_hd__buf_4 fanout276 (.A(net279),
    .X(net276));
 sky130_fd_sc_hd__buf_2 fanout277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__buf_4 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__buf_2 fanout279 (.A(\top0.cordic0.vec[0][5] ),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_4 fanout280 (.A(net284),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_2 fanout281 (.A(net284),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_4 fanout282 (.A(net284),
    .X(net282));
 sky130_fd_sc_hd__buf_2 fanout283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__buf_2 fanout284 (.A(\top0.cordic0.vec[0][4] ),
    .X(net284));
 sky130_fd_sc_hd__buf_4 fanout285 (.A(\top0.cordic0.vec[0][4] ),
    .X(net285));
 sky130_fd_sc_hd__buf_2 fanout286 (.A(\top0.cordic0.vec[0][4] ),
    .X(net286));
 sky130_fd_sc_hd__buf_2 fanout287 (.A(net293),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_2 fanout288 (.A(net293),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_4 fanout289 (.A(net293),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_4 fanout290 (.A(net293),
    .X(net290));
 sky130_fd_sc_hd__buf_4 fanout291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__buf_4 fanout292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_2 fanout293 (.A(\top0.cordic0.vec[0][3] ),
    .X(net293));
 sky130_fd_sc_hd__buf_2 fanout294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__buf_2 fanout295 (.A(net297),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_4 fanout296 (.A(net297),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_4 fanout297 (.A(\top0.cordic0.vec[0][2] ),
    .X(net297));
 sky130_fd_sc_hd__buf_2 fanout298 (.A(net299),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_4 fanout299 (.A(net301),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_4 fanout300 (.A(net301),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_4 fanout301 (.A(\top0.cordic0.vec[0][1] ),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_4 fanout302 (.A(net305),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_2 fanout303 (.A(net305),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_4 fanout304 (.A(net305),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_2 fanout305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_4 fanout306 (.A(\top0.cordic0.vec[0][0] ),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_8 fanout307 (.A(\top0.pid_d.mult0.b[15] ),
    .X(net307));
 sky130_fd_sc_hd__buf_2 fanout308 (.A(net309),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_4 fanout309 (.A(net310),
    .X(net309));
 sky130_fd_sc_hd__buf_4 fanout310 (.A(\top0.pid_d.mult0.b[14] ),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_4 fanout311 (.A(net312),
    .X(net311));
 sky130_fd_sc_hd__buf_2 fanout312 (.A(net313),
    .X(net312));
 sky130_fd_sc_hd__buf_2 fanout313 (.A(\top0.pid_d.mult0.b[13] ),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_4 fanout314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_4 fanout315 (.A(\top0.pid_d.mult0.b[12] ),
    .X(net315));
 sky130_fd_sc_hd__buf_2 fanout316 (.A(net317),
    .X(net316));
 sky130_fd_sc_hd__buf_2 fanout317 (.A(net318),
    .X(net317));
 sky130_fd_sc_hd__buf_1 fanout318 (.A(net319),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_4 fanout319 (.A(\top0.pid_d.mult0.b[11] ),
    .X(net319));
 sky130_fd_sc_hd__buf_2 fanout320 (.A(net1023),
    .X(net320));
 sky130_fd_sc_hd__buf_1 fanout321 (.A(net322),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_4 fanout322 (.A(\top0.pid_d.mult0.b[10] ),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_4 fanout323 (.A(net324),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_2 fanout324 (.A(net325),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_4 fanout325 (.A(net326),
    .X(net325));
 sky130_fd_sc_hd__buf_2 fanout326 (.A(\top0.pid_d.mult0.b[9] ),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_4 fanout327 (.A(net1022),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_2 fanout328 (.A(net329),
    .X(net328));
 sky130_fd_sc_hd__buf_4 fanout329 (.A(\top0.pid_d.mult0.b[8] ),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_4 fanout330 (.A(net331),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_8 fanout331 (.A(net332),
    .X(net331));
 sky130_fd_sc_hd__buf_4 fanout332 (.A(\top0.pid_d.mult0.b[7] ),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_4 fanout333 (.A(net335),
    .X(net333));
 sky130_fd_sc_hd__buf_4 fanout334 (.A(net336),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_2 fanout335 (.A(net336),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_4 fanout336 (.A(\top0.pid_d.mult0.b[6] ),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_4 fanout337 (.A(net339),
    .X(net337));
 sky130_fd_sc_hd__buf_4 fanout338 (.A(net339),
    .X(net338));
 sky130_fd_sc_hd__buf_4 fanout339 (.A(\top0.pid_d.mult0.b[5] ),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_4 fanout340 (.A(net342),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_4 fanout341 (.A(net342),
    .X(net341));
 sky130_fd_sc_hd__buf_4 fanout342 (.A(\top0.pid_d.mult0.b[4] ),
    .X(net342));
 sky130_fd_sc_hd__buf_2 fanout343 (.A(net344),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_4 fanout344 (.A(net345),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_4 fanout345 (.A(net346),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_4 fanout346 (.A(\top0.pid_d.mult0.b[3] ),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_4 fanout347 (.A(net348),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_4 fanout348 (.A(net350),
    .X(net348));
 sky130_fd_sc_hd__buf_2 fanout349 (.A(net350),
    .X(net349));
 sky130_fd_sc_hd__buf_2 fanout350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_4 fanout351 (.A(\top0.pid_d.mult0.b[2] ),
    .X(net351));
 sky130_fd_sc_hd__buf_2 fanout352 (.A(net354),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_2 fanout353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_4 fanout354 (.A(net355),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_4 fanout355 (.A(net356),
    .X(net355));
 sky130_fd_sc_hd__buf_4 fanout356 (.A(\top0.pid_d.mult0.b[1] ),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_4 fanout357 (.A(net358),
    .X(net357));
 sky130_fd_sc_hd__buf_2 fanout358 (.A(net359),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_4 fanout359 (.A(net360),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_4 fanout360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__buf_4 fanout361 (.A(\top0.pid_d.mult0.b[0] ),
    .X(net361));
 sky130_fd_sc_hd__buf_4 fanout362 (.A(net367),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_2 fanout363 (.A(net367),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_4 fanout364 (.A(net367),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_4 fanout365 (.A(net367),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_2 fanout366 (.A(net367),
    .X(net366));
 sky130_fd_sc_hd__buf_2 fanout367 (.A(\top0.pid_d.mult0.a[15] ),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_4 fanout368 (.A(\top0.pid_d.mult0.a[14] ),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_2 fanout369 (.A(\top0.pid_d.mult0.a[14] ),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_4 fanout370 (.A(\top0.pid_d.mult0.a[14] ),
    .X(net370));
 sky130_fd_sc_hd__buf_2 fanout371 (.A(net372),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_4 fanout372 (.A(\top0.pid_d.mult0.a[13] ),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_4 fanout373 (.A(\top0.pid_d.mult0.a[13] ),
    .X(net373));
 sky130_fd_sc_hd__buf_4 fanout374 (.A(net376),
    .X(net374));
 sky130_fd_sc_hd__buf_2 fanout375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__buf_4 fanout376 (.A(\top0.pid_d.mult0.a[12] ),
    .X(net376));
 sky130_fd_sc_hd__buf_2 fanout377 (.A(net379),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_4 fanout378 (.A(net379),
    .X(net378));
 sky130_fd_sc_hd__buf_2 fanout379 (.A(net380),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_4 fanout380 (.A(\top0.pid_d.mult0.a[11] ),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_4 fanout381 (.A(net382),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_4 fanout382 (.A(net384),
    .X(net382));
 sky130_fd_sc_hd__buf_4 fanout383 (.A(net384),
    .X(net383));
 sky130_fd_sc_hd__buf_2 fanout384 (.A(\top0.pid_d.mult0.a[10] ),
    .X(net384));
 sky130_fd_sc_hd__buf_2 fanout385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_2 fanout386 (.A(net387),
    .X(net386));
 sky130_fd_sc_hd__buf_2 fanout387 (.A(net389),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_4 fanout388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_4 fanout389 (.A(\top0.pid_d.mult0.a[9] ),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_4 fanout390 (.A(net391),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_4 fanout391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_4 fanout392 (.A(net394),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_4 fanout393 (.A(net394),
    .X(net393));
 sky130_fd_sc_hd__buf_2 fanout394 (.A(\top0.pid_d.mult0.a[8] ),
    .X(net394));
 sky130_fd_sc_hd__buf_2 fanout395 (.A(net397),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_4 fanout396 (.A(net397),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_2 fanout397 (.A(\top0.pid_d.mult0.a[7] ),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_4 fanout398 (.A(\top0.pid_d.mult0.a[7] ),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_2 fanout399 (.A(\top0.pid_d.mult0.a[7] ),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_4 fanout400 (.A(net401),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_2 fanout401 (.A(net402),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_2 fanout402 (.A(\top0.pid_d.mult0.a[6] ),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_4 fanout403 (.A(\top0.pid_d.mult0.a[6] ),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_4 fanout404 (.A(\top0.pid_d.mult0.a[6] ),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_4 fanout405 (.A(\top0.pid_d.mult0.a[5] ),
    .X(net405));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout406 (.A(\top0.pid_d.mult0.a[5] ),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_4 fanout407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_4 fanout408 (.A(\top0.pid_d.mult0.a[5] ),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_2 fanout409 (.A(\top0.pid_d.mult0.a[5] ),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_4 fanout410 (.A(net414),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_2 fanout411 (.A(net414),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_4 fanout412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_4 fanout413 (.A(net414),
    .X(net413));
 sky130_fd_sc_hd__buf_2 fanout414 (.A(\top0.pid_d.mult0.a[4] ),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_4 fanout415 (.A(net417),
    .X(net415));
 sky130_fd_sc_hd__buf_2 fanout416 (.A(net417),
    .X(net416));
 sky130_fd_sc_hd__buf_4 fanout417 (.A(\top0.pid_d.mult0.a[3] ),
    .X(net417));
 sky130_fd_sc_hd__buf_2 fanout418 (.A(net420),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_2 fanout419 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__buf_4 fanout420 (.A(net421),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_2 fanout421 (.A(\top0.pid_d.mult0.a[2] ),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_4 fanout422 (.A(net423),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_4 fanout423 (.A(net424),
    .X(net423));
 sky130_fd_sc_hd__buf_4 fanout424 (.A(\top0.pid_d.mult0.a[1] ),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_4 fanout425 (.A(net427),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_4 fanout426 (.A(net427),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_4 fanout427 (.A(\top0.pid_d.mult0.a[0] ),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_4 fanout428 (.A(\top0.matmul0.beta_pass[14] ),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_4 fanout429 (.A(net430),
    .X(net429));
 sky130_fd_sc_hd__buf_2 fanout430 (.A(\top0.matmul0.beta_pass[10] ),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_4 fanout431 (.A(\top0.pid_d.state[5] ),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_4 fanout432 (.A(net434),
    .X(net432));
 sky130_fd_sc_hd__buf_2 fanout433 (.A(net434),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_4 fanout434 (.A(\top0.pid_d.state[4] ),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_4 fanout435 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__buf_2 fanout436 (.A(\top0.pid_d.state[2] ),
    .X(net436));
 sky130_fd_sc_hd__buf_2 fanout437 (.A(net440),
    .X(net437));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout438 (.A(net440),
    .X(net438));
 sky130_fd_sc_hd__buf_2 fanout439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_2 fanout440 (.A(\top0.pid_d.state[2] ),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_4 fanout441 (.A(\top0.pid_d.state[1] ),
    .X(net441));
 sky130_fd_sc_hd__buf_2 fanout442 (.A(\top0.pid_d.state[1] ),
    .X(net442));
 sky130_fd_sc_hd__buf_4 fanout443 (.A(\top0.pid_q.mult0.b[15] ),
    .X(net443));
 sky130_fd_sc_hd__buf_4 fanout444 (.A(\top0.pid_q.mult0.b[15] ),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_4 fanout445 (.A(net446),
    .X(net445));
 sky130_fd_sc_hd__buf_4 fanout446 (.A(\top0.pid_q.mult0.b[14] ),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_4 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_4 fanout448 (.A(\top0.pid_q.mult0.b[13] ),
    .X(net448));
 sky130_fd_sc_hd__buf_4 fanout449 (.A(net451),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_2 fanout450 (.A(net451),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_4 fanout451 (.A(\top0.pid_q.mult0.b[12] ),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_4 fanout452 (.A(net454),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_2 fanout453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_4 fanout454 (.A(\top0.pid_q.mult0.b[11] ),
    .X(net454));
 sky130_fd_sc_hd__buf_4 fanout455 (.A(net457),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_4 fanout456 (.A(net457),
    .X(net456));
 sky130_fd_sc_hd__buf_4 fanout457 (.A(\top0.pid_q.mult0.b[10] ),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_4 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__buf_2 fanout459 (.A(net460),
    .X(net459));
 sky130_fd_sc_hd__buf_4 fanout460 (.A(\top0.pid_q.mult0.b[9] ),
    .X(net460));
 sky130_fd_sc_hd__buf_4 fanout461 (.A(net463),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_4 fanout462 (.A(\top0.pid_q.mult0.b[8] ),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_2 fanout463 (.A(\top0.pid_q.mult0.b[8] ),
    .X(net463));
 sky130_fd_sc_hd__buf_4 fanout464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_4 fanout465 (.A(\top0.pid_q.mult0.b[7] ),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_4 fanout466 (.A(net467),
    .X(net466));
 sky130_fd_sc_hd__buf_2 fanout467 (.A(\top0.pid_q.mult0.b[7] ),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_4 fanout468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__buf_2 fanout469 (.A(net470),
    .X(net469));
 sky130_fd_sc_hd__buf_4 fanout470 (.A(\top0.pid_q.mult0.b[6] ),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_4 fanout471 (.A(\top0.pid_q.mult0.b[5] ),
    .X(net471));
 sky130_fd_sc_hd__buf_2 fanout472 (.A(\top0.pid_q.mult0.b[5] ),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_4 fanout473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__buf_2 fanout474 (.A(\top0.pid_q.mult0.b[5] ),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_4 fanout475 (.A(net478),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_4 fanout476 (.A(net477),
    .X(net476));
 sky130_fd_sc_hd__buf_2 fanout477 (.A(net478),
    .X(net477));
 sky130_fd_sc_hd__buf_2 fanout478 (.A(\top0.pid_q.mult0.b[4] ),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_4 fanout479 (.A(net482),
    .X(net479));
 sky130_fd_sc_hd__buf_2 fanout480 (.A(net481),
    .X(net480));
 sky130_fd_sc_hd__buf_2 fanout481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_2 fanout482 (.A(net483),
    .X(net482));
 sky130_fd_sc_hd__buf_4 fanout483 (.A(\top0.pid_q.mult0.b[3] ),
    .X(net483));
 sky130_fd_sc_hd__buf_2 fanout484 (.A(net486),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_2 fanout485 (.A(net486),
    .X(net485));
 sky130_fd_sc_hd__buf_2 fanout486 (.A(net488),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_4 fanout487 (.A(net488),
    .X(net487));
 sky130_fd_sc_hd__buf_4 fanout488 (.A(\top0.pid_q.mult0.b[2] ),
    .X(net488));
 sky130_fd_sc_hd__buf_2 fanout489 (.A(net492),
    .X(net489));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout490 (.A(net492),
    .X(net490));
 sky130_fd_sc_hd__clkbuf_4 fanout491 (.A(net492),
    .X(net491));
 sky130_fd_sc_hd__buf_4 fanout492 (.A(\top0.pid_q.mult0.b[1] ),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_4 fanout493 (.A(net495),
    .X(net493));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout494 (.A(net496),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_4 fanout495 (.A(net496),
    .X(net495));
 sky130_fd_sc_hd__buf_4 fanout496 (.A(\top0.pid_q.mult0.b[0] ),
    .X(net496));
 sky130_fd_sc_hd__buf_4 fanout497 (.A(net498),
    .X(net497));
 sky130_fd_sc_hd__clkbuf_4 fanout498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__buf_4 fanout499 (.A(\top0.pid_q.mult0.a[15] ),
    .X(net499));
 sky130_fd_sc_hd__buf_4 fanout500 (.A(net502),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_2 fanout501 (.A(net502),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_4 fanout502 (.A(\top0.pid_q.mult0.a[14] ),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_4 fanout503 (.A(net504),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_2 fanout504 (.A(net505),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_4 fanout505 (.A(\top0.pid_q.mult0.a[13] ),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_8 fanout506 (.A(\top0.pid_q.mult0.a[12] ),
    .X(net506));
 sky130_fd_sc_hd__buf_2 fanout507 (.A(\top0.pid_q.mult0.a[12] ),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_4 fanout508 (.A(net509),
    .X(net508));
 sky130_fd_sc_hd__buf_2 fanout509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__buf_4 fanout510 (.A(\top0.pid_q.mult0.a[11] ),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_4 fanout511 (.A(net512),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_4 fanout512 (.A(net1029),
    .X(net512));
 sky130_fd_sc_hd__buf_2 fanout513 (.A(\top0.pid_q.mult0.a[10] ),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_4 fanout514 (.A(net515),
    .X(net514));
 sky130_fd_sc_hd__buf_2 fanout515 (.A(net516),
    .X(net515));
 sky130_fd_sc_hd__buf_4 fanout516 (.A(\top0.pid_q.mult0.a[9] ),
    .X(net516));
 sky130_fd_sc_hd__clkbuf_4 fanout517 (.A(net518),
    .X(net517));
 sky130_fd_sc_hd__buf_2 fanout518 (.A(net1028),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_2 fanout519 (.A(\top0.pid_q.mult0.a[8] ),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_4 fanout520 (.A(net521),
    .X(net520));
 sky130_fd_sc_hd__buf_4 fanout521 (.A(\top0.pid_q.mult0.a[7] ),
    .X(net521));
 sky130_fd_sc_hd__clkbuf_4 fanout522 (.A(net524),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_4 fanout523 (.A(net524),
    .X(net523));
 sky130_fd_sc_hd__clkbuf_4 fanout524 (.A(\top0.pid_q.mult0.a[6] ),
    .X(net524));
 sky130_fd_sc_hd__clkbuf_4 fanout525 (.A(net526),
    .X(net525));
 sky130_fd_sc_hd__buf_4 fanout526 (.A(net527),
    .X(net526));
 sky130_fd_sc_hd__buf_4 fanout527 (.A(\top0.pid_q.mult0.a[5] ),
    .X(net527));
 sky130_fd_sc_hd__buf_4 fanout528 (.A(\top0.pid_q.mult0.a[4] ),
    .X(net528));
 sky130_fd_sc_hd__clkbuf_2 fanout529 (.A(net530),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_2 fanout530 (.A(\top0.pid_q.mult0.a[4] ),
    .X(net530));
 sky130_fd_sc_hd__buf_4 fanout531 (.A(net533),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_2 fanout532 (.A(net533),
    .X(net532));
 sky130_fd_sc_hd__buf_4 fanout533 (.A(\top0.pid_q.mult0.a[3] ),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_4 fanout534 (.A(net535),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_4 fanout535 (.A(net536),
    .X(net535));
 sky130_fd_sc_hd__buf_2 fanout536 (.A(\top0.pid_q.mult0.a[2] ),
    .X(net536));
 sky130_fd_sc_hd__clkbuf_4 fanout537 (.A(net538),
    .X(net537));
 sky130_fd_sc_hd__buf_4 fanout538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__buf_4 fanout539 (.A(\top0.pid_q.mult0.a[1] ),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_4 fanout540 (.A(net541),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_4 fanout541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_4 fanout542 (.A(\top0.pid_q.mult0.a[0] ),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_4 fanout543 (.A(\top0.pid_q.state[5] ),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_4 fanout544 (.A(net545),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_4 fanout545 (.A(\top0.pid_q.state[4] ),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_4 fanout546 (.A(net547),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_4 fanout547 (.A(\top0.pid_q.state[3] ),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_4 fanout548 (.A(net549),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_4 fanout549 (.A(net552),
    .X(net549));
 sky130_fd_sc_hd__buf_2 fanout550 (.A(net552),
    .X(net550));
 sky130_fd_sc_hd__buf_2 fanout551 (.A(net552),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_2 fanout552 (.A(\top0.pid_q.state[2] ),
    .X(net552));
 sky130_fd_sc_hd__clkbuf_4 fanout553 (.A(\top0.pid_q.state[1] ),
    .X(net553));
 sky130_fd_sc_hd__buf_2 fanout554 (.A(\top0.pid_q.state[1] ),
    .X(net554));
 sky130_fd_sc_hd__buf_2 fanout555 (.A(\top0.svm0.delta[0] ),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_4 fanout556 (.A(net557),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_4 fanout557 (.A(net558),
    .X(net557));
 sky130_fd_sc_hd__clkbuf_4 fanout558 (.A(net561),
    .X(net558));
 sky130_fd_sc_hd__clkbuf_4 fanout559 (.A(net561),
    .X(net559));
 sky130_fd_sc_hd__buf_4 fanout560 (.A(net561),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_4 fanout561 (.A(\top0.matmul0.matmul_stage_inst.state[6] ),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_4 fanout562 (.A(net563),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_4 fanout563 (.A(\top0.matmul0.matmul_stage_inst.state[5] ),
    .X(net563));
 sky130_fd_sc_hd__buf_4 fanout564 (.A(\top0.matmul0.matmul_stage_inst.state[4] ),
    .X(net564));
 sky130_fd_sc_hd__buf_2 fanout565 (.A(\top0.matmul0.matmul_stage_inst.state[4] ),
    .X(net565));
 sky130_fd_sc_hd__clkbuf_4 fanout566 (.A(net567),
    .X(net566));
 sky130_fd_sc_hd__clkbuf_4 fanout567 (.A(\top0.matmul0.matmul_stage_inst.state[4] ),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_4 fanout568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_4 fanout569 (.A(\top0.matmul0.matmul_stage_inst.state[2] ),
    .X(net569));
 sky130_fd_sc_hd__buf_4 fanout570 (.A(\top0.matmul0.matmul_stage_inst.state[2] ),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_2 fanout571 (.A(\top0.matmul0.matmul_stage_inst.state[2] ),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_4 fanout572 (.A(net573),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_4 fanout573 (.A(\top0.matmul0.matmul_stage_inst.state[1] ),
    .X(net573));
 sky130_fd_sc_hd__clkbuf_4 fanout574 (.A(\top0.matmul0.matmul_stage_inst.state[1] ),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_2 fanout575 (.A(\top0.matmul0.matmul_stage_inst.state[1] ),
    .X(net575));
 sky130_fd_sc_hd__buf_4 fanout576 (.A(net577),
    .X(net576));
 sky130_fd_sc_hd__buf_4 fanout577 (.A(net606),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_4 fanout578 (.A(net579),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_4 fanout579 (.A(net586),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_4 fanout580 (.A(net581),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_2 fanout581 (.A(net585),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_4 fanout582 (.A(net584),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_4 fanout583 (.A(net584),
    .X(net583));
 sky130_fd_sc_hd__buf_2 fanout584 (.A(net585),
    .X(net584));
 sky130_fd_sc_hd__buf_2 fanout585 (.A(net586),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_2 fanout586 (.A(net606),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_4 fanout587 (.A(net589),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_4 fanout588 (.A(net589),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_4 fanout589 (.A(net606),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_4 fanout590 (.A(net598),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_4 fanout591 (.A(net598),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_4 fanout592 (.A(net597),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_4 fanout593 (.A(net597),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_4 fanout594 (.A(net596),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_4 fanout595 (.A(net596),
    .X(net595));
 sky130_fd_sc_hd__buf_2 fanout596 (.A(net597),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_2 fanout597 (.A(net598),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_2 fanout598 (.A(net605),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_4 fanout599 (.A(net600),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_4 fanout600 (.A(net605),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_4 fanout601 (.A(net602),
    .X(net601));
 sky130_fd_sc_hd__buf_2 fanout602 (.A(net605),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_4 fanout603 (.A(net605),
    .X(net603));
 sky130_fd_sc_hd__buf_2 fanout604 (.A(net605),
    .X(net604));
 sky130_fd_sc_hd__clkbuf_2 fanout605 (.A(net606),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_4 fanout606 (.A(net630),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_4 fanout607 (.A(net608),
    .X(net607));
 sky130_fd_sc_hd__clkbuf_2 fanout608 (.A(net630),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_4 fanout609 (.A(net630),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_4 fanout610 (.A(net630),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_4 fanout611 (.A(net612),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_4 fanout612 (.A(net615),
    .X(net612));
 sky130_fd_sc_hd__clkbuf_4 fanout613 (.A(net614),
    .X(net613));
 sky130_fd_sc_hd__buf_2 fanout614 (.A(net615),
    .X(net614));
 sky130_fd_sc_hd__buf_2 fanout615 (.A(net629),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_4 fanout616 (.A(net620),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_4 fanout617 (.A(net620),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_4 fanout618 (.A(net619),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_4 fanout619 (.A(net620),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_2 fanout620 (.A(net629),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_4 fanout621 (.A(net624),
    .X(net621));
 sky130_fd_sc_hd__buf_2 fanout622 (.A(net624),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_4 fanout623 (.A(net624),
    .X(net623));
 sky130_fd_sc_hd__buf_2 fanout624 (.A(net629),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_4 fanout625 (.A(net629),
    .X(net625));
 sky130_fd_sc_hd__buf_2 fanout626 (.A(net629),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_4 fanout627 (.A(net628),
    .X(net627));
 sky130_fd_sc_hd__clkbuf_2 fanout628 (.A(net629),
    .X(net628));
 sky130_fd_sc_hd__buf_2 fanout629 (.A(net630),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_4 fanout630 (.A(net2),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_4 fanout631 (.A(net635),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_4 fanout632 (.A(net634),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_4 fanout633 (.A(net634),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_4 fanout634 (.A(net635),
    .X(net634));
 sky130_fd_sc_hd__buf_2 fanout635 (.A(net654),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_4 fanout636 (.A(net638),
    .X(net636));
 sky130_fd_sc_hd__clkbuf_4 fanout637 (.A(net638),
    .X(net637));
 sky130_fd_sc_hd__clkbuf_4 fanout638 (.A(net639),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_4 fanout639 (.A(net654),
    .X(net639));
 sky130_fd_sc_hd__clkbuf_4 fanout640 (.A(net645),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_4 fanout641 (.A(net645),
    .X(net641));
 sky130_fd_sc_hd__clkbuf_4 fanout642 (.A(net645),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_2 fanout643 (.A(net645),
    .X(net643));
 sky130_fd_sc_hd__clkbuf_4 fanout644 (.A(net645),
    .X(net644));
 sky130_fd_sc_hd__clkbuf_4 fanout645 (.A(net654),
    .X(net645));
 sky130_fd_sc_hd__clkbuf_4 fanout646 (.A(net649),
    .X(net646));
 sky130_fd_sc_hd__clkbuf_4 fanout647 (.A(net649),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_2 fanout648 (.A(net649),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_2 fanout649 (.A(net654),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_4 fanout650 (.A(net653),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_4 fanout651 (.A(net653),
    .X(net651));
 sky130_fd_sc_hd__buf_2 fanout652 (.A(net653),
    .X(net652));
 sky130_fd_sc_hd__buf_2 fanout653 (.A(net654),
    .X(net653));
 sky130_fd_sc_hd__buf_2 fanout654 (.A(net687),
    .X(net654));
 sky130_fd_sc_hd__clkbuf_4 fanout655 (.A(net663),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_4 fanout656 (.A(net658),
    .X(net656));
 sky130_fd_sc_hd__clkbuf_4 fanout657 (.A(net658),
    .X(net657));
 sky130_fd_sc_hd__clkbuf_2 fanout658 (.A(net661),
    .X(net658));
 sky130_fd_sc_hd__clkbuf_4 fanout659 (.A(net660),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_4 fanout660 (.A(net661),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_2 fanout661 (.A(net663),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_4 fanout662 (.A(net663),
    .X(net662));
 sky130_fd_sc_hd__clkbuf_4 fanout663 (.A(net687),
    .X(net663));
 sky130_fd_sc_hd__buf_4 fanout664 (.A(net666),
    .X(net664));
 sky130_fd_sc_hd__clkbuf_4 fanout665 (.A(net666),
    .X(net665));
 sky130_fd_sc_hd__clkbuf_4 fanout666 (.A(net669),
    .X(net666));
 sky130_fd_sc_hd__clkbuf_4 fanout667 (.A(net669),
    .X(net667));
 sky130_fd_sc_hd__clkbuf_4 fanout668 (.A(net669),
    .X(net668));
 sky130_fd_sc_hd__buf_2 fanout669 (.A(net687),
    .X(net669));
 sky130_fd_sc_hd__clkbuf_4 fanout670 (.A(net673),
    .X(net670));
 sky130_fd_sc_hd__clkbuf_4 fanout671 (.A(net673),
    .X(net671));
 sky130_fd_sc_hd__buf_2 fanout672 (.A(net673),
    .X(net672));
 sky130_fd_sc_hd__clkbuf_2 fanout673 (.A(net674),
    .X(net673));
 sky130_fd_sc_hd__clkbuf_2 fanout674 (.A(net675),
    .X(net674));
 sky130_fd_sc_hd__clkbuf_4 fanout675 (.A(net687),
    .X(net675));
 sky130_fd_sc_hd__clkbuf_4 fanout676 (.A(net686),
    .X(net676));
 sky130_fd_sc_hd__clkbuf_4 fanout677 (.A(net678),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_4 fanout678 (.A(net679),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_4 fanout679 (.A(net686),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_4 fanout680 (.A(net681),
    .X(net680));
 sky130_fd_sc_hd__clkbuf_4 fanout681 (.A(net686),
    .X(net681));
 sky130_fd_sc_hd__clkbuf_4 fanout682 (.A(net685),
    .X(net682));
 sky130_fd_sc_hd__buf_2 fanout683 (.A(net685),
    .X(net683));
 sky130_fd_sc_hd__clkbuf_4 fanout684 (.A(net685),
    .X(net684));
 sky130_fd_sc_hd__buf_2 fanout685 (.A(net686),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_4 fanout686 (.A(net687),
    .X(net686));
 sky130_fd_sc_hd__clkbuf_8 fanout687 (.A(net2),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_4 fanout688 (.A(net689),
    .X(net688));
 sky130_fd_sc_hd__clkbuf_2 fanout689 (.A(net693),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_4 fanout690 (.A(net692),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_2 fanout691 (.A(net692),
    .X(net691));
 sky130_fd_sc_hd__buf_2 fanout692 (.A(net693),
    .X(net692));
 sky130_fd_sc_hd__buf_2 fanout693 (.A(net700),
    .X(net693));
 sky130_fd_sc_hd__clkbuf_4 fanout694 (.A(net695),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_4 fanout695 (.A(net696),
    .X(net695));
 sky130_fd_sc_hd__buf_2 fanout696 (.A(net700),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_4 fanout697 (.A(net700),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_4 fanout698 (.A(net699),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_4 fanout699 (.A(net700),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_2 fanout700 (.A(net1),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk_sys (.A(clknet_3_2__leaf_clk_sys),
    .X(clknet_leaf_0_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk_sys (.A(clknet_3_2__leaf_clk_sys),
    .X(clknet_leaf_1_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk_sys (.A(clknet_3_2__leaf_clk_sys),
    .X(clknet_leaf_2_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk_sys (.A(clknet_3_2__leaf_clk_sys),
    .X(clknet_leaf_3_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk_sys (.A(clknet_3_0__leaf_clk_sys),
    .X(clknet_leaf_4_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk_sys (.A(clknet_3_0__leaf_clk_sys),
    .X(clknet_leaf_5_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk_sys (.A(clknet_3_2__leaf_clk_sys),
    .X(clknet_leaf_6_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk_sys (.A(clknet_3_2__leaf_clk_sys),
    .X(clknet_leaf_7_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk_sys (.A(clknet_3_2__leaf_clk_sys),
    .X(clknet_leaf_8_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk_sys (.A(clknet_3_2__leaf_clk_sys),
    .X(clknet_leaf_9_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_10_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_11_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_12_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_13_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_14_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_15_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk_sys (.A(clknet_3_2__leaf_clk_sys),
    .X(clknet_leaf_16_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk_sys (.A(clknet_3_2__leaf_clk_sys),
    .X(clknet_leaf_17_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_18_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk_sys (.A(clknet_3_2__leaf_clk_sys),
    .X(clknet_leaf_20_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk_sys (.A(clknet_3_2__leaf_clk_sys),
    .X(clknet_leaf_21_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk_sys (.A(clknet_3_2__leaf_clk_sys),
    .X(clknet_leaf_22_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_23_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_24_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_25_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_26_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_27_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_28_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_29_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_30_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_31_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk_sys (.A(clknet_3_6__leaf_clk_sys),
    .X(clknet_leaf_32_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk_sys (.A(clknet_3_6__leaf_clk_sys),
    .X(clknet_leaf_33_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk_sys (.A(clknet_3_7__leaf_clk_sys),
    .X(clknet_leaf_36_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk_sys (.A(clknet_3_7__leaf_clk_sys),
    .X(clknet_leaf_37_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk_sys (.A(clknet_3_7__leaf_clk_sys),
    .X(clknet_leaf_38_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk_sys (.A(clknet_3_7__leaf_clk_sys),
    .X(clknet_leaf_39_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk_sys (.A(clknet_3_7__leaf_clk_sys),
    .X(clknet_leaf_40_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk_sys (.A(clknet_3_7__leaf_clk_sys),
    .X(clknet_leaf_41_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk_sys (.A(clknet_3_7__leaf_clk_sys),
    .X(clknet_leaf_42_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk_sys (.A(clknet_3_7__leaf_clk_sys),
    .X(clknet_leaf_43_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk_sys (.A(clknet_3_7__leaf_clk_sys),
    .X(clknet_leaf_44_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk_sys (.A(clknet_3_7__leaf_clk_sys),
    .X(clknet_leaf_45_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk_sys (.A(clknet_3_7__leaf_clk_sys),
    .X(clknet_leaf_46_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk_sys (.A(clknet_3_7__leaf_clk_sys),
    .X(clknet_leaf_47_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk_sys (.A(clknet_3_7__leaf_clk_sys),
    .X(clknet_leaf_48_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk_sys (.A(clknet_3_6__leaf_clk_sys),
    .X(clknet_leaf_49_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk_sys (.A(clknet_3_6__leaf_clk_sys),
    .X(clknet_leaf_50_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk_sys (.A(clknet_3_6__leaf_clk_sys),
    .X(clknet_leaf_51_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk_sys (.A(clknet_3_6__leaf_clk_sys),
    .X(clknet_leaf_52_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk_sys (.A(clknet_3_6__leaf_clk_sys),
    .X(clknet_leaf_53_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk_sys (.A(clknet_3_6__leaf_clk_sys),
    .X(clknet_leaf_54_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk_sys (.A(clknet_3_4__leaf_clk_sys),
    .X(clknet_leaf_55_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk_sys (.A(clknet_3_6__leaf_clk_sys),
    .X(clknet_leaf_56_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk_sys (.A(clknet_3_4__leaf_clk_sys),
    .X(clknet_leaf_57_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk_sys (.A(clknet_3_4__leaf_clk_sys),
    .X(clknet_leaf_58_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk_sys (.A(clknet_3_4__leaf_clk_sys),
    .X(clknet_leaf_59_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk_sys (.A(clknet_3_4__leaf_clk_sys),
    .X(clknet_leaf_60_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk_sys (.A(clknet_3_4__leaf_clk_sys),
    .X(clknet_leaf_61_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk_sys (.A(clknet_3_4__leaf_clk_sys),
    .X(clknet_leaf_62_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk_sys (.A(clknet_3_4__leaf_clk_sys),
    .X(clknet_leaf_63_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk_sys (.A(clknet_3_5__leaf_clk_sys),
    .X(clknet_leaf_64_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk_sys (.A(clknet_3_5__leaf_clk_sys),
    .X(clknet_leaf_65_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk_sys (.A(clknet_3_5__leaf_clk_sys),
    .X(clknet_leaf_66_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk_sys (.A(clknet_3_5__leaf_clk_sys),
    .X(clknet_leaf_67_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk_sys (.A(clknet_3_5__leaf_clk_sys),
    .X(clknet_leaf_68_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk_sys (.A(clknet_3_5__leaf_clk_sys),
    .X(clknet_leaf_69_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk_sys (.A(clknet_3_5__leaf_clk_sys),
    .X(clknet_leaf_70_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk_sys (.A(clknet_3_5__leaf_clk_sys),
    .X(clknet_leaf_71_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk_sys (.A(clknet_3_5__leaf_clk_sys),
    .X(clknet_leaf_72_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk_sys (.A(clknet_3_5__leaf_clk_sys),
    .X(clknet_leaf_73_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk_sys (.A(clknet_3_5__leaf_clk_sys),
    .X(clknet_leaf_74_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk_sys (.A(clknet_3_4__leaf_clk_sys),
    .X(clknet_leaf_75_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk_sys (.A(clknet_3_4__leaf_clk_sys),
    .X(clknet_leaf_76_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_77_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_78_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_79_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_80_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk_sys (.A(clknet_3_4__leaf_clk_sys),
    .X(clknet_leaf_81_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk_sys (.A(clknet_3_4__leaf_clk_sys),
    .X(clknet_leaf_82_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk_sys (.A(clknet_3_4__leaf_clk_sys),
    .X(clknet_leaf_83_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_84_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_85_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_86_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_87_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_88_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk_sys (.A(clknet_3_3__leaf_clk_sys),
    .X(clknet_leaf_89_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_90_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_91_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_92_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_93_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk_sys (.A(clknet_3_0__leaf_clk_sys),
    .X(clknet_leaf_94_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_96_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_97_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_98_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk_sys (.A(clknet_3_1__leaf_clk_sys),
    .X(clknet_leaf_99_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk_sys (.A(clknet_3_0__leaf_clk_sys),
    .X(clknet_leaf_100_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk_sys (.A(clknet_3_0__leaf_clk_sys),
    .X(clknet_leaf_101_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk_sys (.A(clknet_3_0__leaf_clk_sys),
    .X(clknet_leaf_102_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk_sys (.A(clknet_3_0__leaf_clk_sys),
    .X(clknet_leaf_103_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk_sys (.A(clknet_3_0__leaf_clk_sys),
    .X(clknet_leaf_104_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk_sys (.A(clknet_3_0__leaf_clk_sys),
    .X(clknet_leaf_105_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk_sys (.A(clknet_3_0__leaf_clk_sys),
    .X(clknet_leaf_106_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk_sys (.A(clknet_3_0__leaf_clk_sys),
    .X(clknet_leaf_107_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk_sys (.A(clknet_3_0__leaf_clk_sys),
    .X(clknet_leaf_108_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk_sys (.A(clknet_3_2__leaf_clk_sys),
    .X(clknet_leaf_109_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk_sys (.A(clknet_3_2__leaf_clk_sys),
    .X(clknet_leaf_110_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_sys (.A(clk_sys),
    .X(clknet_0_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk_sys (.A(clknet_0_clk_sys),
    .X(clknet_3_0__leaf_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk_sys (.A(clknet_0_clk_sys),
    .X(clknet_3_1__leaf_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk_sys (.A(clknet_0_clk_sys),
    .X(clknet_3_2__leaf_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk_sys (.A(clknet_0_clk_sys),
    .X(clknet_3_3__leaf_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk_sys (.A(clknet_0_clk_sys),
    .X(clknet_3_4__leaf_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk_sys (.A(clknet_0_clk_sys),
    .X(clknet_3_5__leaf_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk_sys (.A(clknet_0_clk_sys),
    .X(clknet_3_6__leaf_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk_sys (.A(clknet_0_clk_sys),
    .X(clknet_3_7__leaf_clk_sys));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_mosi (.A(clk_mosi),
    .X(clknet_0_clk_mosi));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk_mosi (.A(clknet_0_clk_mosi),
    .X(clknet_3_0__leaf_clk_mosi));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk_mosi (.A(clknet_0_clk_mosi),
    .X(clknet_3_1__leaf_clk_mosi));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk_mosi (.A(clknet_0_clk_mosi),
    .X(clknet_3_2__leaf_clk_mosi));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk_mosi (.A(clknet_0_clk_mosi),
    .X(clknet_3_3__leaf_clk_mosi));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk_mosi (.A(clknet_0_clk_mosi),
    .X(clknet_3_4__leaf_clk_mosi));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk_mosi (.A(clknet_0_clk_mosi),
    .X(clknet_3_5__leaf_clk_mosi));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk_mosi (.A(clknet_0_clk_mosi),
    .X(clknet_3_6__leaf_clk_mosi));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk_mosi (.A(clknet_0_clk_mosi),
    .X(clknet_3_7__leaf_clk_mosi));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\spi0.cs_sync[0] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\spi0.cs_sync[1] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\top0.kpq[13] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net4),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(_00439_),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net6),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_00441_),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net5),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_00440_),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\top0.kpq[12] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\top0.matmul0.matmul_stage_inst.b[15] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\top0.cordic0.sin[3] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\top0.kpq[11] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\top0.matmul0.matmul_stage_inst.c[13] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\top0.cordic0.cos[1] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\top0.matmul0.matmul_stage_inst.a[7] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\top0.matmul0.matmul_stage_inst.a[4] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\top0.cordic0.cos[3] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\top0.kpq[6] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\top0.cordic0.sin[9] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\top0.cordic0.sin[1] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\top0.pid_d.curr_error[15] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_00325_),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\top0.cordic0.sin[8] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\top0.matmul0.matmul_stage_inst.d[7] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\top0.cordic0.sin[6] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\top0.cordic0.sin[4] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\top0.pid_q.prev_error[14] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\top0.svm0.tB[0] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\top0.matmul0.matmul_stage_inst.a[13] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\top0.cordic0.cos[4] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\top0.cordic0.cos[0] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\top0.cordic0.sin[11] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\top0.kpq[9] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\top0.matmul0.matmul_stage_inst.c[6] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\top0.svm0.tC[0] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\top0.periodTop[15] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\top0.cordic0.cos[6] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\top0.matmul0.matmul_stage_inst.d[8] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\top0.cordic0.sin[13] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\top0.periodTop[4] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\top0.matmul0.matmul_stage_inst.d[13] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\top0.c_out_calc[5] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\state[1] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\top0.cordic0.sin[0] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\top0.matmul0.matmul_stage_inst.d[12] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\top0.matmul0.matmul_stage_inst.d[4] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\top0.matmul0.matmul_stage_inst.start ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\top0.cordic0.sin[2] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\top0.matmul0.matmul_stage_inst.d[2] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\top0.kpq[4] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\top0.matmul0.matmul_stage_inst.d[11] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\top0.matmul0.matmul_stage_inst.d[10] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\top0.periodTop[14] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\top0.matmul0.matmul_stage_inst.d[6] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\top0.cordic0.cos[2] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\top0.kpq[1] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\top0.pid_q.prev_error[15] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\top0.matmul0.matmul_stage_inst.d[0] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\top0.pid_d.curr_error[11] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\top0.cordic0.cos[12] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\top0.cordic0.cos[5] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\top0.cordic0.cos[7] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\top0.matmul0.matmul_stage_inst.b[6] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\top0.pid_d.curr_error[14] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_00324_),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\top0.matmul0.matmul_stage_inst.a[5] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\top0.matmul0.matmul_stage_inst.a[1] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\top0.cordic0.sin[7] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\top0.matmul0.matmul_stage_inst.a[3] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\top0.cordic0.cos[8] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\top0.pid_q.curr_int[15] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_00434_),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\top0.svm0.tB[10] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\top0.kpq[7] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\top0.svm0.tB[7] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\top0.svm0.tA[13] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\top0.matmul0.matmul_stage_inst.b[14] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\top0.matmul0.matmul_stage_inst.c[7] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\top0.svm0.tA[6] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\top0.svm0.tA[10] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\top0.periodTop[3] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\top0.svm0.tA[2] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\top0.matmul0.matmul_stage_inst.b[4] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\top0.cordic0.cos[9] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\top0.matmul0.matmul_stage_inst.b[13] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\top0.kpq[2] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\top0.svm0.tA[7] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\top0.kpq[3] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\top0.svm0.tB[11] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\top0.matmul0.matmul_stage_inst.c[8] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\top0.matmul0.matmul_stage_inst.b[7] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\top0.kpq[5] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\top0.cordic0.cos[10] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\top0.svm0.tA[1] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\top0.kpq[10] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\top0.svm0.tB[9] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\top0.c_out_calc[2] ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\top0.matmul0.matmul_stage_inst.c[5] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\top0.svm0.tA[15] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\top0.c_out_calc[8] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\top0.currT_r[15] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\top0.kpq[14] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\top0.svm0.tB[13] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\top0.matmul0.matmul_stage_inst.c[9] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\top0.svm0.tA[11] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\top0.svm0.tC[10] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\top0.matmul0.matmul_stage_inst.b[10] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\top0.svm0.tB[12] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\top0.svm0.tC[7] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\top0.svm0.tA[3] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\top0.pid_q.prev_error[8] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\top0.matmul0.matmul_stage_inst.b[12] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\top0.svm0.tB[8] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\top0.pid_d.prev_int[15] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_00132_),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\top0.svm0.tC[9] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\top0.pid_q.prev_error[7] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\top0.matmul0.matmul_stage_inst.b[3] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\top0.pid_q.prev_error[9] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\top0.svm0.tB[5] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\top0.matmul0.matmul_stage_inst.c[4] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\top0.svm0.tB[4] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\top0.svm0.tC[14] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\top0.matmul0.matmul_stage_inst.c[11] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\top0.pid_q.prev_error[10] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\top0.kpq[8] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\top0.pid_d.curr_int[10] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_00127_),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\top0.svm0.tA[0] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\top0.svm0.tB[1] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\top0.periodTop[11] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\top0.c_out_calc[0] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\top0.svm0.tB[6] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\top0.svm0.tB[2] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\top0.matmul0.matmul_stage_inst.d[5] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\top0.svm0.tB[3] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\top0.svm0.tB[14] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\top0.svm0.tB[15] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\top0.c_out_calc[10] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\top0.matmul0.matmul_stage_inst.c[12] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\top0.pid_q.prev_error[6] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\top0.kpq[0] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\top0.c_out_calc[11] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\top0.periodTop[5] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\top0.matmul0.matmul_stage_inst.d[1] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\top0.matmul0.matmul_stage_inst.c[3] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\top0.svm0.tC[8] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\top0.pid_q.prev_error[5] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\top0.matmul0.matmul_stage_inst.d[9] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\top0.svm0.tC[13] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\top0.svm0.tC[1] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\top0.svm0.tC[2] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\top0.matmul0.matmul_stage_inst.c[10] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\top0.svm0.tC[3] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\top0.matmul0.matmul_stage_inst.b[8] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\top0.svm0.tC[11] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\top0.svm0.tC[15] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\top0.matmul0.matmul_stage_inst.c[2] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\top0.pid_q.prev_error[4] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\top0.svm0.tC[6] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\top0.matmul0.matmul_stage_inst.b[0] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\top0.cordic0.cos[13] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\top0.svm0.tC[5] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\top0.pid_q.curr_error[14] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\top0.matmul0.matmul_stage_inst.b[5] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\top0.c_out_calc[6] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\top0.svm0.tC[12] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\top0.svm0.tC[4] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\top0.matmul0.matmul_stage_inst.c[1] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\top0.matmul0.matmul_stage_inst.b[2] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\top0.pid_d.prev_error[3] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\top0.pid_q.prev_error[13] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\top0.pid_d.prev_error[10] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_00320_),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\top0.pid_d.prev_error[8] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_00318_),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\top0.pid_d.prev_error[4] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\top0.pid_d.prev_error[6] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\top0.pid_d.prev_error[7] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_00317_),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\top0.svm0.tA[12] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\top0.svm0.tA[4] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\top0.pid_d.prev_error[5] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\top0.pid_q.curr_error[15] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\top0.periodTop[13] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\top0.matmul0.matmul_stage_inst.b[1] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\top0.c_out_calc[7] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\top0.pid_d.prev_error[9] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_00319_),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\top0.matmul0.matmul_stage_inst.b[11] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\top0.pid_d.prev_error[2] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_00312_),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\top0.svm0.tA[5] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\top0.periodTop[12] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\top0.svm0.delta[2] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\top0.pid_q.prev_error[2] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\top0.pid_q.prev_error[11] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\top0.pid_q.prev_error[3] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\top0.periodTop[10] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\top0.cordic0.slte0.opA[0] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\top0.svm0.calc_ready ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\top0.pid_d.prev_error[12] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_00322_),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\top0.currT_r[5] ),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\top0.matmul0.matmul_stage_inst.b[9] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\top0.currT_r[0] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\top0.svm0.tA[14] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\top0.pid_q.prev_error[12] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\top0.pid_d.curr_error[13] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\top0.pid_d.curr_int[7] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_00124_),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\top0.cordic0.slte0.opA[10] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\top0.pid_q.prev_int[11] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\top0.cordic0.out_valid ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\top0.c_out_calc[14] ),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\top0.pid_d.prev_int[13] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\top0.currT_r[4] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\top0.currT_r[1] ),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\top0.cordic0.sin[5] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\top0.c_out_calc[15] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\top0.currT_r[12] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\top0.pid_d.curr_error[8] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\top0.pid_q.curr_int[8] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\spi0.data_packed[44] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_05378_),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\top0.pid_d.curr_error[7] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\top0.cordic0.sin[10] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\top0.pid_q.curr_error[4] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\top0.svm0.tA[8] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\top0.pid_d.curr_error[10] ),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\top0.cordic0.slte0.opA[8] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\top0.svm0.delta[7] ),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\top0.currT_r[3] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\top0.currT_r[11] ),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\top0.c_out_calc[13] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\top0.kpq[15] ),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\top0.pid_d.prev_int[6] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\top0.c_out_calc[12] ),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\top0.pid_d.curr_error[0] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\top0.pid_d.prev_int[14] ),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\spi0.data_packed[43] ),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\top0.matmul0.b[15] ),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\spi0.data_packed[34] ),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_05368_),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\spi0.data_packed[40] ),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_05374_),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\top0.currT_r[8] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\spi0.data_packed[45] ),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_05379_),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\top0.matmul0.b[10] ),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\top0.currT_r[9] ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\spi0.data_packed[38] ),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_05372_),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\top0.svm0.delta[6] ),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\spi0.data_packed[42] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_05375_),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\spi0.data_packed[33] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\top0.svm0.delta[11] ),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\top0.currT_r[6] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\top0.pid_d.prev_error[1] ),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\top0.currT_r[7] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\spi0.opcode[7] ),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\top0.pid_d.prev_int[4] ),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\top0.b_in_matmul[5] ),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\top0.b_in_matmul[6] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\spi0.data_packed[39] ),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\top0.pid_d.prev_int[0] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\spi0.data_packed[46] ),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\top0.pid_q.prev_int[9] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\top0.pid_d.prev_int[2] ),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\top0.svm0.delta[12] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\spi0.data_packed[37] ),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_05370_),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\spi0.data_packed[35] ),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\top0.pid_q.prev_int[7] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\top0.pid_q.prev_int[3] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\top0.pid_d.curr_int[12] ),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\top0.a_in_matmul[2] ),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\top0.b_in_matmul[11] ),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\top0.cordic0.slte0.opA[4] ),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\top0.pid_q.prev_int[4] ),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\top0.pid_q.curr_error[1] ),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\top0.pid_q.prev_error[0] ),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\top0.a_in_matmul[8] ),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\top0.pid_d.curr_error[2] ),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\top0.matmul0.a[3] ),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\top0.pid_q.prev_int[10] ),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\top0.svm0.tA[9] ),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\top0.pid_d.prev_int[9] ),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\top0.pid_q.prev_int[0] ),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\top0.cordic0.slte0.opA[2] ),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\top0.matmul0.matmul_stage_inst.a[0] ),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\top0.b_in_matmul[14] ),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\top0.pid_q.prev_int[2] ),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\top0.cordic0.sin[12] ),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\top0.matmul0.state[0] ),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\top0.b_in_matmul[1] ),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\top0.cordic0.sin[9] ),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\top0.cordic0.sin[7] ),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\top0.cordic0.sin[8] ),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\top0.cordic0.cos[4] ),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\top0.cordic0.sin[1] ),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\top0.b_in_matmul[5] ),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\top0.cordic0.sin[6] ),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\top0.periodTop[15] ),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\top0.cordic0.sin[13] ),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\top0.cordic0.cos[6] ),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\top0.b_in_matmul[14] ),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\top0.cordic0.sin[3] ),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\spi0.data_packed[43] ),
    .X(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_01123_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_02352_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_02367_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_03020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_05444_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_09593_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_12739_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_12739_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_12739_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_12812_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\top0.periodTop_r[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\top0.pid_d.state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\top0.svm0.out_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_08403_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_10561_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_11094_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\top0.c_out_calc[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\top0.matmul0.matmul_stage_inst.e[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net687));
 sky130_fd_sc_hd__clkbuf_1 wire1 (.A(_11850_),
    .X(net1012));
 sky130_fd_sc_hd__buf_4 fanout2 (.A(_11548_),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_4 fanout3 (.A(_11439_),
    .X(net1014));
 sky130_fd_sc_hd__buf_4 fanout4 (.A(_05518_),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_4 fanout5 (.A(_11517_),
    .X(net1016));
 sky130_fd_sc_hd__buf_4 fanout6 (.A(_03020_),
    .X(net1017));
 sky130_fd_sc_hd__buf_2 fanout7 (.A(_08403_),
    .X(net1018));
 sky130_fd_sc_hd__buf_4 fanout8 (.A(_05444_),
    .X(net1019));
 sky130_fd_sc_hd__buf_4 fanout9 (.A(_11651_),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_4 fanout10 (.A(_12744_),
    .X(net1021));
 sky130_fd_sc_hd__buf_4 fanout11 (.A(net328),
    .X(net1022));
 sky130_fd_sc_hd__buf_4 fanout12 (.A(net321),
    .X(net1023));
 sky130_fd_sc_hd__clkbuf_8 fanout13 (.A(net75),
    .X(net1024));
 sky130_fd_sc_hd__buf_4 fanout14 (.A(net55),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_4 fanout15 (.A(net530),
    .X(net1026));
 sky130_fd_sc_hd__buf_4 fanout16 (.A(net53),
    .X(net1027));
 sky130_fd_sc_hd__buf_4 fanout17 (.A(net519),
    .X(net1028));
 sky130_fd_sc_hd__buf_4 fanout701 (.A(net513),
    .X(net1029));
 sky130_fd_sc_hd__buf_4 fanout702 (.A(net29),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_8 fanout703 (.A(net117),
    .X(net1031));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_812 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_870 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_983 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1087 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1066 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1095 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1064 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_871 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1064 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_190_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_194_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1193 ();
endmodule
