VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_wrapper
  CLASS BLOCK ;
  FOREIGN fpga_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 563.495 BY 574.215 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 563.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 563.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 563.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 563.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 557.760 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 557.760 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 557.760 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 489.570 557.760 491.170 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 563.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 563.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 563.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 563.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 557.760 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 557.760 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 557.760 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 557.760 487.870 ;
    END
  END VPWR
  PIN clk_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 559.495 231.240 563.495 231.840 ;
    END
  END clk_mosi
  PIN clk_sys
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END clk_sys
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 559.495 234.640 563.495 235.240 ;
    END
  END cs
  PIN pwmA
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 418.690 570.215 418.970 574.215 ;
    END
  END pwmA
  PIN pwmB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 405.810 570.215 406.090 574.215 ;
    END
  END pwmB
  PIN pwmC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 409.030 570.215 409.310 574.215 ;
    END
  END pwmC
  PIN ready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 559.495 285.640 563.495 286.240 ;
    END
  END ready
  PIN rstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END rstb
  PIN spi_mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END spi_mosi
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 557.520 563.125 ;
      LAYER met1 ;
        RECT 4.670 10.640 558.830 563.280 ;
      LAYER met2 ;
        RECT 4.690 569.935 405.530 570.930 ;
        RECT 406.370 569.935 408.750 570.930 ;
        RECT 409.590 569.935 418.410 570.930 ;
        RECT 419.250 569.935 558.810 570.930 ;
        RECT 4.690 10.695 558.810 569.935 ;
      LAYER met3 ;
        RECT 4.000 545.040 559.495 563.205 ;
        RECT 4.400 543.640 559.495 545.040 ;
        RECT 4.000 541.640 559.495 543.640 ;
        RECT 4.400 540.240 559.495 541.640 ;
        RECT 4.000 286.640 559.495 540.240 ;
        RECT 4.000 285.240 559.095 286.640 ;
        RECT 4.000 279.840 559.495 285.240 ;
        RECT 4.400 278.440 559.495 279.840 ;
        RECT 4.000 235.640 559.495 278.440 ;
        RECT 4.000 234.240 559.095 235.640 ;
        RECT 4.000 232.240 559.495 234.240 ;
        RECT 4.000 230.840 559.095 232.240 ;
        RECT 4.000 10.715 559.495 230.840 ;
      LAYER met4 ;
        RECT 23.295 27.375 23.940 553.345 ;
        RECT 26.340 27.375 174.240 553.345 ;
        RECT 176.640 27.375 177.540 553.345 ;
        RECT 179.940 27.375 327.840 553.345 ;
        RECT 330.240 27.375 331.140 553.345 ;
        RECT 333.540 27.375 481.440 553.345 ;
        RECT 483.840 27.375 484.740 553.345 ;
        RECT 487.140 27.375 490.065 553.345 ;
  END
END fpga_wrapper
END LIBRARY

